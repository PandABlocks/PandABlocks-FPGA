library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.support.all;

entity pulse is
port (
    -- Clock and Reset
    clk_i               : in  std_logic;
    -- Block Input and Outputs
    trig_i              : in  std_logic;
    enable_i            : in  std_logic;
    out_o               : out std_logic;
    -- Block Parameters
    TRIG_EDGE           : in  std_logic_vector(31 downto 0) := (others => '0');
    TRIG_EDGE_WSTB      : in  std_logic;
    DELAY_L             : in  std_logic_vector(31 downto 0);
    DELAY_L_WSTB        : in  std_logic;
    DELAY_H             : in  std_logic_vector(31 downto 0);
    DELAY_H_WSTB        : in  std_logic;
    WIDTH_L             : in  std_logic_vector(31 downto 0);
    WIDTH_L_WSTB        : in  std_logic;
    WIDTH_H             : in  std_logic_vector(31 downto 0);
    WIDTH_H_WSTB        : in  std_logic;
    PULSES              : in  std_logic_vector(31 downto 0) := (others => '0');
    PULSES_WSTB         : in  std_logic;
    STEP_L              : in  std_logic_vector(31 downto 0);
    STEP_L_WSTB         : in  std_logic;
    STEP_H              : in  std_logic_vector(31 downto 0);
    STEP_H_WSTB         : in  std_logic;
    -- Block Status
    QUEUED              : out std_logic_vector(31 downto 0);
    DROPPED             : out std_logic_vector(31 downto 0)
);
end pulse;

architecture rtl of pulse is

-- The pulse queue; keeps track of the timestamps of incoming pulses
component pulse_queue
port (
    clk                 : in std_logic;
    srst                : in std_logic;
    din                 : in std_logic_vector(48 DOWNTO 0);
    wr_en               : in std_logic;
    rd_en               : in std_logic;
    dout                : out std_logic_vector(48 DOWNTO 0);
    full                : out std_logic;
    empty               : out std_logic;
    data_count          : out std_logic_vector(10 downto 0)
);
end component;

-- Variable declarations

-- Attached to architecture inputs

signal DELAY            : std_logic_vector(47 downto 0);
signal DELAY_wstb       : std_logic;
signal STEP             : std_logic_vector(47 downto 0);
signal STEP_wstb        : std_logic;
signal WIDTH            : std_logic_vector(47 downto 0);
signal WIDTH_wstb       : std_logic;


-- Constants

constant c_number_zero          : std_logic_vector(1 downto 0) := "00";
constant c_number_one           : std_logic_vector(1 downto 0) := "01";
constant c_number_two           : std_logic_vector(1 downto 0) := "10";

constant c_timestamp_max        : unsigned(47 downto 0) := (others => '1');
constant c_timestamp_min        : unsigned(47 downto 0) := (others => '0');


-- Standard logic signals

signal enable_i_prev            : std_logic := '0';

signal fancy_delay_line_started : std_logic := '0';
signal first_pulse              : std_logic := '0';

signal got_first_pulse          : std_logic := '0';
signal got_pulse_program        : std_logic := '0';

signal had_falling_trigger      : std_logic := '0';
signal had_rising_trigger       : std_logic := '0';
signal had_trigger              : std_logic := '0';

signal pulse                    : std_logic := '0';
signal pulse_queued_empty       : std_logic := '0';
signal pulse_queued_full        : std_logic := '0';
signal pulse_queued_rstb        : std_logic := '0';
signal pulse_queued_wstb        : std_logic := '0';
signal pulse_value              : std_logic := '0';

signal queue_has_been_empty     : std_logic := '0';
signal queue_pulse_value        : std_logic := '0';

signal reset                    : std_logic := '0';

signal start_delay_countdown    : std_logic := '0';
signal signal_val               : std_logic := '0';
signal trig_fall_prev           : std_logic := '0';
signal trig_i_prev              : std_logic := '0';
signal trig_rise_prev           : std_logic := '0';
signal trig_same_prev           : std_logic := '0';

signal trig_fall                : std_logic := '0';
signal trig_rise                : std_logic := '0';
signal trig_same                : std_logic := '0';

signal value                    : std_logic := '0';

signal waiting_for_delay        : std_logic := '1';


-- Standard logic vector signals

signal program_progress         : std_logic_vector(1 downto 0) := (others => '0');

signal pulse_queued_din         : std_logic_vector(48 downto 0);
signal pulse_queued_dout        : std_logic_vector(48 downto 0);
signal pulse_queued_data_count  : std_logic_vector(10 downto 0);


-- Unsigned integer signals

signal delay_i                  : unsigned(47 downto 0) := (others => '0');
signal delay_i_prev             : unsigned(47 downto 0) := (others => '1');
signal delay_remaining          : unsigned(47 downto 0) := (others => '0');

signal edges_remaining          : unsigned(31 downto 0) := (others => '0');

signal gap_i                    : unsigned(47 downto 0) := (others => '0');
signal gap_i_prev               : unsigned(47 downto 0) := (others => '1');

signal missed_pulses            : unsigned(31 downto 0) := (others => '0');

signal pulses_i                 : unsigned(31 downto 0) := (others => '0');
signal pulse_gap                : unsigned(47 downto 0) := (others => '0');
signal pulse_ts                 : unsigned(47 downto 0) := (others => '0');
signal pulse_width              : unsigned(47 downto 0) := (others => '0');

signal queued_din               : unsigned(47 downto 0) := (others => '0');
signal queue_pulse_ts           : unsigned(47 downto 0) := (others => '0');

signal step_i                   : unsigned(47 downto 0) := (others => '0');
signal step_i_prev              : unsigned(47 downto 0) := (others => '1');
signal signal_ts                : unsigned(47 downto 0) := (others => '0');

signal timestamp                : unsigned(47 downto 0) := (others => '0');
signal timestamp_fall           : unsigned(47 downto 0) := (others => '0');
signal timestamp_prev           : unsigned(47 downto 0) := (others => '1');
signal timestamp_rise           : unsigned(47 downto 0) := (others => '0');

signal width_i                  : unsigned(47 downto 0) := (others => '0');
signal width_i_prev             : unsigned(47 downto 0) := (others => '1');

begin

-- The pulse queue; keeps track of the timestamps of incoming pulses, maps to component above, attached to this architecture
pulse_queue_inst : pulse_queue
port map (
    clk         => clk_i,
    srst        => reset,
    din         => pulse_queued_din,
    wr_en       => pulse_queued_wstb,
    rd_en       => pulse_queued_rstb,
    dout        => pulse_queued_dout,
    full        => pulse_queued_full,
    empty       => pulse_queued_empty,
    data_count  => pulse_queued_data_count
);

-- Code that runs outside of a process architecture (i.e. not executed in sequence, all executed in parallel)

-- Bits relating to the FIFO queue

queue_pulse_ts <= unsigned(pulse_queued_dout(47 downto 0));
queue_pulse_value <= pulse_queued_dout(48);


-- Other output assignments
DROPPED <= std_logic_vector(missed_pulses);
QUEUED <= ZEROS(32-pulse_queued_data_count'length) &  pulse_queued_data_count;


-- Bits relating to timings

-- Take 48-bit time as combination of two for:
-- 1) The delay width
DELAY_WSTB <= DELAY_L_WSTB or DELAY_H_WSTB;
DELAY(31 downto 0) <= DELAY_L;
DELAY(47 downto 32) <= DELAY_H(15 downto 0);

-- 2) The pulse width
WIDTH_WSTB <= WIDTH_L_WSTB or WIDTH_H_WSTB;
WIDTH(31 downto 0) <= WIDTH_L;
WIDTH(47 downto 32) <= WIDTH_H(15 downto 0);

-- 3) The overall step width
STEP_WSTB <= STEP_L_WSTB or STEP_H_WSTB;
STEP(31 downto 0) <= STEP_L;
STEP(47 downto 32) <= STEP_H(15 downto 0);


-- For those not requiring mathematics

-- If 0 < DELAY < 5, it should be set to 5
delay_i <=  (unsigned(DELAY) - 1) when (unsigned(DELAY) > 5) else
            (2 => '1', others => '0');

-- Make sure that if we recieve a pulse and the PULSE variable is accidentally set to zero we don't punish a hapless user
pulses_i <= unsigned(PULSES) when (unsigned(PULSES) /= 0) else
            (0 => '1', others => '0');

-- Set an internal width value
width_i <=  unsigned(WIDTH);


-- For those requiring mathematics

-- Calculate the minimum gap given all the other parameters
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        gap_i <= (others => '0');
        gap_i_prev <= (others => '1');
    elsif (rising_edge(clk_i) and enable_i = '1') then
        gap_i_prev <= gap_i;

        if (width_i /= width_i_prev or step_i /= step_i_prev) then
            if ((signed(step_i) - signed(width_i)) > 1) then
                gap_i <= step_i - width_i;
            else
                gap_i <= (0 => '1', others => '0');
            end if;
        end if;
    end if;
end process;


-- Calculate the minimum step given all the other parameters
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        step_i <= (others => '0');
        step_i_prev <= (others => '1');
    elsif (rising_edge(clk_i) and enable_i = '1') then
        step_i_prev <= step_i;

        if (width_i /= width_i_prev) then
            if (unsigned(STEP) > width_i) then
                step_i <= unsigned(STEP);
            else
                step_i <= unsigned(STEP) + width_i + 1;
            end if;
        end if;
    end if;
end process;


-- Code that runs inside process structures (i.e. code that runs in sequence with the blocks running in parallel)

-- Free running global timestamp counter
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        timestamp <= (others => '0');
    elsif (rising_edge(clk_i) and enable_i = '1') then
        timestamp <= timestamp + 1;
    end if;
end process;


-- Free running edge watcher
process(clk_i, trig_i)
begin
    if (rising_edge(clk_i)) then
        trig_fall <= '0';
        trig_rise <= '0';
        trig_same <= '1';
    elsif (falling_edge(trig_i)) then
        trig_fall <= '1';
        trig_same <= '0';
    elsif (rising_edge(trig_i)) then
        trig_rise <= '1';
        trig_same <= '0';
    end if;
end process;


-- Free running delay countdown block
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        delay_remaining <= (others => '0');
    elsif (rising_edge(clk_i) and enable_i = '1') then
        if (delay_remaining /= 0) then
            delay_remaining <= delay_remaining - 1;
        elsif ((start_delay_countdown = '1') and (pulse_queued_empty = '1')) then
            delay_remaining <= delay_i - 2;
        end if;
    end if;
end process;


-- Variable storage for comparison next clock cycle
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        delay_i_prev      <= (others => '1');
        enable_i_prev     <= '0';
        step_i_prev       <= (others => '1');
        timestamp_prev    <= (others => '1');
        trig_i_prev       <= trig_i;
        trig_fall_prev    <= '0';
        trig_rise_prev    <= '0';
        trig_same_prev    <= '0';
        width_i_prev      <= (others => '1');
    elsif (rising_edge(clk_i) and enable_i = '1') then
        delay_i_prev      <= delay_i;
        enable_i_prev     <= enable_i;
        step_i_prev       <= step_i;
        timestamp_prev    <= timestamp;
        trig_fall_prev    <= trig_fall;
        trig_i_prev       <= trig_i;
        trig_rise_prev    <= trig_rise;
        trig_same_prev    <= trig_same;
        width_i_prev      <= width_i;
    end if;
end process;


-- Filling the queue
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
        -- In case of a reset we'll need to reset these values from this process
        fancy_delay_line_started <= '0';

        got_first_pulse <= '0';

        had_rising_trigger <= '0';
        had_falling_trigger <= '0';

        missed_pulses <= (others => '0');
        
        pulse_queued_din <= (others => '0');
        pulse_queued_wstb <= '0';
        
        start_delay_countdown <= '0';

        timestamp_rise <= (others => '0');
        timestamp_fall <= (others => '0');

        value <= '0';

    elsif (rising_edge(clk_i) and enable_i = '1') then
        -- Bits that need resetting every clock cycle
        pulse_queued_wstb <= '0';
        value <= '0';
        start_delay_countdown <= '0';

        if (trig_rise = '1') then
            timestamp_rise <= timestamp;

        elsif (trig_fall = '1') then
            timestamp_fall <= timestamp;

        end if;

        if (waiting_for_delay = '0') then
            had_falling_trigger <= '0';
            had_rising_trigger <= '0';
        end if;

        -- If check to make sure that we should be storing this event at all
        if (trig_same /= '1') then
            -- First up, event rejection criteria:
            -- 1)   Queue full condition flags an error, and ticks missing pulse counter
            -- 2)   Pulse period must obey Xilinx FIFO IP latency following the first pulse
            -- 3)   Can't accept more pulses if we're processing them already
            if (fancy_delay_line_started = '0' and (pulse_queued_full = '1' or waiting_for_delay = '0' or edges_remaining /= 0)) then
                if(((TRIG_EDGE(1 downto 0) = c_number_zero) and (trig_rise = '1')) or
                   ((TRIG_EDGE(1 downto 0) = c_number_one) and (trig_fall = '1')) or
                    (TRIG_EDGE(1 downto 0) = c_number_two)) then
                        missed_pulses <= missed_pulses + 1;
                end if;

            -- Next, if we have a width (i.e. no timestamp maths required)
            elsif (width_i /= 0) then
                if(((TRIG_EDGE(1 downto 0) = c_number_zero) and (trig_rise = '1')) or
                   ((TRIG_EDGE(1 downto 0) = c_number_one) and (trig_fall = '1')) or
                    (TRIG_EDGE(1 downto 0) = c_number_two)) then
                        pulse_queued_din <= '1' & std_logic_vector(width_i);
                        pulse_queued_wstb <= '1';

                        start_delay_countdown <= '1';
                end if;

            -- If we have a step but no width
            elsif (width_i = 0 and unsigned(STEP) /= 0) then
                if (TRIG_EDGE(1 downto 0) = c_number_zero) then
                    if (trig_rise = '1' and had_rising_trigger = '0') then
                        had_rising_trigger <= '1';
                    elsif (trig_fall = '1' and had_rising_trigger = '1') then
                        had_rising_trigger <= '0';

                        if (timestamp_fall - timestamp_rise > 2) then
                            pulse_queued_din <= '0' & std_logic_vector(timestamp - timestamp_rise);
                        else
                            pulse_queued_din <= '0' & std_logic_vector((timestamp_prev - timestamp) + 1);
                        end if;

                        pulse_queued_wstb <= '1';
                        start_delay_countdown <= '1';
                    end if;
                end if;

                if (TRIG_EDGE(1 downto 0) = c_number_one) then
                    if (trig_fall = '1' and had_falling_trigger = '0') then
                        had_rising_trigger <= '1';
                    elsif (trig_rise = '1' and had_falling_trigger = '1') then
                        had_falling_trigger <= '0';

                        if (timestamp_rise - timestamp_fall > 2) then
                            pulse_queued_din <= '0' & std_logic_vector(timestamp - timestamp_fall);
                        else
                            pulse_queued_din <= '0' & std_logic_vector((timestamp_prev - timestamp) + 1);
                        end if;

                        pulse_queued_wstb <= '1';
                        start_delay_countdown <= '1';
                    end if;
                end if;

            -- If we have no step and no width
            elsif ((width_i = 0) and (unsigned(STEP) = 0)) then
                if (fancy_delay_line_started = '0') then
                    start_delay_countdown <= '1';
                    fancy_delay_line_started <= '1';
                end if;

                if (trig_rise = '1') then
                    pulse_queued_din <= '1' & std_logic_vector(timestamp + delay_i);
                    pulse_queued_wstb <= '1';
                elsif (trig_fall = '1') then
                    pulse_queued_din <= '0' & std_logic_vector(timestamp + delay_i);
                    pulse_queued_wstb <= '1';
                end if;
            end if;
        end if;
    end if;
end process;


-- Process to pass edges
process(clk_i, enable_i)
begin
    if (rising_edge(enable_i) or reset = '1') then
            edges_remaining <= (others => '0');
            
            pulse <= '0';
            pulse_queued_rstb <= '0';
            pulse_ts <= (others => '0');
            pulse_width <= (others => '0');
            pulse_value <= '0';

            waiting_for_delay <= '1';

    elsif (rising_edge(clk_i) and enable_i = '1') then
        pulse_queued_rstb <= '0';

        if (fancy_delay_line_started = '0') then
            if (delay_remaining = 1) then
                waiting_for_delay <= '0';
                pulse_queued_rstb <= '1';
            else
                if (pulse_queued_empty = '1' and (timestamp >= pulse_ts)) then
                    waiting_for_delay <= '1';
                end if;
            end if;
        else
            if (delay_remaining = 1) then
                waiting_for_delay <= '0';
            elsif (delay_remaining = 2) then
                pulse_ts <= queue_pulse_ts;
                pulse_value <= queue_pulse_value;
            end if;
        end if;

        --- If we're running as a fancy delay line
        if ((width_i = 0) and (unsigned(STEP) = 0)) then
            if (waiting_for_delay = '0' and timestamp = pulse_ts) then
                out_o <= pulse_value;
            end if;

            if (timestamp = (queue_pulse_ts - 2)) then
                pulse_queued_rstb <= '1';
                pulse_ts <= queue_pulse_ts;
                pulse_value <= queue_pulse_value;
            end if;
           
        --- Otherwise let's process some pulses
        else
            if (edges_remaining = 0) then
                if (waiting_for_delay = '0' and (timestamp >= pulse_ts)) then
                    if (width_i = 0 and unsigned(STEP) /= 0) then
                        if ((signed(step_i) - signed(queue_pulse_ts)) > 1) then
                            pulse_gap <= step_i - queue_pulse_ts;
                        else
                            pulse_gap <= (1 => '1', others => '0');
                        end if;

                        pulse_width <= queue_pulse_ts;
                    else
                        pulse_gap <= gap_i;
                        pulse_width <= queue_pulse_ts;
                    end if;

                    edges_remaining <= unsigned(pulses_i) + unsigned(pulses_i) - 1;
                    pulse_ts <= timestamp + queue_pulse_ts;
                    pulse <= '1';
                    out_o <= '1';
                end if;
            else
                if (timestamp = pulse_ts) then
                    if (unsigned(edges_remaining mod 2) = 0) then
                        edges_remaining <= edges_remaining - 1;
                        pulse_ts <= timestamp + pulse_width;
                        pulse <= not pulse;
                        out_o <= pulse;
                    else
                        edges_remaining <= edges_remaining - 1;
                        pulse_ts <= timestamp + pulse_gap;
                        pulse <= not pulse;
                        out_o <= pulse;
                    end if;

                    if (edges_remaining = 1) then
                        pulse_queued_rstb <= '1';
                    end if;
                end if;
            end if;
        end if;
    elsif (rising_edge(clk_i) and enable_i = '0') then
        out_o <= '0';
    end if;
end process;

end rtl;