--------------------------------------------------------------------------------
--  File:       pcap_dma.vhd
--  Desc:       Position capture module
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.support.all;

entity pcap_dma is
generic (
    AXI_BURST_LEN       : natural := 16;        -- AXI3 standard
    AXI_ADDR_WIDTH      : natural := 32;
    AXI_DATA_WIDTH      : natural := 32
);
port (
    -- Clock and Reset
    clk_i               : in  std_logic;

    -- Block Input and Outputs
    pcap_dat_i          : in  std_logic_vector(31 downto 0);
    pcap_wstb_i         : in  std_logic;
    pcap_done_i         : in  std_logic;
    pcap_status_i       : in  std_logic_vector(2 downto 0);
    dma_error_o         : out std_logic;
    irq_o               : out std_logic;

    -- Block Registers
    DMA_RESET           : in  std_logic;
    DMA_INIT            : in  std_logic;
    DMA_ADDR            : in  std_logic_vector(31 downto 0);
    DMA_ADDR_WSTB       : in  std_logic;
    TIMEOUT             : in  std_logic_vector(31 downto 0);
    TIMEOUT_WSTB        : in  std_logic;
    IRQ_STATUS          : out std_logic_vector(31 downto 0);
    BLOCK_SIZE          : in  std_logic_vector(31 downto 0);

    -- AXI3 HP Bus Write Only Interface
    m_axi_awready       : in  std_logic;
    m_axi_awregion      : out std_logic_vector(3 downto 0);
    m_axi_awaddr        : out std_logic_vector(AXI_ADDR_WIDTH-1 downto 0);
    m_axi_awvalid       : out std_logic;
    m_axi_awburst       : out std_logic_vector(1 downto 0);
    m_axi_awcache       : out std_logic_vector(3 downto 0);
    m_axi_awid          : out std_logic_vector(5 downto 0);
    m_axi_awlen         : out std_logic_vector(3 downto 0);
    m_axi_awlock        : out std_logic_vector(1 downto 0);
    m_axi_awprot        : out std_logic_vector(2 downto 0);
    m_axi_awqos         : out std_logic_vector(3 downto 0);
    m_axi_awsize        : out std_logic_vector(2 downto 0);
    m_axi_bid           : in  std_logic_vector(5 downto 0);
    m_axi_bready        : out std_logic;
    m_axi_bresp         : in  std_logic_vector(1 downto 0);
    m_axi_bvalid        : in  std_logic;
    m_axi_wready        : in  std_logic;
    m_axi_wdata         : out std_logic_vector(AXI_DATA_WIDTH-1 downto 0);
    m_axi_wvalid        : out std_logic;
    m_axi_wlast         : out std_logic;
    m_axi_wstrb         : out std_logic_vector(AXI_DATA_WIDTH/8-1 downto 0)
);
end pcap_dma;

architecture rtl of pcap_dma is

-- Bit-width required to represent maximum burst length (5)
constant AXI_BURST_WIDTH    : integer := LOG2(AXI_BURST_LEN) + 1;
-- Number of byte per AXI burst
constant BURST_LEN          : integer := AXI_BURST_LEN * AXI_ADDR_WIDTH/8;

component fifo_1K32_ft
port (
    clk                 : in std_logic;
    srst                : in std_logic;
    din                 : in std_logic_vector(31 DOWNTO 0);
    wr_en               : in std_logic;
    rd_en               : in std_logic;
    dout                : out std_logic_vector(31 DOWNTO 0);
    full                : out std_logic;
    empty               : out std_logic;
    data_count          : out std_logic_vector(10 downto 0)
);
end component;

signal BLOCK_TLP_SIZE       : unsigned(31 downto 0);
signal M_AXI_BURST_LEN      : std_logic_vector(AXI_BURST_WIDTH-1 downto 0);
signal reset                : std_logic;

type pcap_fsm_t is (INIT, ACTV, DO_DMA, IS_FINISHED, IRQ, COMPLETED);
signal pcap_fsm             : pcap_fsm_t;

signal IRQ_STATUS_T         : std_logic_vector(31 downto 0);
signal first_data           : std_logic;
signal timeout_counter      : unsigned(31 downto 0);
signal pcap_timeout         : std_logic;
signal pcap_timeout_latch   : std_logic;

signal dma_start            : std_logic;
signal dma_done             : std_logic;
signal dma_irq              : std_logic;
signal dma_error            : std_logic;
signal tlp_count            : unsigned(31 downto 0);
signal last_tlp             : std_logic;
signal axi_awaddr_val       : unsigned(31 downto 0);
signal axi_wdata_val        : std_logic_vector(AXI_DATA_WIDTH-1 downto 0);
signal next_dmaaddr_valid   : std_logic;
signal switch_block         : std_logic;
signal pcap_wstb            : std_logic;
signal writing_sample       : std_logic;

signal fifo_data_count      : std_logic_vector(10 downto 0);
signal fifo_count           : unsigned(10 downto 0);
signal transfer_size        : unsigned(AXI_BURST_WIDTH-1 downto 0);
signal fifo_rd_en           : std_logic;
signal fifo_dout            : std_logic_vector(AXI_DATA_WIDTH-1 downto 0);
signal fifo_full            : std_logic;

signal irq_flags            : std_logic_vector(7 downto 0);
signal sample_count         : unsigned(23 downto 0);
signal pcap_completed       : std_logic;

signal pcap_error           : std_logic;

begin

-- Assign outputs.
irq_o <= dma_irq;

-- DMA engine reset
reset <= DMA_RESET;

-- DMA error occurs when fifo is full or AXI transaction error
-- This flag is used to abort ongoing pcap operation along with other flags
dma_error_o <= fifo_full or dma_error;

-- TLP_COUNT = BLOCK_SIZE/BURST_LEN
BLOCK_TLP_SIZE <= to_unsigned((to_integer(unsigned(BLOCK_SIZE)) / BURST_LEN),32);

-- Pcap status information
--  pcap_status_i[0] : user disarmed
--  pcap_status_i[1] : framing error
--  pcap_status_i[2] : dma error
pcap_error <= pcap_status_i(2) or pcap_status_i(1);

--
-- 32bit FIFO with 1K sample depth
--
dma_fifo_inst : fifo_1K32_ft
port map (
    srst            => reset,
    clk             => clk_i,
    din             => pcap_dat_i,
    wr_en           => pcap_wstb_i,
    rd_en           => fifo_rd_en,
    dout            => fifo_dout,
    full            => fifo_full,
    empty           => open,
    data_count      => fifo_data_count
);

fifo_count <= unsigned(fifo_data_count);
transfer_size <= to_unsigned(AXI_BURST_LEN, AXI_BURST_WIDTH)
                   when (fifo_count > AXI_BURST_LEN) else
                     unsigned(fifo_data_count(AXI_BURST_WIDTH-1 downto 0));

--------------------------------------------------------------------------
-- PCAP Main State Machine
--
-- Order of actions are as follows for Initialisation, and IRQ handling
--
--
--                INIT         IRQ
--              ----------- ----------
-- RESET       | 1.w       |          |
-- ENABLE      | 3.w       |          |
-- ADDR        | 2.w, 4.w  | 3.w      |
-- IRQ_FLAGS   |           | 1.r      |
-- SMPL_COUNT  |           | 2.r      |
--

-- DMA_ADDR_WSTB strobe is used as a handshake between PS and
-- PL logic. If PS can not keep up with the DMA rate by setting
-- next DMA address on irq, DMA will be aborted.
--------------------------------------------------------------------------
process(clk_i) begin
    if rising_edge(clk_i) then
        if (reset = '1') then
            next_dmaaddr_valid <= '0';
        else
            if (DMA_ADDR_WSTB = '1') then
                next_dmaaddr_valid <= '1';
            -- Clear flag on every IRQ
            elsif (pcap_fsm = IRQ) then
                next_dmaaddr_valid <= '0';
            end if;
        end if;
    end if;
end process;

--------------------------------------------------------------------------
-- Timeout Counter is used to issue an interrupt @ TIMEOUT rate for very
-- slow acquisition.
-- TIMEOUT = 0 disables the counter, otherwise counter is active only in
-- ACTV state.
--------------------------------------------------------------------------
writing_sample <= pcap_wstb_i or pcap_wstb;

process(clk_i) begin
    if rising_edge(clk_i) then
        if (reset = '1') then
            first_data <= '0';
            pcap_timeout <= '0';
            timeout_counter <= (others => '0');
            pcap_timeout_latch <= '0';
            pcap_wstb <= '0';
        else
            pcap_wstb <= pcap_wstb_i;
            -- Wait until first data received to prevent empty timeout IRQs
            if (pcap_fsm = INIT) then
                first_data <= '0';
            elsif (pcap_wstb_i = '1') then
                first_data <= '1';
            end if;

            -- Reset timeout on start-up and interrupts, and synchronise to
            -- first incoming sample
            if (pcap_fsm = INIT or pcap_fsm = IRQ or first_data = '0') then
                pcap_timeout <= '0';
                timeout_counter <= (others => '0');
            else
                timeout_counter <= timeout_counter + 1;
                if (unsigned(TIMEOUT) = 0) then
                    pcap_timeout <= '0';
                elsif (timeout_counter = unsigned(TIMEOUT) - 1) then
                    pcap_timeout <= '1';
                end if;
            end if;

            -- Latch timeout flag for interrupt status
            if (pcap_fsm = ACTV and pcap_timeout = '1') then
                pcap_timeout_latch <= '1';
            elsif (pcap_fsm = IRQ) then
                pcap_timeout_latch <= '0';
            end if;
        end if;
    end if;
end process;

process(clk_i) begin
    if rising_edge(clk_i) then
        if (reset = '1') then
            pcap_completed <= '0';
        elsif (pcap_done_i = '1') then
            pcap_completed <= '1';
        end if;
    end if;
end process;

--------------------------------------------------------------------------
-- Main State Machine
--
-- tlp_count       : # of TLPs DMAed per IRQ.
-- sample_count    : # of samples (DWORDs) DMAed per IRQ.
-- M_AXI_BURST_LEN : # of beats in individual AXI3 write.
--------------------------------------------------------------------------

switch_block <= '1' when (tlp_count = BLOCK_TLP_SIZE) else  '0';

PCAP_STATE : process(clk_i)
begin
if rising_edge(clk_i) then
    if (reset = '1') then
        pcap_fsm <= INIT;
        IRQ_STATUS_T <= (others => '0');
        dma_irq <= '0';
        last_tlp <= '0';
        dma_start <= '0';
        axi_awaddr_val <= (others => '0');
        M_AXI_BURST_LEN <= (others => '0');
        tlp_count <= (others => '0');
        sample_count <= (others => '0');
    else
        case pcap_fsm is
            -- Wait Initialistion by kernel driver
            when INIT =>
                axi_awaddr_val <= unsigned(DMA_ADDR);
                if (DMA_INIT = '1') then
                    pcap_fsm <= ACTV;
                end if;

            -- Wait until FIFO has enough data worth for a AXI burst
            -- (AXI_BURST_LEN beats).
            when ACTV =>
                dma_irq <= '0';
                -- An unrecoverable error occured, no need to continue 
                -- finishing off the buffer
                if (pcap_completed = '1' and pcap_error = '1') then
                    last_tlp <= '1';
                    pcap_fsm <= IRQ;
                -- Timeout occured, transfer all data in the buffer before
                -- raising IRQ.
                elsif (pcap_timeout = '1' and writing_sample = '0') then
                    if (fifo_count = 0) then
                        pcap_fsm <= IRQ;
                    else
                        dma_start <= '1';
                        sample_count <= sample_count + transfer_size;
                        M_AXI_BURST_LEN <= std_logic_vector(transfer_size);
                        pcap_fsm <= DO_DMA;
                    end if;
                -- At least 1 TLP in available the queue
                elsif (fifo_count > AXI_BURST_LEN and writing_sample = '0') then
                    dma_start <= '1';
                    sample_count <= sample_count + transfer_size;
                    M_AXI_BURST_LEN <= std_logic_vector(transfer_size);
                    pcap_fsm <= DO_DMA;
                -- Position compare completed
                elsif (pcap_completed = '1' and writing_sample = '0') then
                    last_tlp <= '1';
                    if (fifo_count = 0) then
                        pcap_fsm <= IRQ;
                    else
                        dma_start <= '1';
                        sample_count <= sample_count + transfer_size;
                        M_AXI_BURST_LEN <= std_logic_vector(transfer_size);
                        pcap_fsm <= DO_DMA;
                    end if;
                end if;

            -- Waits until DMA Engine completes. Also keeps tracks of TLPs
            -- for Buffer switching.
            when DO_DMA =>
                dma_start <= '0';
                if (dma_done = '1') then
                    tlp_count <= tlp_count + 1;
                    pcap_fsm <= IS_FINISHED;
                end if;

            -- Decide what to do next.
            when IS_FINISHED =>
                -- Timeout or buffer full, should switch buffers
                if(pcap_timeout_latch = '1' or switch_block = '1') then
                    pcap_fsm <= IRQ;
                -- Block buffer is not consumed and Pcap is still active
                else
                    pcap_fsm <= ACTV;
                    axi_awaddr_val <= axi_awaddr_val + BURST_LEN;
                end if;

            -- Set IRQ flag, and either continue or stop operation
            when IRQ =>
                -- Raise the interrupt to PS
                dma_irq <= '1';

                -- Switch to next given buffer and reset sample counter
                axi_awaddr_val <= unsigned(DMA_ADDR);
                sample_count <= (others => '0');
                tlp_count <= (others => '0');

                -- Latch IRQ status flags
                IRQ_STATUS_T(31 downto 8) <= std_logic_vector(sample_count);
                IRQ_STATUS_T(7 downto 0) <= irq_flags;

                -- Next state
                if (last_tlp = '1' or next_dmaaddr_valid = '0') then
                    pcap_fsm <= COMPLETED;
                else
                    pcap_fsm <= ACTV;
                end if;

            -- Either End-Of-Experiment or Abort-on-Error happened.
            -- Requires full DMA reset-init cycle.
            when COMPLETED =>
                dma_irq <= '0';

            when others =>

        end case;
    end if;
end if;
end process;

--------------------------------------------------------------------------
-- Keep track of system status
--------------------------------------------------------------------------
-- PCAP completed or next buffer is not ready on interrupt
irq_flags(0) <= last_tlp or not next_dmaaddr_valid;
-- Completion reason (0 = Successful)
irq_flags(3 downto 1) <= pcap_status_i;
irq_flags(4) <= not next_dmaaddr_valid;
irq_flags(5) <= pcap_timeout_latch;
irq_flags(6) <= switch_block;
irq_flags(7) <= '0';

--
-- AXI DMA Master Engine
--
WORD_SWAP_32 : if (AXI_DATA_WIDTH = 32) generate
    axi_wdata_val(31 downto 0) <= fifo_dout(31 downto 0);
end generate;

WORD_SWAP_64 : if (AXI_DATA_WIDTH = 64) generate
    axi_wdata_val(63 downto 32) <= fifo_dout(31 downto 0);
    axi_wdata_val(31 downto 0) <= fifo_dout(63 downto 32);
end generate;

dma_write_master : entity work.axi_write_master
generic map (
    AXI_BURST_WIDTH     => AXI_BURST_WIDTH,
    AXI_ADDR_WIDTH      => AXI_ADDR_WIDTH,
    AXI_DATA_WIDTH      => AXI_DATA_WIDTH
)
port map (
    clk_i               => clk_i,
    reset_i             => reset,

    m_axi_burst_len     => M_AXI_BURST_LEN,

    m_axi_awready       => m_axi_awready,
    m_axi_awregion      => m_axi_awregion,
    m_axi_awaddr        => m_axi_awaddr,
    m_axi_awvalid       => m_axi_awvalid,
    m_axi_awburst       => m_axi_awburst,
    m_axi_awcache       => m_axi_awcache,
    m_axi_awid          => m_axi_awid,
    m_axi_awlen         => m_axi_awlen,
    m_axi_awlock        => m_axi_awlock,
    m_axi_awprot        => m_axi_awprot,
    m_axi_awqos         => m_axi_awqos,
    m_axi_awsize        => m_axi_awsize,
    m_axi_bid           => m_axi_bid,
    m_axi_bready        => m_axi_bready,
    m_axi_bresp         => m_axi_bresp,
    m_axi_bvalid        => m_axi_bvalid,
    m_axi_wready        => m_axi_wready,
    m_axi_wdata         => m_axi_wdata,
    m_axi_wvalid        => m_axi_wvalid,
    m_axi_wlast         => m_axi_wlast,
    m_axi_wstrb         => m_axi_wstrb,

    dma_addr            => std_logic_vector(axi_awaddr_val),
    dma_data            => axi_wdata_val,
    dma_read            => fifo_rd_en,
    dma_start           => dma_start,
    dma_done            => dma_done,
    dma_error           => dma_error
);

IRQ_STATUS <= IRQ_STATUS_T;

end rtl;

