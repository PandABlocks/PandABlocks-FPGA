library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.top_defines.all;
use work.support.all;

package register_map is

constant OUTTTL0_VAL    : std_logic_vector := TO_STD_VECTOR(0, MEM_AW);
constant OUTTTL1_VAL    : std_logic_vector := TO_STD_VECTOR(1, MEM_AW);
constant OUTTTL2_VAL    : std_logic_vector := TO_STD_VECTOR(2, MEM_AW);
constant OUTTTL3_VAL    : std_logic_vector := TO_STD_VECTOR(3, MEM_AW);
constant OUTTTL4_VAL    : std_logic_vector := TO_STD_VECTOR(4, MEM_AW);
constant OUTTTL5_VAL    : std_logic_vector := TO_STD_VECTOR(5, MEM_AW);
constant OUTTTL6_VAL    : std_logic_vector := TO_STD_VECTOR(6, MEM_AW);
constant OUTTTL7_VAL    : std_logic_vector := TO_STD_VECTOR(7, MEM_AW);
constant OUTLVDS0_VAL   : std_logic_vector := TO_STD_VECTOR(8, MEM_AW);
constant OUTLVDS1_VAL   : std_logic_vector := TO_STD_VECTOR(9, MEM_AW);



end register_map;


package body register_map is


end register_map;

