--------------------------------------------------------------------------------
--  File:       panda_pgen.vhd
--  Desc:       5-Input LUT.
--
--  Author:     Isa S. Uzun (isa.uzun@diamond.ac.uk)
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity panda_pgen is
generic (
    AXI_BURST_LEN       : integer := 256;
    DW                  : natural := 32
);
port (
    -- Clock and Reset
    clk_i               : in  std_logic;
    reset_i             : in  std_logic;
    -- Block Input and Outputs
    enable_i            : in  std_logic;
    trig_i              : in  std_logic;
    out_o               : out std_logic_vector(31 downto 0);
    -- Block Parameters
    CYCLES              : in  std_logic_vector(31 downto 0);
    TABLE_ADDR          : in  std_logic_vector(31 downto 0);
    TABLE_LENGTH        : in  std_logic_vector(31 downto 0);
    TABLE_LENGTH_WSTB   : in  std_logic;
    -- DMA Engine Interface
    dma_req_o           : out std_logic;
    dma_ack_i           : in  std_logic;
    dma_done_i          : in  std_logic;
    dma_addr_o          : out std_logic_vector(31 downto 0);
    dma_len_o           : out std_logic_vector(7 downto 0);
    dma_data_i          : in  std_logic_vector(DW-1 downto 0);
    dma_valid_i         : in  std_logic
);
end panda_pgen;

architecture rtl of panda_pgen is

component pgen_dma_fifo
port (
    clk                 : in std_logic;
    rst                 : in std_logic;
    din                 : in std_logic_vector(31 DOWNTO 0);
    wr_en               : in std_logic;
    rd_en               : in std_logic;
    dout                : out std_logic_vector(31 DOWNTO 0);
    full                : out std_logic;
    empty               : out std_logic;
    data_count          : out std_logic_vector(10 downto 0)
);
end component;

type state_t is (IDLE, WAIT_FIFO, DMA_REQ, DMA_READ, IS_FINISHED, FINISHED);
signal pgen_fsm         : state_t;

signal reset            : std_logic;
signal TABLE_WORDS      : unsigned(31 downto 0);

signal table_cycle      : unsigned(31 downto 0);
signal table_ready      : std_logic;

signal fifo_reset       : std_logic;
signal fifo_rd_en       : std_logic;
signal fifo_dout        : std_logic_vector(DW-1 downto 0);
signal fifo_count       : integer range 0 to 2047;
signal fifo_full        : std_logic;
signal fifo_data_count  : std_logic_vector(10 downto 0);
signal fifo_available   : std_logic;

signal trig             : std_logic;
signal enable           : std_logic;
signal trig_pulse       : std_logic;
signal enable_fall      : std_logic;

signal count            : unsigned(31 downto 0);
signal dma_len          : unsigned(8 downto 0);
signal dma_addr         : unsigned(31 downto 0);

begin

-- Assign outputs
dma_len_o <= std_logic_vector(dma_len(7 downto 0));
dma_addr_o <= std_logic_vector(dma_addr);
out_o <= fifo_dout;

-- Reset for state machine
reset <= reset_i or not table_ready or enable_fall;

--
-- 32bit FIFO with 1K sample depth
--
dma_fifo_inst : pgen_dma_fifo
port map (
    rst             => fifo_reset,
    clk             => clk_i,
    din             => dma_data_i,
    wr_en           => dma_valid_i,
    rd_en           => fifo_rd_en,
    dout            => fifo_dout,
    full            => fifo_full,
    empty           => open,
    data_count      => fifo_data_count
);

fifo_reset <= reset;
fifo_rd_en <= trig_pulse;
fifo_count <= to_integer(unsigned(fifo_data_count));
fifo_available <= '1' when (fifo_count < 768) else '0';

--
-- Input registers
--
process(clk_i) begin
    if rising_edge(clk_i) then
        trig <= trig_i;
        enable <= enable_i;
    end if;
end process;

-- Trigger pulse pops data from fifo and tick data counter when block
-- is enabled and table is ready.
trig_pulse <= (trig_i and not trig) and enable_i and table_ready;
enable_fall <= not enable_i and enable;

--
-- Table ready controls state machine reset. The table is un-validated once
-- LENGTH=0 written.
--
TABLE_WORDS <= unsigned(TABLE_LENGTH) srl 2;  -- Byte -> Dword

process(clk_i) begin
    if rising_edge(clk_i) then
        if (reset_i = '1') then
            table_ready <= '0';
        else
            if (TABLE_LENGTH_WSTB = '1') then
                if (TABLE_WORDS = 0) then
                    table_ready <= '0';
                elsif (TABLE_WORDS /= 0) then
                    table_ready <= '1';
                end if;
            end if;
        end if;
    end if;
end process;

process(clk_i) begin
    if rising_edge(clk_i) then
        if (reset = '1') then
            dma_req_o <= '0';
            count <= (others => '0');
            dma_addr <= (others => '0');
            dma_len <= (others => '0');
            table_cycle <= (others => '0');
            pgen_fsm <= IDLE;
        else
            case pgen_fsm is
                when IDLE =>
                    -- Wait following fifo reset by monitoring full flag.
                    if (fifo_full = '0') then
                        table_cycle <= table_cycle + 1;
                        count <= TABLE_WORDS;
                        dma_addr <= unsigned(TABLE_ADDR);
                        pgen_fsm <= WAIT_FIFO;
                    end if;

                -- Wait until enough space available in the fifo.
                when WAIT_FIFO =>
                    if (fifo_available = '1') then
                        dma_req_o <= '1';
                        pgen_fsm <= DMA_REQ;

                        -- Determine dma length in samples.
                        if (count < AXI_BURST_LEN) then
                            dma_len <= count(8 downto 0);
                        else
                            dma_len <= to_unsigned(AXI_BURST_LEN, dma_len'length);
                        end if;
                    end if;

                when DMA_REQ =>
                    if (dma_ack_i = '1') then
                        dma_req_o <= '0';
                        pgen_fsm <= DMA_READ;
                    end if;

                when DMA_READ =>
                    -- Wait until DMA completes, and keep track of total count.
                    if (dma_done_i = '1') then
                        count <= count - dma_len;
                        dma_addr <= dma_addr + dma_len * 4;
                        pgen_fsm <= IS_FINISHED;
                    end if;

                when IS_FINISHED =>
                    -- Is table finished?
                    if (count = 0) then
                        -- Are there more table cycles?
                        if (table_cycle = unsigned(CYCLES)) then
                            pgen_fsm <= FINISHED;
                        else
                            count <= TABLE_WORDS;
                            dma_addr <= unsigned(TABLE_ADDR);
                            pgen_fsm <= WAIT_FIFO;
                            table_cycle <= table_cycle + 1;
                        end if;
                    else
                        pgen_fsm <= WAIT_FIFO;
                    end if;

                -- Wait for re-enable to start over.
                when FINISHED =>
                    dma_req_o <= '0';
                    count <= (others => '0');
                    dma_addr <= (others => '0');
                    dma_len <= (others => '0');
            end case;
        end if;
    end if;
end process;

end rtl;

