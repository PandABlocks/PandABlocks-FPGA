library ieee;
use ieee.std_logic_1164.all;
package slow_version is
constant SLOW_FPGA_VERSION: std_logic_vector(31 downto 0)   := X"23021700";
end slow_version;
