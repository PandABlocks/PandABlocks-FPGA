`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rD+dVeClxa5UKiAeGPSos59e0yGruYVZi+W/E+0q3fZeAjTB+esh7TgdUdHfBjzrqSij4ITE13SB
S2JTA0+Lxw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gOFW7NYGrBefbvEmNP/RoKVgAM+JPbz39U+/GYb30Z575UtDQulr9SX4XJnY7uSV40YUJ2ArXd24
OY4Z5AB9fiMNGA76bpOHLvGgHnu6l/objBS/Wz5AG5Y605zXoFjje4C6kA6X3UqKBfHsY0jz0hsC
vz2foTkPJrLM12y3Edg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fLzV/2Lx//cfK0x/bUaUV2CBkd86pxFH92BuYuZcuFu1oHBj7L8oMae44nU6anOJ0bbfks8lhzQC
b8Cj35a+SBYIfMz+sN9vYNunT7rmzw/eE8HnmaJuglw7ycr07dmRuTnvJKlhMpMQtBeQIl8CHPnK
eBV7OPQuSxPWiDRYJx2Rj0mYaDEUCB/UHXHbdM1har3rDftLp4or1Gta45jMXe53D6DwgVHTmFQ0
QX4V5IcmNfof9+Pp6TeaA7jiYyecJUx8c5VkS+MsJvtyKpgT7BvlsO9oZknCfvRvQBu8sKk+Vsrc
XVF26jvVYm5WKyAgbsLkZIc7Sw8V1Z+tu2Cx9g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Hk0C5QdySjsdnqNSf/TQ0ywVrxMSePJS+YXzTTuNiNV3smgIh3MuTQCTxDwEtkQBwTirzdj0UAY6
UcL2Z+7AQAECIESNxFE9S7mQNtq+KnQMLsg+PkS6RgxdeGsVZ79GnzMmQZ5zFxMVyu4g4OgrrCNb
gvnN9Czy5GSbkjvKbHk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nkoloWRMWd2XlHh/zsh4/7c8WPJ2mRzQLi/+v3Fs1TviBbuQPYRFHjFiQZAFZg1bkP7UIGFs8fOT
K7j8xmPkWDnFlSLPFJ1VXXiwngN+K7IqRaqeJPl7mfp+Ll+BfRHfZ47EzOyQil9Wb2u+9lYytH2h
NT04IiYZ2Mpra6Mx/+uc0FwWwrOMXIjqneysNBX+iMgpzEl2h3LnGTr1JSMXjKmK/VoO5ZFfdFd/
XnppjEUCeylPd+dlYiGH/kbBASgoUXJ7mt2nQ9ThPtuojx/qVb52/sS6tCp/oCehxkf9cRKD8PA3
psxBGy4Qs2dEwMkU3RphG9PLPzc2nwbZUA5PTQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1459520)
`protect data_block
EUukn7t7KP/vTXvThjEUCK5/p7vo9htgmGCbpD3Ay2TwToCa1Qs8IuKSBgbgUxpXZKsQrKZZmF6U
m1GEJ5i0neG8hHLaZSQ8tPeHLdqFPU+6gBVUPRm6IoCiN6gf3COdtzmy79b6GcY6sZ4wpVoBwxdq
qKtK37USS1zK06olFLg12jC/DLQfaEoxDouegnt04RPdll1U70LM+lnsHCJA5zFyeUrS4+yTC8qK
0y/RcJ1tLKhYctOZmRWBuLlGN6UCQzcE7RtTqSs6RwZ8IHmSuEbcGJNdYKDIiABzPCbqXn2WkwRr
SO0gOTvL+rWV1gZ9KVoE/qmEAXCupXu6AZuAk3bE5i8LK460HS2PbzGhD2OvGl+Gckk98KMbH479
Pg80t+d/r+qrJ55CSbPX4pl0Z4kKydTBm93izQ+UJojalAPiSqIfpf16eOsPifeyyk1NDgSOxSVh
g1EfA6OB47bI8TOGf/GH/08szYODstNbANsC+V0Drix2QNPu4h6FpwTlbo8VRn7VJ7MlT990lTDn
6IuoYL0A8kwQgmBGn2FL42+0pZ/7INUZ7Q0lquoyo6CFe9WNgxtMQPRjnk2WekVf6sHlCY9nYI6d
AuVks0YqZdjKO/XXU4MYoak2X9bI4EWK4djBFY/UyCQrhsTIgPTJZl9GYUudZlKtGT/JVY3uR2o+
QIODfm5HGIKyTLc6Y1ktgcR3yr5YfmXccKtn4c1WEfVICTOoJb1GX6rmPhfzuZLt/Um5RgH7Nswn
NCUjKsDWqNs0ljiP3MR54SEzEB9t1KN7hjyk8aDyldxQs+KODLgKpz1bt0agSeEw/AXRgLyXJ2az
ZqG5cCtMoUS71qSABAktQEx/b+TWAyls0QD4tO29nBpclUzLs/uTmULOy039LJKrvzKz2yh97ogo
vjh90Ezps1wM9kkj6jd64/GMrpDe5PWD5yknIOg8fDmIROO8JLQte00a/F7NXeSlZQLn682JSf51
EPKa6DSuvfC6DJ/BeGxC56yJobPEaWFfVopnR7PkH2Bj4B9XtcKt2Wy21Jg2Wf4dQ6nH9HQ5+gKD
Bx7AfQ2HKymLIKw3NP/nlOlGaf8cKAubrr5Eq6Dcd6iVVFTiO8FNwDlGLo1Ec1i5eckswJqfb8fS
vP8dkx15S82gfYH/yd7H4riiO9Z+UlmmN4653MVcBprDsb0/Hq9QCgE30RmPsfb4LTjwcxRtfBdZ
qAbhNDM1KksHax5IO+9kBlo5yt0vtZjnhL1zdN+29NTvoVV57MrCEAwMxDLhXw8s9FviWz9yxDWp
fNmjKRX/feoMwKFfLN1Xg9A2kAJpmHpIB/C3pOdMvLV6EM5sT17pucop8651EMiyRG+aqOA1VjHv
6mnFf+RE2VJ+rUX6NVtFt87WckQMaApXO64GWhyHTce9rz5NR9SuXXkQBQovm1+RAbitT3fu8r/a
DfaD4lQ4TQg7JwS90KX1cuO6hXdlNwQ/GfRJODLcXX+aoKxq8+euy7nSFznTMJ2Iicvfem7TXSUp
j7TiTMLBb2YCOM5X05P9g7CsU0qfIsAbUaHAIDfUezyy4zmKuz/0IIGKWORofm51uWPXybmWK5gi
Ug+0NWP7Dg1fnI7gJTMvwHEgI6VbpMyvVLtlZsViz3ZC/yXCWBECU/M63ZAHklEnuA5rHpIqIyxx
Ub5M3T8hTV4KC6OJ84X3AfU7ZaQ40FYT3WvsKVct1yv/spm/3JJLPRq2wLyWlYtbIKu+7KdTA9v5
+/ifPXKeJ5Gvj67bJ8Tsav7TK7G32w4lvrP0psAO0Hikdp8ItNwABk8oj0gohcOE1+qhCURNMDH9
Cplr3BjwHoZ8bzrJnNcKsm6KSJjS0Ta50QB5T2iILyaNCOq+c6cfieYFtPNlFrARXv76Pa34ZfTf
DHP/A9dHKfz6RUbMzAteq3Y1kq65b+jzpq8Rw26Y++6wTMmq3xsgy+AhTBFmvisaYpMUcbypVUO1
vRwv8KGEiQ6INJqKOMuN8jLU20EmOEd2r5QWYG+2q9axkzE2p+nuDKp1VLnRg5/APjHOWOlpDsxI
JJ9h4UIz/Smpjg6fozr0w9wTIWggV6X3wM7C8WWcW44TEj9GSJq1OYhOkYX1W9ZwqiVLDPfVO2mp
7mI3qihTE9tOoexxcQVGW4HAqui7oQXDnbBQ9vqNoU7t5xYAQpdA2P4rvbtKfW6/kopnqivIpX0s
9UaMz9Y+eajMneiRPfFLXsXuYhsM+YEX+Ve0rzlfKQd9d4QrGRYuKulTwSYdtggaD0LQhjCs81S4
YkjDb+NuyoIDiAgU8eRqmLodmWFcu1Q0Qc834HHr4AXPSL3qTFeVphZJtxb07hLox1ZVR31PjnoI
rsP9+rNMpXNknXIZkVLcsX+d8aTlCrpn11lDTZIiZVR7aZEFvuplzATL9zZ6Ih7G2dMCJBNK8tTz
/xy+0MtTmMT2mXnUtLMJAVm0SEPAL9RwJ7PDuJxCn9F0+XPHxeJYN7gXW6cJPHTDJhvyuj/mzIkp
Eenkdqb47tcXfGwV8DuEpcdLiGkhKgh9vpHAo9mFksR5UhaQqxv53+5Km5aUPDoiDrWGCyCyfASw
D+NiMVKS5C4Zvto5UBJ2HsFZFjKj8IAfyIIRpWuuPAMNhgySkCy/UG+2PE0NN0Zf3enVv7O1Kyih
ik4KDTCZ0NXdAqZSueTGhi+PQ4aQKA4eJ8mrPBwXnQ/6GjvSDZAOxCOeXR/1H1YGKWd3Inpeoq79
GhBBxZzdUXt0qkQRWa4oQz6wGgk8YQ7Oo21nhMCcq94s08wb9Yp6GY8r2SlVomPwGMK28ApfBFcf
hjmxBv4ZuTdsECqQ0pTGcV5GLls/6fyxM7en2O11SYhCtNFwtspUANmIOmJB7HLCMVpxfZbP3nYC
SvpGfgzxIG9H6o/d8Oom8K7DqvwXl5aLSQ4jNTYBnKNI2DLkJ1T4V/We3KH/s4M/eSYBQ7hZTfvj
HysAVQSs/izIWEr51iOQEQngzetWpdkQvgMoLaefxutU6FWEHIt7c3Fd+RgzZQfPWsqBEDHilB5h
JBB1DUGW3FcUy18V4aG88L61G6nsfSi9a8e/nbfo2vLfBGeuPtexJqgmC6ZtxXOaUIdGKEpg9dDP
B98HoCZomw74TIgk7+pSVQAPi0VnePOKkkVZXbhEMtF/kpQvdNMTLF7XJ20KHMrSAjNsFPqtdM8X
rsvqhHvZ7uPzU5/GaVdKaGADDkILYzsPq1k5ImEjmHvLmcbvuh+TjAIMspvwgq0d+UFcIKr3kKIQ
f6cnPoaE8mFIII2/IPMOgb1gTW5Ow6ntq0PXOcn7hCHKWwMUbJz4HjEABXVfapXFdp5DZ+eU59qV
HmV8ABYg7meRlZoTf/DteDinb6pBqT3rKmd2O5gz9UQ+XHwN6+dZKELrPRktX0e7EdQKEI9YHj7n
mUc5IHMIu8Wfxvual24/vNH4nv+kgg/kHiSJuo1hh0h3xUQFUHzo/DMmLwPx+ruFSyPF5kDTKo0O
FpDhzJ4VPJ+0NFdokup+AXP++M8zzuGjwaUc+yXKw6zICYpKTzngUs+BlteH0jxXE31BuxAV+Iyh
wvdmJp+G3lqQozr4QdDJHtJugPWRs+qoKYHwBMcl7r4ROVmhYorOzVykP7JT2llVJDIddjbj0T8i
3jIh6aDZ+9GJPG/pzYAHfp57nUkZSjHDcnAFHhVfaDdkI4K8pv0M7TgeiTq2rOqnpbr6rMBrzC5u
cXeEL78h7qRjoKA9vM7HhW3syZxL2GkCOJW1WL8A7Wd28mUJ8dGb7Gf3axjrktj7QUPUgfzDaaG+
nzlK+/a/zuKBp/SFGva9iv4PoiaEgk37r27mBKuwRZRZl0qTavOaakVt8bdzKWcLKAkLzItX7qkn
kPDJDXavAWQcNITMQhVbu5VoFhrZ9CrAGRr17JZc0sBB2aPdt2bfQDZspMRCwB5ItFXAe9YVd4pg
w9CyLeNcxa9LxHQVAcAloVrg3VhQ+SwNgIXFkKdCtPtqXswLIlPAwlW2cKkDGPW9mzc05btz7+Ro
1uTmLVLZ+uIeooSXoDFCcvvJ4RmndB1gRcFMYZaS3XvtFpfWgdZ0Rp4T4O7+4ibQfRLKym0Q8wVY
WQhH8Axbx2jsaEFtDmGyCW8vTAJ7gFg8URM8JJWA9HKc6muY1NhrrYQNUi6gUNixLArqreQsmh1s
x6B9yzK5o4LpnnHYUFlC8Yj8dIVhUTRrjR7jZy9xYsYG1FdCEta0i9B7O8QbDXTQwWNNd6zsPWR9
PhpVpAInhNqoWlhvPjg2v4EIxXOoaVWLipe/NjcYYyaa0kZ8U6znTEhxk1KUCel7fCU6Oy3QZuQS
l05ixRg1WbwsyuGj8Y2vo9srslVaisRKgX2GQD3MUvvGfZ25jk0cRGdRejNm7RpHv1G4h/t95JDW
4d2HOi14BUWhZKIilbhKE4D0jJqDGaXI11XifeN+dQWPai4Nxf4UNCoSHkDAjcthHza4R811ppXW
uKyfIIHPB5POX4JO7TkO+sZztZRHU+YxTUKOCqKPsmQ4tsfjmOor6FM1PI9tMXbxe4J6YT1L+K0+
ZTdIU9wNhWL+eOn6P7GD6mPxxVyg+TnyLuB1MUK6Xw+8b8QPVkVuA+lEiws9JZzPgYgGnnjhx9UN
yfv++OrSB4xVitlegDYmu6MrvCAPyUfgr6v4RX6oIlXTe1tSt+x2bmdLd8yvopEqWVg0TiJUXrX7
nqxGr2jHpnNSPSa3iGKFIUG3qHIxgbnNGXlSwr5QqgLyOve+0Fm3X+uSvBcRSEUswhvo2IdFyBD/
Vx+IjyJ1/LSjr3ReE+bnbjMZdpP4Z08adkKPVSKOEjBcBdacC5D2s/qFfWuJCOF2EueA/mMRXgPE
zQKAyoMCk7yX8BSGc9ILU7ESiSns4/pXoZl5ljvlRy1LQlbPwyFNojBkcXT1syvnRBQO/ScpGL1E
CCUSb8x+MXEWlyusMdM1mAQuxV1aE7ctBKCqzDYXFLNUr4YXXMC+YTRG7PoJ3oMvOIexIrefCJ++
e7qdzkhDuvaUGD8n9bv8OmHQx45PiQMR5rJ0O/1xNJAn5Y8C2n3wP5GM/XoEGAPdZjGnEfptYNki
cm4WvnQskRBVxMdjB60rHUYLrCoobFADo4MmtQQaJrVKnXnuzDqItm8oy71cmOnREMx7x9YII477
cRl8LYfe/dwif8aCRmhBHMgyEPk5KSlFupr8KQtzAD93z/YGCxgJspNSQhLkOmdwKDTbbDueh+zG
yY0mcG7BRQJulixuU6U+F8Vzoi2E4Gox6SFAChTWNJ6vQ0G5Uq0G5ERPAhg/WhVFV3UZYP6xxwNE
uBgwmRKc/JHEdrqbSviL6w/Z9+p9gMg92qeE2LvvbowxCv7k3P4eGbgwnslCX8Ggqh9NZBLP252Q
qlDegtM8b/TbVOl4D05xLrKwQHOaNA7VZLo/IuR6B1Te3Rsm2em2VBMNjDjhM3zcBu0eiM6VJxJc
/3eBqOi+FdrIGMPGbNB3w1mXhY63luIWE7vg2xU+IG9IF+j6N0rQsQtCzOVQpilLHUwbDkRYK+Zp
9l+RFQCc6+i/i7UUXEUjv7iIHoXRtgK+SFldOc65/XgybiyREzf4S4fD0xhw4AHpMuIoFLB2tp3R
rQtqXcMamoCMM9hbDlBI57VNL4JLW42eUzaKzcUpNxO82CQj2Z5firgy9j/lwp3zILN/b6sU4VAb
cbzn5u4XrP9kz7m5nVD2QZOkumQ0SA5WK5HUVqWtKp5Z3oQpLB1PpsMu6sC7p1EFn290fFaUIO9H
sZ0btsr7zG9lkQ54yafWxPxml1WtecoO5sjPDbmY5YqBWXR+zXg3xmEtN0rxWWV3zaLjAHtJqtjx
YSzBZbBPwv7t9xM9HLvIYp277g7Npfh4TydQwTeou4fuzp2LvE6PePChDMCOCdAqbxzdqP9Yb2X4
PZ96/j2Kl5/76B+pYLDqydIDyi7HeQZ0g2LIOXCXvhDvIQ51/aW9IN/oZRxXSVEji3AV/Avag30s
krkiyWvZ6W1U6X/IUd8Wzdm6bpjY1wxDrcNOHFSxP+xENLNu8zLUizE3JsIHYg1k7k0jG0cY4sLK
EBcFFo9ICQtkZuGw4KJiUgjkeAIx12NiwiAt6qXyuXCD8EpFYX6apR9zFahb3HPuFCj6Lp/r6n1s
Zvvaz7cbPd/gaAEvVbBFHtLi2sNvVi6qGne26zTiGHXIIBQKQSArXvrQJZ47gO/u3kyXzQjXX4k+
txm80vQvjJlzjVFQ7z7MZezEtfe3wu8KxDcZKl9cWHwWcvXcqlw8Dz1qcM19tGt0S6x5pOKxJ+LB
VjXZKYLVx64iUGMDvh5G8vixeYoyxtRY/b9clJfhhYAf7CzC5M7lYCTvNz8rUlUWSf+c1uWOBsWA
X4SJAwOsq7Kq6ScBPb3oPp4Hd2VcGwHSpv0AdvWDEtYQ1tAflVKhZhzVsdhVNdxHhMMiatYAosow
U91ZLYkVnZnlKHfsUaDymcKdqJEmmusepwCboH4MCy6/+vtBZmowQp1zH3jcU4nmpjTGKh0tty+J
j6NTrVrcYtDAxIxwU8tQGZ3YV8T6yp2h85DCt/rqgI534gjwXv1QnRXLaA0Sl+jeHdciUH+KnCfn
4YuV3YPHc71wYC40L3Jkf8ZJvICjgzl0Go5bD9Q2wa/AYLfC0SH0rv/QDxrskpNZ1akS1q1vjnir
l07sWaxwAPbsoYhNB8PXMZldn4UqWvedfHyCm8yqgKm7ErpFpY8UXNwDme769kS12DuIfXKfRe7I
uodofMEIALceuWDID/VrvWD27ozjJ6QlDTFD7RY8OUT67jEIMSkah0bouwnnQRkphovpPhslHRI4
hsJhZkqiM1wVR0P29FOXIvRXzJKjR6lOX8F4kgldChAUhW2ROebutK7mRL5tnKzAtvNXSVrCpRDe
NzPu2UNT4ZWFeynRQCI9XmlVbROXbneyqQ7maFVuDcA6F8FKxkJuMpmhwgjgrRk/MilT42m51rLP
g49fiSYP/84WdUxlhqEb/bsJv6osUgVRTam42VYTZN3w9IaoDieq+yyWiHxTAJJlbz1juZPKxyow
g0P3o8ZfBIC/YD4FwCEuby9z1CYcZbsvO/f6Au9e1SFsUJPshk9iTbpZe+79OI/eqeWw81lEREOV
rvpFE/k11dO0ZmxzSKLNP0lP8E3sd5US5R1Y18yGYmRwnFTfsC8ZXdAlAlw1v6ijLgTokJ8WT1Eb
WwnT6Skun6tT6MYvYuSlaBxKCIm4ARodyI+WEE8tmc9lQKbzQpZnh2w35WWZ++zjsCKdq3xQ6UPU
JQHSMvCQuaB30fcVU8oRBaVlppl9Ukg+lFqD8LwjgeO2DMlx9YgA1gReYxnOrlxI2PLa9Uj5nUPK
3vojuaXUcp6qufGbW6ybsibBzGJhzyH2CcdJfJ8h9cwAMiQe2CFzVBP6h+rdzae0FLXdrXRL5Ej0
miEWlP5rNSWo6GsSrpuqtJFoN1y8G9uiXfSrHwmYqHzhpzqFxitvPEfSrUr7191VRgF4wwBgShq+
/cQJ4Dy5avLAVYOV22ilLbJxx4nWWP9Y2lfRw6qIeNiK5XEbqzXKtaJheYynPtj8zWHJz8e1MAiK
8LdBsqG8/essmRiCaJITUKl1tzD2icoko9KOIGOlXTFTYo2yZQZxv2mdhimbPdrv/9XCC9sY6K9h
JBrLU+boCl6D56X5v6mCDPHEVX7g4/eh5aWgz/IgGokj+WY+faqvgls6ws0H2b8wZHZvLA36iGAm
FP6HD98Snbm2mrgX6TQ69P9nUq0DNM3zWzMd6LZEXkjpec1dxPD/1HNV2eYO9z3tCoROheWvXYWP
W4lafqn9SUEIVqeLJH721njmYyy5YnaKG8aUa9AkH8LmrMprXRKh44Y8PUDs/A4p5iN804ewSGqI
XfgaMqc1I9MbURlHmaMMoHl4lOkUatxQpU4/zirxosYHicW/KDtS9p0fu4q3sl/scEfgpFH25yH8
IZtPhdjZccgZvrfZKT0bMNA0AjRYFM8zh1dQRhV9NylxwbTm+JfrdQ4UV91hXbXxfZfbUsbhRhv+
cUg4hGee9QUMwT3ecaxU36yFH7LdzYSCtjgztAcPYV7ZFcq4dgoYpizMYZ4vAGOFSi1Naj/bs1Xo
d6i3Cc6n6BOlBdyMKGs0L27BPC7WvloPpUnkYa+NqdkWTazoeDsr+7NEUTnp1C+m86eXmEZtVRfh
DfH1CGEIbFGt5bq9JQB9ckSDVjvAoaeIrrLcNzWwdgNe5ZkQq3rL7q73zh6AKDzj3Kwsl0rhyh81
dQlWkctLNtTHv9VybjI4PMsTXF8IOG71odjabnORW8GmGp3IEJok6cYoRWGqAZdp/Rwj2hUqkCsw
MTxw90XTwdhR4GbqeVMaKwP9+tWZDwgEdT6FZF2cZ5d/V49kH41t2gJpHBosCKeLKXmOO86ituid
xu3atyv+7wYm9kVf91qmlQNdQ/kYJiz8ZFVs6Fku9hQQOGLEVh7i3n5eI1842bkuk0O95ePgldVV
lkuUN6xmqug3pVf25anOylR0Jb/tmfJy9+ndZQBEDpYREJ/0ZReQrNA6DRo5vTp/bWTvn/DYrjUg
NqPk4UDuyi0V7Fg9jMteFeT3WjK43gysPTkXZ+T0kZ/Aj7Ati01HCaBnUIQggclhR/I7gUUEHSJX
6CA7AEG4FwUNfLNopJUcPfcSdGCY7xHa8UoW+hdVuCOI9nRwlAyM3KK2tizKBG56aC7pekXQuX4P
jRL2KcIlRLUQUk6tUPJ5MQumLzWgm+fOmOSFSLKEgJkt/XR3d5oeza/NfPG4DxR+tjxEcPbVpKpw
wF3DZlm3mVekD5HQagAF2nGKjE1kAZyEkp91xXBOvHhltMldNcaIjHW2yEvAFmlju2uP4JvM0wyB
9nM4ekq52EmTZe1wE7wMfY9k5WBZUtpYbJZ+dqqJwPFHa1bioUqmk8QozbEEXhmKRRjhtryIvKCH
yuY4QXZg/uSV7ANAuLzXXlVCYddYrs0MtaZxl0FsuZfoFK4k8jhzys1+fP+oy1eFaYV95L5mAero
J78blf3bcly/ofK3BZm8AVFGwwwp1J/m+8o4N7x5Q4LTXofH4s13cutPt/5Jn2+Y8qVWjEap9691
nfq2q0YS404fVBH9BTbYgyeXbvCWe8292HWR2JmzrmwOFim+q9pTTUMnR/HSoWDH+V42nk6QjoeW
+yTIp4iFAZ4uzfSUFIYkyBucdQBed973U9Kc4G2KWH2eW3V8sap/cDyAyuFZz5DcJJDSRDjhzuAj
EsAJ5abu6EvcMzn/JHSDohDhd4zdmMMBbfa1ratj/vCXPEfw5+ZUx8YxQD3LqlacI3EYV2AGxTfF
qY3i9aX/NnOrIqql7iH6o41dvDapA3OVGTk4FtBc0IPUx0rXN3L8jz0YtX9ixJbjkYmEgXwAdX+e
4fNgvCKTu5zdPtSEgTpdXZaZtB6CDOeOF6g/mi19VaeA0AMN+blHP/+I/blSEvBXdPMzttLqmOam
e5jCU+AUoLyGpDQPgXv9o79idiruxr97YRGuTThW89OMp4VNmolywX0IfmOcUpAjNzP3+it7u28b
iTWEE+qPQIDHCOVybHamR4e1ZoBdNdNdqZcPzUGcKjurFfEI+lVnweIXHQGlnx26EU0fIlLpocGz
Nxl0+DLGHyAyaeJOe9bUHn5O7cMK8SG5+oa4WxX+PQMNVyxnkGC5foUzolRuzdN78486zVZos7JO
PgNCVGZD9ClG55NbG+JRMMxwvcVQsNHvAMXKg22UvFwd0cNQ/MVmDJSE6gBQ4QBKdXy1biPf0eFw
hwluYknUss1vPqqBiUCwaayjEH/KhaXYMQX+R09u51ViiYZLJ27oNBucuyQo84vtpKkA8b7L3i1d
U9qQbN69UfgrX4Ya23whyVqo8GdtYffw9nQ7ZGLAITVBUiFWuUwRXnO0z87MDO+A5ENU/YEIqu3w
gOSNthF148fRbh7AlaF+UKsBw3C7YdsgYuVpZMijx1y0zZtE9uSK5KzMy8WLjZQVgint8tS7uFTt
Kd0Eim7sEpb+INtK4yWFv0Q881Id5qJi++Dnd8KZK1bi8eyrYeAepbUl4RPivekKLca8Z+yDlRX6
aH+/O0j2aLkFv57585AdOm76ks7ktRonrhvwZFQ5Gihl0aDMdzgDcTydFk9/1poQ3MWGeCyrLSIJ
LZ2D8F85Lq97vQXuApLmU4fkTC0108CJfu0KiY4n3IeCMxT8e3iC1kSugDflwI3cxO/g9Ea3j9ht
AH+2FmjiCrR+SUFM1WJ9x6VhwkncaABNxp/Rq/5T6YRQ/06+SInhooG+C8Rdiq/qmy1R4D71Q1tZ
jH2i5Juuxr/cQNUF8M1wxra/btYlSZAK8NSRO8+TPo8Ur43Ue6aTKeo/dB+WhHuL2JU7aGgBPEKn
mGTWQ+3WvwGV7r6RzttWKwJ2DVI98uDv3SPZDDJQLvM1D6TArguDRnQBysw1ExIyloeUeCdH/hnr
K+1Z9sWdkzzfasjgANQ8Nmxc6nSXCxBYi4PKKF3K8ueChIVrPyaos9KYjoVoZwz3vcLM6e0DwII4
e5PDVxhwxLqqgBNe7qQwnfvj8ILDRBanZzyZYRYFglxGSiC0dzn7dGMRcXpM1LvjExtK18fb85k5
IDAs3yD69XCNacBnLfpYPluS0WNtBlgcfdZ6c0NRsN60ll8+9hr86IOppMTMFUzl0j1n/0/XQEHl
m3IypCBxsBLovW3BxEFPf2IicDCto7290PqssUHkutcr4M+hYVapaiUtMDLkbGnMrRRg9CM7Gy/E
hIJjdOr98SwR6kAQES2WR4Jn+mIDRNQ6H82mXY1ZFmvBnimoKR/e8inE8iq6ieqRkM4i4MBsKHwS
gVAWdQM1p0vPCwbDVoDqU31DTZS0n6jsr9Bhqb2DWk/fMhYMv7vMYKve8Go1dfHLnb+u2I5WxV/0
u9qb3W6grK8kCqpxgcAvP1q0I9lUG7Lar0ifdrEX73JgoMmhcZNh30SmXCuFIDEVB20MVdqIUwVb
GmMfQ9tiWv/xHk58T2YEXZQhzqMH28R34Idj6go2zWX8/n6bpWQdmbrjgN33gdxC2jFmTKd8rGEC
5oYc+xbYpb1Jpfy+yhlkVm88DqAg8KAAvD4yR5IkU6mRh2OmYofSLyzI7Nhthxqz9MR+6g22FaTe
w+qPjnk5wdzlg98M97+lsEz7f7AoP9y9gOOIAGIlnZ83x2aiameRVoFqPdDsz3mskzyBSvUSYZUn
5+e+iNcF8B3TXaahVawLXM68/9cEHX8YoQxqzeB3PJVS0LKuFcSvDEHYwPeVw3EZsdzrExaDqGTp
dJt9PDxCAufyoMLD5s2xc9lw48G9VgJOo4RQltsqfNBXvCDxwDsFFIB/gWi4Z+Qjb+AiiDt8M2C+
dZlKNIgYihBAOXcuuKKtOqQS5jMC/vhlS2rWOUbhaHw/xzG+sN6rx6s7niKmo6+d4JH7xcDvU68F
PlhdWfFcz8MopywV73nmPPgZaAn+w+bAM9RE6CsoWlhPZkkeniSocRrhEmozJ5kKZJiZqitJFRWs
38URvSj0+t+3IP3Pyq3jCr0lSaKAHj8MxR/mJTy2+WbGHnfLZ2fC8dCl5xvg9Hr5a+Gtvn245NR1
ESWbnKLvflxrm3fseCl0mZ/jLnRtajGSHeWHWSa7MtR/iAVwkPpXmOMPi7/JFnkUhCFXlgACfKlF
Y4NDzexiztVlddDHgutEwOdXa1XtH8+OFzt7n6L4YuZl7yZZPPnCMYX6qZycqaAVRF/TgSDZVDRl
obBF7EzjeGU7NjChckObnPQ81ifQz8ZlQ6DZhodFZeJR63QVTK0zrGClFeKykBOyhRCfGuFeiCIR
28YUI3yTFYEHwfk1k+sXLccnqCfIEo6Q7s5i0XQJxj+K5yB2Ghl8PpvEmzonCDpC7FHw86vGe3kT
50hOET5ZCVxyu/Wa6p+9SXtwBDT4tAPsTM7NFGu8bVR2HJogxhGcaMkNe56Z1jKXCjRuyw2ybJP8
p3rflAHBeriJWRuELI3PKwXaynQFzzNQ57Dgx5Cc0L9N2Z48WR9Jl6tW+FRNauAVuFdatxUi3z0V
DL3bDDy3zfQp9WQ3JK1uNaZQMuIAcWPigDTAfKCXEhPLbwf07lopQzpkJgZz5LsgMcVL4dCqiKao
dTkLqfvSyxAJHDAEYbIOMQeQQjhbX5u2T7hTPT04fQsRG//8HEEZ2gd39wd8MbEsz2N2f+g6ly2O
jNEPR5LilJTk6vfpn3i1v+OFtobXWL81vtOfwbqiAozHBMvDdomzMO85NeGkrbh+V3hszfvE+nl3
OK/CUZ7Elpm7a5o+TkxxvIc90nWiEJVYi41jHMoyRJ5RaLL0OUaOK83vu7AoQLbd/FsRTBF5gT9g
rhN+3JVfh43n5Sa1U220rCI7GzVejtFxeMfYW07Lphy0MKFDERbsu02lBSlQ2u1kopFjW/EsWeyO
P7oQmvKbe8u0BB5rlGDNH+dvzS+ltxJeRBAoem3PIpCu8fjkQn3XZKdsykOxIahz1ZI6dH5ouxeQ
g5CFLBZwiAosAwtqEXjfajWFuTrLeGIyAdtc9BKJuFtFDxR0qddEhchzp2AoPM64ZYIfa0kOLSb+
xCjZDPRrb1mYPWdLb9t1mnN5Uy3LfELocqssPqlKM3UZ+v+PuLaukFSiP25woZPQ367iskWs7bWg
71f0Tc31ewqibk8KNyJPXK3b9oZ5bykhkAK/UnpsLIsbj/otJdN1XE9buC8FhVZKmozHRR0DmILV
R7Pl2QmP6x5pTgbLTyxrw9zzh7oSGA1heQoWWS43ek/yo8OQBJBp5Gxn06JF0W5sXv2bw8r4CUvV
5eir1NyQnEfHYKLpoL1PE6F07xXcI8m5ATCaFHmzCBPq/+pTmI28l48xt/UKQLY6fqP3GCoxNQoF
a5hcgZjei4S57W81m+gzJaMu7op66IKnXOMU1a4DP840dkJfsMb9I7y8IQ6kaos48RnrnIqgyfCX
J5cDinhz50jdzXFIWkr6wIKDDFqjQXC9q1a2wHYMte1W7qZvT+28O4H62gA1NoNZKyRel5ix1iso
VX/imWO2DliIoW4w6tkArD+gAWPDWHuhwHXesEu/2V2+5xeEgY8r7djSw0LIlYp1CiLIWQ3NWFwQ
QFbd1iOax1ni7oBCQOgEN0sEmSOOjCdPLzM/wQnXsQflonTV+AC3VyxkXVO0RhacD/YNtgUbfGq/
y9qt8TenEBL4f/AH1YO7/PLs4YDxBCe89DalcTmlgbfJic2Y+aNBsvtlu0COZdGhUGBFe7nbd8UV
FdG0PdWIivtWY+P3k+wGgXOukuK24bPTp8y5FL+0ylmtFc4JUxlskQlXdCIvoZOCkeZ+Udgtdjg/
t8pJOISApL7NPjP/6RFyoXBfHpmsqQg08owpxqimqCrLx0FHnSh1MRWH2rITTgQNhmIh02OxbNfe
Nbn1TrkiIHTSruvkX69w5d/gWcnltbbrhOBGYZ//juHmqvzLLzrJGcTs4Pi/BMaX2+tea5lLfBeX
LjlLku2/pz2QmDV+IU8WgDJ2JIOMB/tFg5kDnykjfentVts3PzDdtfXOIUCEr55Hzk9qNhT9BOxE
5pQB4BbT9xE1NTIkBApzwOJtZ/EfBqKWwqkp165MUWsr8AFsuTxqM1FOmUydW+OJ111aHDV1y3fV
jAg8E347se8qJuSFmbgmknm578sZ4Y6lPaOelK9T1jivuehxDSfg5ydg6oiu6RZQPSBE8OqGRqud
9c7vDT98eSoutSA9XuXF/ql3n0nfglRfFhiwRPmsW9RolAp0379ZD7FnsIxNzmRLqUTnxIsIaajC
0MXzDHWz2hVMXOxXmmIn1ab/+wBFi1KnDisVtRKO8zbacEvsGQXSNPywBUhn+v8xIqIqClcb3Ugn
3XLicezYR9Oqr/mL33+5m4ayD3+Yx7l5v1y65z2f79EaVS/Na4tiI4ljwPqPjo4+2UbdGYQVmmXN
bK8dyolnu/YS7Isjua+pQxmmBsaYkUhWm8I2qMfSNrwAcxfF7jPkMVhbT6CCYWurYfJF6U2VdUoJ
CDm2qb6rWwSucKqAzoQAdgVFjnD+fDJ98bkH8zCDAw0oHKl5G2DqSPQduCNCmUQGYZqzYBKgYyfH
C8SzCQYQszuOzdYbYh4zAllkIP0Ca8NjUbsDqBHxzx6PC1UhkBV2Zev3KJ9fEzFi9rvRn9GCPEmX
8JHFObxsK7h0+7o/pM23B9R/x3Gc3Mg7g7d72EWL6r94vrMC/GbVvVdH3L3rehv2/qJfYSdjY37Y
xqTwYvcOA/IhwypBoP4HkPrQ39bBEChSzHAZOMDHN+xIaL/Vf6Opgrz7KCEvRzntP8tqbl5aX0Z/
g9+GkI8DtwxCD/0653uLvijWzWq9gG67tgDtxV9dYvc0rUWEtlzWyRRCRgYoi0BRz57+X9DaIz6T
4e55IW40umXwOqI2Ulch7S7DB7/FHXC0L4kx++0EyMUCpPIzgIsiDYPECn5QlLXqkMu0ud3Nu8Jj
MOfBDHY305+rrb1wjuMQN7MbPbnvmp6R3UZlTPjEHhAv7bWvAug1f3j/a/qzZEazhQQ3rvdWyrPD
Uwzgv/MQ1hjFCaeLmM8ffce9G5HIajQiGsOwg+JaGiHbo35EvhblOeB6rMuGXbf2blr0xio0rbAS
MPjnorIX9bxC6mxsU/4da2A9OqDGX44f4Pjt/EPKoUOFWQm88z6zlrMYQ9meuHLya2VJFBB7ue1d
4a9qCB+vba87Fr0zbM/cVNt6w5zgqHkQzu3iKtfdIht9x7c/NPVdO6CsO5OkOmxawosAdrIO507f
+ZM+RPd0+jUsKqFtu4u4g9yw6yNfu9aPEfIP53C8g1tO4enX5MINYrQAOONkH3I5jvPOAMcXELUH
1sO8ddDQaxf93YWpIBVPvA1Q1EJoJIqy9t68GdInhDICNIWWx2djmBebud7Tx60I/X5b06AhXHoW
E7cdehtQrcBhlosqQ9obxtZfTbpwKHjdsGELg7vUP8GFpDK1TuGNAo0lV6D5RJb7KL30dk2/K6Fd
SYGnYfN2EK1rTbTR2VmCXXH2bCGDxWXs72FTS8ZL1NC/7DgXp3QszOf/VsjQ9DXKOPfV8hosbXmd
WFrhmAIfmD3x+4jh6OjjFXTEf5xtCfC0gQ3+cMvEKsx39JRyO3QomZraXN/KSTJ7nK20GFu+PaSs
0MRVZWQPhSmjMkZrSIICzVoiTIC5wG3kingfMH21PzwM6lurIKwXUCOhEiu+FGRCfI5KTew64qkL
qlxk5s0/XsYbSbNGL3lE2WTTZDfwGBSu+2phBKtj+JX5tYzB8Y5Mr/yRbSNBwcqIItFT2XBMY0+R
NinKy70GedmuxEh6YDHETw8QarqRtuGQWWvzA90aviSD4556NMk11h43NGoMT6NpICz64DC98pSb
ZeXQV8knjE5maSckNfuCMqkZrNybuFfpWmmZd+737Jmiy+EQiIwIrlssM05snZLq79zJYZ4M6g9I
/Kl6RAlUipXjrDXafNHtI359QTvO5w+44zz6MJL+6RB9lXlLkqRbHdO878RUSND5XpjzV+DiUmUP
Q6W69iUbyacmEcwRK+TxA0/wwIUhEK5zE0BKQ8EkGAp6GTTH9FEX1aBRT1EOrHIIuyj1CTm5fmwj
12/jJlEu2Ww050PA9RMAaFkeBKkc2oL0relit47aSikXKWpk4ko4Zy+cCgU7HIiF30oAU23g4jFh
3i0FheI5c6/V0PzK0exOXhoTs51Wc71TBkjxW8+Anlk9lWvYHTRuOdhqCdDNzEm6YUx+KELA/7ah
Js73I0JHSDKVoHtmxcuFWQug2Hys5qQQY/XdBHtCcQlVttwuR3IdY3Gqf9G+RjHefpI7g9S2tho4
skUD4hUt/PZGtfY395e/D5ielngH5+24YuHR897ExX270ouLco68+Ulk0nZl/ZiLl3bOibp4BTuo
yaTnBZNYUb8xmaV0UIXKV1CdF7MWMimaM3MUtXKVXHFwsqcEPUtscafv+HanTcJrKNxFCHSzuRA0
Ur/AixYXADUDGZ3lM9pXSVF+HRpRE8d0ccVO2f/SVuSGHYxRHwhVGNwDzHaHxrMg/xjLbhBtBqUN
Eq1gpSEvCc+J7jGiq9r9ho3UnKEtIWdzw+fZvugrnmhJWBnZ73VlDHdWoAQuooVRAFSgvU/Mb0hs
zKyJrliMeeRm/ibeAk6PXrgq50gjqg1KsnQmalA7zzmbu29nmBI46I0X44U80zaFpG4uzpXaSzUc
XlNcWmKx7cY5Zdg3waWV7NRTdkLpfsUoJLCh/xyONMja8q5+Zxpq/LYtyorRIlgICvH51bLTaNVy
JQu7LKthuN3iQ9JR4Zyoz0Sx1zu/ZSkZAD04Z2rQ+Q/u4olhMsqVQJX5a3rY62UnLP7eT+kJGzEo
Hk5TFKSUtyQcxhVvoZXGR5MB3RjVBjxtIQUyNkUGq15fwg0IWJ9n+c4pgT9rEPEouB3ogBOIZHJ4
6aR0qpUxiSyALNr9oZfb/fWguny88hu/uDi1ceGdPWovDXgXD+5xWILFr+NwwRq1XIQ1Yp3nP5Ib
3mvR9ZgYP0L0Ton2DdlEkXj3tk+2aHhcGfxuM6t9lR6saYkDp9Q1vaaAi+DahY50bTmpsmZs6/p3
9C4yfBROY30x+DJlY/o5rmqT1AHI945roYUkt9WAoWwFefDF/1z6FqaG4Ln4DYVJ9PxAxIFsOf5B
zZUQRQ0HxkqIQSMHp/prXDy3QdW7H4aJbskT0PQsM8Ert3EhNiHa34TyRl0v4wWrP2BXN0wbRMvf
znmym/ODhQche8kQ2QBMXN6NoHfhZp1ME3F6oM30adhQwT3mW5oaZsVE3ZDPqVCiO4wjPBySOdxx
G+5IPSAf5jdxp6zlhyy/JsVjy+NxNvn6NJQIDAL3B+Emrbj7Wb4JylYo/l4XCgsAzTbWycm+kIcq
nRtWJQL2CqBRNJl63DfmQFqPC5YCc9Fxad9wnUWs8jUKE7bMuNH0/4lHz1TaV6uoxbuPpCMc6lI3
hZFKdciE3DgyOTVGsQAqqG1P4599ZNDN7y+jQ6hHxXFlKMYCtwRyWhheXNjQXWOcKdawcHdOiB6F
1rnOIF7ycJ2y6iPwIguwqPGiEuTn7QeHzi1wEZXQQsBkMjc9td/lMKyGtAZMcsUBcpOva4Qcm+Op
ebwzssrryp7EfvPouK2QRDqfk0FrXShfnaUdb7ZB9a3kpQETxa9VksJdAvlH9tt1GBrvqaMkgTcG
GepGNq63AehRtRdAtBZeOSDZXcG2AZZlT98YGSd2fdyxgA3ND0OpneHz/9o1nY6yKBuAHItgFqt4
7AADheIZrpbOvFpBRfJG+9/mi9E0Y/PMVtInX/l6v5Qr6MG7FoReOhHw+SZEmFdOsnVW66msRhzo
hLXata7zI28J/i6n3Osr1YhFqzPavdmWZLD+ZJa8Cjd5fTKpZIF0A00R11ze5nhNv35RO/yxWikw
zwigJ1eMvKljo4plP5jbTa5zIq5C3vnHnSLeCxUkwrfpvw6KqSa5/SBfoeOOZIYefJPMMwphWiQ1
8iLGNgZav+IKDKIK1W3hJY1G2ke4HoadjMibrUvMVEB9tgYGoy0EVmJWwGVoDIgsOsfdqAxIClDE
1r5gVWemkWsUEZ0n01aTKB3CAWLzPc26gWB6sqPo7sIhobgGHNtET3shTCPWO+qZKvy60roDv56d
kEeOCvqRj15ZOfjvmQDQ6N+60A5OZGpZkzD+2RYotjsGVtwda2y09IWao54o3LA6OS987OBCPeFK
Izq20ulCz8V1M+TrFWlHiWPn/zgULpBjERrakv74eML2l/tUukPYv/43DIQVY4KC5GkoL1cGcBAL
Rr+dfrSbv97PNs+qmMr78Uo4mYcHo5fshBZQBd7gu4WT0Jn+xj63TIVNphelVNw61fp64vrp2EZL
CzpXhdKVGq5TcMAo8Hb2RJ/iGCx6XD81SGnNMF6+SHNSLchLA1A0TWZ400PZUJFzABgNEkHFjLE5
aOoreKlwAHwbtu/67KTlKVPIqNo9kyGwrJmk8geQQQUY4tTrH2ZxNXjC2+y5+0FZmxPI1wzFc5o3
RTla8XTHDBNYYB31Orqot5oGU8QiJnt8rUopNVbwkqwXKEsqZFnDas2M7jlH4RI0d7yeHCxJqyVJ
AjSEaf+/QkEEcmjvF0zHnrOHCQXYIXNVxZ2h1b4PWt5rI2L6Q1b7mTTxJUQEmHPmYb8pkTprrfSA
BwK2ULBSASpNwA87cc37gIVbGWkLcpQ3hns4yvhbwwCXuQsT2a8D9dwLWz2TbAJOdhG0kYgnfWWF
aebA1dGGhprntDkX2SBXPs1BMUTMIN8RFlOoMeyDWpKtX0MFvpYSqdFSajc8GA1cOWkjWjUS5ld0
G0bg3wAF0WfGCS+mdT4pSpOFobzDEAXIr4Z6BTg20yRn77iDHAuoK8prZ06zByuP5QJYfTIGY1NG
yMXFnK+MdBKn8r2826+Zy+fPX5gNoTvhMmMh0MEpQSrhew+fVrpUmt0gXMNz4FJYUWyHe4mUcXSb
lPCpioT8D7i9s6IY4F6roO80MgW0ykKLq3uViYOtno3VWd6mE3boNDnrPLPHL+g+Yf+KA0nodvpd
bcdRzAloQg4J5i4NInQEfpbutIYjOGLZml9xLY1QvjJANrZ3j1oXUUndIB+yw7EZJNX/JirEYKy+
/Oe7LJErPWcqYEzf7lwp5b5z/7ShRhchSAr/UE+y7oMvsrwah5LDhdDjkT5/OmxtWMgEO3I89zWl
r9Au54NBDs6JIYSkY0eUkfZL/5Z88uW3nzfy8tIOW7C8A+Y9saLKhPHsNR4UTH/pw/S0QFfVF1uK
nLBlkuszGo+jdORp6wJu4RMGy8QJXC/FgCxZlealKKa6vSIMY7CxGJhV36vbXp9VSJcHNphbzAoA
A1bNwCCeez78bJBkv0qQmebIleJHi8V1UhxEaTI6JbtppZm/9o2rlnc1oOhDsPCQbgoFXOPlxA1i
Cu1E5+i6NBL5zcC9hT+NQYsKMed8SVWmfq0deqFElc7OTTTSf9xTKyX4URIRYQEJ29PzpbA02AC6
lWiuqqARkTOK3K/C/97iwQVaifEchyV5iPCHCY1SzIDr8hYdqKnuiC75dit5x3vKrmcPKE4GYyy0
/3iLF8g4tTKX7GALJvGJwWiBpxNkwZshqfAdMVwGZjkZrg+6giolrT45NkhVoY3IOC0NxfKmSk6K
YN1r5OvdwxkhEUEPhPrFP6fZijThrLZsIt2g0fN/BJZ3OIEKLYqgEyETyLseUyjPVSvyZ4aYpG3v
fg9fNtty1i7zRsXFNGlnPhEWhx8y0wi3Ek6uFeabkaCT89KYrJQNKvAhdXKMCg1wUhbv9W+zUayW
6kRH8QC9nBOn/VPI1BDs/jTX4WwPdzTzZTljE/Qp9ZmbDQUMUdHvMC0qGqiaWYx+eNvxhdydPWBC
7FDrNLQfWBxs+vVO2rQjMnh2+NaNbRePz86FuOIkLWc8kOHNH+nVk7iw8ayHtebc9vh49UOeSDkv
Xv7hOCEq8uj5k2CnY0XhPAv92jwj2ZZr/6GWBK9pcCGDyqgefardEQkOdTErLwHEO5SZBPHHQPM5
Dc56mQ1cliYxnptClBh2Ejx78aZB1cgqEiDhQEKNNsQuD1e3O92Y+qvtsODKM8h/Qus3aiYoMs6k
lZTeDscGqNmLl5TLzHoRHWdv96YGBl6mukqyHyrbOU6jPU7VOlkYOJdc22wKGPs6kX6GXdwmEADD
+1cTlVwAVS3fWNHsoCdHRs8lMymX+pKkWX+z+Lv/g+OsBjR35SHYLko6jgVIrMEvEXX3nJhBvjzm
VPd236qGdyS/DaKgp86WhT5rQly9KWlm2PFQpqLDdtJ6J5QrjWNBtdheuHrTlTZrnxPiZl9Se+bu
YtbVI7X+cNJ7YxOrH8UcaXoyqCvfLyuM1aKPUFudlgMtokWi/8h58IbSSX5qPdcjSx6oVxDneCKj
shBPXtI/xJJaMOm5q5iz+CQdW70+DL9FAL5Xynq1DHqVUSuDAfYDqJy6Wh2FXC+26sIevjTSh6pz
eVAEG3z7aSA7s7U3cEVCTxTJVPf4bmI9X3PP60/dNOTFjL7j7/wT9FBxc+/2tVQz2Bk0e61omHy6
7P89eC+WfbdJkUxhU7C/Hte+IKEgc7/BfkqkySdbjV/nLLL17JFHqJHJ9/cuKb2wp9wUmcNhF0p6
hB/+Ppy5FLplwM4r24OlXiEwv77X4zsp+VRb7SEpk+++10jBWOJG5OGyszLbN6WibZKCjLnct8v1
ZKtJHEmWnEBWTqpCQlJO205g78q/VYhheWQ5SugfpFtnNsqmmUOz9oVbZ1WzVevJeZtI/WwEgbpw
XIMKUJYLTJZ4wgjOZIbslLnWjnwoQhOoWffWuEM8kfamUE5SzSF+ThWO0uq2GYxm3aZalBygmHN3
DZ7bSXPB0gagARq1C04GAK4/KMuuCK7VCIKs4JQzQ1cWfEY3X5P1F/ysUNGX1EuOOM2Ba2zfe2+T
40pZmqsqj/1dyHxZloPhWiSIzFXwBkXmIYekmL7pSYRkDc5x9fE0n40rmEBEsWzMBaV+mjdhBUQ/
sFF+WdLyop+1bFPKy6lx9HFM9LM87rvX+Gk5wWIypkNqhUvCRaO8uu2aIVufmAQbygjYHfW2fNY/
IyAP2cdEZsZBYhEvhZCSFvX+jIHvxnxen25b7Vg6S02p4F38VWZ4HiVJQaZ1ysA8ATodkhh89QHR
1Op5ljSwfiZnmYJlG41LwUS9fwrKudVc93Igiw0hVOYtZqTstpKrt0RtiQCG2lrmKnLBXQ+X2mhC
hfpNWWXLCGv1l5lv3c43AX0DlE8wpyk7fQZSCRDrc940g6pEisFndJZq8PdTvk+VRCGufKJAqIOe
x9NmduTY9lH7PGjYY81FPTgUiFWzMzUX2biGMjD+eKHm/lj5A54Q4YQOFdHv4JDTlP+KJ9KyShsm
w2JSyo1Ui+EsU0LiitLLCDFRra2YaWiYiC/yU7XBVlwXLYqP/er6prr/5TtrqVh7iHyjB321dvQv
+DoW2cdVyDLpOeZ9bnSMSnFAppV+rQG/ID9NhD9RNPgU8ludVUe5B311TFtXE9nQsDL6dPQ1K35h
SoERjaeW/ghbCAtzgG4u2UfkwPKNBDXwbNaO7TpOpi5/8bF7pvXVfUh6cnx0+CFXlY0+XaDyAKdW
065g7D73YMXMgxt9KuoNqiLddtPZ5/sN908h9eIC4D5uPT1iHw84E1cKPU3PLVkN3Ivw4P7n+C7T
fTIPivQYG4YmbSdbns96btIRGBUvjG0YLAIHv2CjB3oG40EEXBVE7PS+50YJZD+shCg/zttq4Apl
oWFn7n6DMLaAGtp4u6fdHd/aRoIqlGvHJRVROB94JtL9MBnIEBWxCyV8KGnKwBQKnhxOKnH61P7l
oOa1Xs6EjRV6oEdXpJFc42AlpfSg8gzORbAo4IvLmZlTaVdUg+yg91wzxis0IhXK81N2wq32N2ad
nIvTtjTxhUkE/QKLo/Cpd5qywH4l2+e1Z8/0nhKlthTWuc4cuyDDuZERkwacjTtAJAvdTe7Q6oaV
byXVLrDDIMVJWyEoUQIvcrFEMSNvByg4qPaEUjWU6P78qm9LrnFZTq/lXkEKOVyAMzOhyDq1tIZG
CVJzmZQcbyTKxT04H1VzGT8+p/iN2M4QMbDRM02cR6uOGbJFZf5GptNuIoTsCLh8L777JcAjTckH
kgoGWCS+oswCyi5cF+DTGiDme9uA6uSPxnSn75tRwuq5MDA6ZlOlxThi4l7f/X+7TJ6X738CVB7F
jWtGumAEOFGnkNFbW21vu41uRBIKIq4ODpicXVmf26C9X+Bvg7Bd7W7XYTzl3t0jUYANJSjInY3b
YfMvadSXgEWOX3E8+IlcVz8gr9Im78VrDvGlLAG7C9FDO1kn1L/7CNlExlBPrix8MoSmWKu0yRuu
U1hrdXjA+2l6g1+5OJEATvwZyLUs3nVXDlNY+6uUpqDUIFb/HwagI1PsGFN7yleFjV/p6GSkyetK
8MiDNcpi22/s/gGYLuCZibvEgBA43iDjJrd9SqAABmc96us2J+AuLtpHjArusiqXuFu82TOxLaPn
yFpvYzFeEBnHxW6rci9zvvynQxLShIQK9CcLnePZCSevOdZj2DFwr8PG26E9L3/uQZKb9x/XLz03
phTf7ainYAnwO22T9M6EPUS1GvVn6Oq0wIiTSrNVl4Nkh3sdbHHIJC6l7L45jmeiHYtjPKNWXlRU
9e9kM+NXXJIcqwYv2I1zET/QxRSya/Nt9SQmhOZAkntiIDBdVUa5X1l6vGE352CHCmJHxh16E/Wx
Mfdxor9XS1HQeyekMiqQXVhp4l8DvYvGWGTbTVoyKf9RabKpOYFAST+AfUv5Hc7+O2N5j27Arp9s
MvhtYqtZLG50msTYHn2SJfc7LFC1x/8vUI9JFiRdhdcxE82C7hSOEd8qVr4gpGvTHxxGXHC4AV5M
OzAz5FGGz14bLTdTfSGKism00vkL42nDzVQafcVKpH/miFPHdDg6ijJLAcBs9LXPRAhNdeEHO1l6
XHVUf2KdvjQvdXuKA+qAF5amYkWf0DTnTjSyymhu8NnkH6qwHFShYBZK44M1Mq1jjR8HHWkP4Lbi
MtN2NzQLBPF7vT37m/TwyxRFWTToMeTZYvA6t/inY/HL27C36Y+oyTP0urIGSXZls4Inzubcymjo
hf3HkPFSaNf6MQJU80/8Un4MKSzBBtgGRc1Ut9jl+v+rYLNP2qvGWXUyPrqYPw0jfVXOiy0YZK5E
0swBsuquLJu/BxYa/PYix3jh1ZujoMBDMYBVkdgR1Hznek3Z2Aw/C+KPq7PrDr9Lx/ZKT5t9oibz
klrxjo2St4xT1b+7v/VqWu725xe6lu+237WNijEZsCWsmV2OFXFYWgNELWkhugy5s3oL8oUvTDbm
gVDz5DdU6dIubI1/RlgIjTc7by7w40e9qjb/S1zHX6w9plBXKp2BBxg7/0hgdZ46BbtduCqLgfTn
z3CCuKGSvQyoVRDY97oPuRS6TBzv+VrpF8SrRjCFXH8S1SBqKnVO3FIyr/pqlzEAV5kQPAOAvVqO
1u+FUInbyIlRY4Nu91Noh/nz4HqY7ZQIbGMNylTCHFsZrhP1DLyn9ntOeWCnbr7QQFAwcK7XeCoj
3kyYKQ6jSSnOZaruqj2LpZgJ7Xm5jndmKkbW6Z6If2psCAQQxjk837GpE24ni35hxteTJyZniC6f
j+ShdEoEloyP8rbEoEQgy/6UnplnkoRD0SbPMfG016LlZCd4Unzqn790+wKf0k0iqGC5ZFeS5Q9l
TrJDSYD2r0sd6Y6ZIBcWS6N0Y+WRNgnI4Kj8poLRm6Lved36Z0rYd2+MWzAaF6cvv7a79ZLs9Skf
dJDC7/qmuEMFs2lzaF6ljIWezhOgRoLXU8nnx4FWLJEtDEkKy3gxpKIOHXX4eHEF16eAYMN2spjv
Mg+tFU+JDtbItvDPs3mglrKQlKBwjCg6AopmldB+xcZHX/OmxRdzpHR+6A/1R4e4QlgCqYzCTt4D
DPxLDHNOpTDHvFmbK7uFWcQ/NEXKfO96h0U10duBBzsoOheRH0JCjR3A2VCHSpvLoQVCf2LtTgk+
WhxakIaFP2nphrmtVta7h2R+9NFqv2HLhTJGizDPfIICdIC1UV8vyOZNsx3lQrJ9BjbiWhwkp8Kh
u9aONHX77CgdaNh6In3XKKPGJH0KyMixwlqeT7wFcM5mFYM+b9Xrb8OTRCmj5JmTutxy/dhXP034
ppjdl2MsphbiIiPC3fSdKJiJqkb9AHlOYlIEOA7fS+DBmVByrYci3iCYGzlq6W+qHLu9XG4p81tJ
EjsZ9IztAHoCOV3+klglxPzsK8bFbzipZdwPvCGT8wHxaMhcyR6rtkhXRGHcp6uAcqQs9CfjsbdQ
AioY8FebFupXCuUjjcC7N/A1mP/ppxWi8EuZlyPFha1PDndCisLUE/U3qQUOhwYMvWLA2xxVWGk0
rMaLdtIbvJFV6GkpjY7kFeIwzwDJz4k0bsIrgel9j0y0Ho3HC5iJsdrKS6tkl7GIgZpeTxl7MIVc
ML3FUG1FILnBibKaH/sj7x+333IkeZWwoORVEqzIitGt8RqXKPy1dh5jmx38HwPvfJQ7zg1Fx2gL
PL4i1TGpyvF0uoY9GSkrP0tNN67vOPpzIFrw1nJ3xotxlvzURFZJB1rYBBGITmDbbTHt4bBg+voD
gWNGgM8oulR3xipzsyC3sTscx5w6oTro7uEmRhLJZ4tv4BqYtt9phjRtLl6AZVxoiZtVId7APtzv
9mLS3uCspAWq5txnPw2q7eYGYu14mkKiansTC85W3+jg0ASEp51Y1zmqXD9v6dCOLVFHbYaXzft9
+I8uxT+ZKqG8pg5ArkqgEvpVK7jSIZiHxR9IBYsBJIyRIV/Kg6T/DPZ7ttSTsbNeTLc7rShtGTRL
+Bc0/lutwyjbfK9ESfQ16uilZTVeV+GTgTsn+knZ3ob1wQPxn+iEZ5jjWBddoKQynY8CaQonSOS2
uDJjyhyBYrrxxLNcX/fyvE/Fnkhzhbdjb/Ve/dSAmIGnPl0+CQjdtY3I7W5Rhq2N4/LN3etmgWCD
iAwzgY0IUQf7Kvsj4qiQwD56xe/YJzR5we8ruTJDoA0ItMkISum3X2wCEhC3dvfXCBqxsoluSH6q
J8mXnW5gai/FSxFDVtejiPY5R41JMYu+V3MkY/HqsgJfmnHmArT1eauKhrI9wkgJXTiBvhusjh/X
dN/oco8HfdMiVV+ZsqsLcDGi8G8YbPMbutWq70aa0tuXJh6FeU+MhA0jYtfbS8kajb3sf/B+f+ih
6Tng4nwcV4au9DMk0SBbGo2UxTBEU5EQw36AGNdQijG2PkOQURroM43XggzhUoxSQ0DsogzedQtW
3/kN/aHPAdk0Pr5yjrV3eUB4I0fvZiwSA6uFgg7Muf/Cf/hyaY2GUCjSixyTBVtnXPexLF4qDv0p
lMWwdiROeR+MJZ4fTyH2aj4/CYyZfBdwXpdy8cDLDUq1KfUVEcgzRrvyYez54RSqtyuO/RD4eVBb
QrLZHbDoHwT+WJfE0GwwR4JJUloqM7TeQ2s5UOcKbJ2I1kuiOVmfMpetYXxwjaA9QDv9GOCONGuP
HOEx8ihZ+o5pkBHQAViV6/TbWpR7Q2Xqx9AUgJXwKY+rq5pfRL8ATGp+7mUJJ3x7lIuLxoH2jQ0s
vrDpq9aNaLpekrbEti28J2DxJjwn2nQS1VahR0FxnnO0FUg9m9nITymTmknUYHwcnLL/Tz6J0xSM
qFF2NR+tfOSPtHsVyJDq7K2t2Stdtv9UZiEzsL9dDbh6fuIct24N8aqUonCQI8o2PxAOLZhMVxOl
l4dUYq9eG7vds7ivhhdJT59lBnAjgH6Dyk3loDLrNv7xfBknX/bJYoYCEQ1tm9EEJYdSbxGiF9qH
em5fIkxywvuayrugUodGlfn2D5OaLNAvmzvgkd5FcNzUlcmTO81KVNeB6pacorQn2MunEggGSmME
e4kVdINwwBgXtkBvyDM/qZgdSdevO+cYd5hFPzSEc6WpBPlsEG/nzi6Z6rhzuPdREkWoLI0fdzJH
qVAQPU7E0Tupn+djY69SkLM5vO7LKylzyMS0X0xYOeGzzOxdNvYDtvlRBZTBs1K/uumjL5WJDpiZ
qLxZxDfTEFEh2//eL6qAajY9p3fis5Xtd3SK5PdJjl1JoADFiM7OkDrtnAAlKAw4BbC3ny9MEqVq
38yyWIwZpgmcf9cIvVvrP5lST07aSNX51v3+zSj4uQztJzlxuMzFqqTX01Q9qhDoWVD7y69zzrhv
/tVRxKYvM9o6Nv18ronh183mXv/VpPCcjnG63fqws+rHc7GpPuN0SJf2fDqLSSYQyyf8DEmca3a2
7nb8ohITX0aQ6KNXj9bQ2x1lQGywkNVllEAklOWcVjyCcXvdKzUz4A6jtkEOKm+UIa1CWGAMob7n
Fkp22c/I5Ozz/aFdo3SBT/5RJrug5FIhQ7juJM2oguynzXz0jEApcE1+CLmTVrrzfcdFuD20qT/D
SudKEV9Q921zFRKyS6tJA6pC14piRzvRJe7QM89vBYftxLNotzuYgXMMwvUYnyme2rk3sMcXN0Wb
9C6lgbCgdDx0gR75WbcdVgjzBu7yctclHfOqgh3cHeOYo8X//rG+LyoeGLIYAdLgoT7B0tN8hcrJ
opnm+kjasdpyBIiCnPwaU62AkEfKRP6+5wOBo8B/1D5lZJenU1Rf1VEBouVStRwcvQRgfj52LIUJ
YQfjn7t8i/lgJZfqLwQ9IMB1I6XirtsMB3qG3BPaK87r6Vf1lkI4zaDQO6yWcxCYqvTZcoIAq6HE
+Zrxe2EEups0IEG9urr6NMES4MlSdJlV1Nzd8Hig18vhjbWhB94+vg2/6i0BpYdYXImCbvc7PxrC
W3zCXj7s01Bdyr/mhy4CJq4ePFfztOY9xi8nsMl/Z9yQBvE0Vp6vDARf4r5pzY5bpvY5Wyn6z1qa
gOgMelYzUbEBuT4TVkS/icvkUsoqwC6MJ9ZZGtjgocToMQY1InJJH4Z7673jlsPKjRl8gPOWGD0J
a8M7tl+wXeu6XieQYEkKocuEFyhJPASAS506S43e+SZp7LXEQUS/o/xwRZ25M2dzclnu5KVIerh3
t1+xcVmy5lNXDpcH/tX6YLVLHsMGYfdODhp/3raGpOhDrLmgjDzpuwxEVrlfZqz7QaRHj6qENEKr
0NNomn0IJvbmGOkPZIyg0eBad2voKFAkDL0GAt+1kmmiLrBcKG36Pa56G/n+rw2H51elrVAzxieU
5ZdN9cxcWdA+gBtnOLteKZ+O5l/YPPz96M248snalPrOGypBbNG5Z7y4KEKR4SutYD5SMJFS5fmP
RZUG0rnQWXKrO63QSL92qg1gl17yQ+0hDka0WTSmUdUQ5XqrgEoFR8NICsMFS06D+Hg5AqLc9iNC
6DI+syfp5FoCBag6bva+om0dA+mE13AkUTc2VpefpMD8FehvnSMsRv3SrEn/nJPsA0vOszgBLr4Y
2JmJoe4OIqbIHXspQtlt5Om5pBdpB1olF4I6bF094VKvdBS1gYYdHvlHhE9vfAN4wMEclBnDiU1G
v5w4cfSxVy0cP7Fe8ze4xy4/OSff3hp5WoUaXkgcirjFSpzl2PiBYNOmiUIwr5QJZZn27jxVAu41
Cfn7ZQUG8SSjLyyMMsFCaTTpsL9AltxQx+SfyRx53VEHjorT0kr+DBRar2W5EgDrfU9EqrS3Zncg
jbSksj6nIzCTQmm4RvmPbFx3glwUWvXcbaLNvK9NRsfFtn8uGx5YUqfSfd97vYDcgFrIfFUGAFYy
BO8eB/jxveF1IczkmZnM35EajMGAdQZOunjLw+BYyAGmIAYiRVtToo1oreI4f7F08rkVH0QXD8vG
pSUBG+zGDyX0hCGU1NdoG8jhv7Qpv4TYCVb/q/li+3oc4jXchpc2bcigh4NhBuv+iE4CsW+Gu9Y2
e1xHVppA/MQ+pqg8KTrc/JMXvnH0NuUlHfiHRWl3RrLvnQ+YCdwyiwbeloB0sO12Wg876vn18Oal
JX/tvEDI9f/soRnJC3NHsGts0mKF96E/PsaXlvBx5FHg6tGTv2LdCzg2ifiwfAP7OOSSh5Gegsd4
9Jli6CQ3DU89STxtkUEwwHgIGhE9+typbzBcswuLU8HrJadU0tV8pslu0YnqotwXlstRWwy9aZSb
SPOKRNWtq9oUh4DpQgptbh7QOPKD68jYxWQhnF4fogb+O0vg2CaJl+eG4sXEoE94z35uALBujHqU
vEeCzjx9P27QD1oWdJJVVxBM/dDm8mJTc5MDxHMu9Db4H+bZ5hbetg8Y8E3LihPk87ZnZ3wQnlR3
cBtCTZ7zb1pJUIKwWf9ZFsRmA3FHD1CjPNrCgDRBUez0sKx7bvyIWH/5Av5pNv3m6y1SILj4Gv4j
om4QGkLe/aviOzxoiU89eSokSfBGlrkBXEbaLYWw94JGytIo3Ca1XGp8j55UlZttAWlldVbNbK8W
ltlPRf9XNFvusGNvmLw4k6PtRl0dameDOLuol0LLIwjvgPral+jPCYWbg3W8VNYzaF0mmeSrlmId
UbBcov2KE05dwnjIdr2ybfkH5tQ+04+Z+iVMEQRzZGTkoKW8RNho1lXrl5WbXuQDkkLQEbp9o1bc
3sMdeXkCxKM0Slx136WV2YTkxoMEQPwIDQoBBMopSaobgSSGvVTnJSivjp1lOSzh2XAGnasabPcc
Z6UY9Wz+vBPOi6+nr3sGhEyYqyAZyGJVMZWC4zuYfTzK4BHq/RvMwrmDIUhwTxgSyi7WDA+hVuBz
7Za6H81YQ+enDSiUPIEoH3t0kRaibz6Aberx0OQ5ZHtxHKFgXtZnrovWNR9JxM2o8o9KuDjJQO4s
+KTGeSnw36tBFx+PnBeDOWAi1WYyo21J7WHB/aI8vcZ9W4FuNPFh8yUVATeuyVkc2iN4UxHB9AwC
+botKvtY7zks8JGsbYSzxoH4t0v8pwbyDB/kJjoQzeie9CswcKJLs5hViewJnRg3XZNDySp22w/5
RXEYY9uEqIg6XC0OxWVjaxtxwXg/SK/L5sVrkhu+MniAQDes9STAxR1ZFhGnyc9W81Bu0LwTkrae
FN8WClMMpsl1NQDw/9SttKUzUxLJnPM5X3cWNPqdm5RKFlmCe7MukiwJ/PeQI4gSqJss//v9QeVo
NOZmvXeoDXn42V50QF4a9r8duVaqGn7RxP4VnAMko0UuRDC1v8kDhSuBAc0lSAr10Ju23en/xCKL
XlNOjhk0tcsk4J2QZ6wDaa+BwVEcE2y4CYuX62xn6XwsqcJjgbdGLw7iNVot61fA1/D/UKH5s34D
j26uvlkTpd46PT6W+mnF91N2UAgSC9KInGsTzsCsT23td+bX1wQdE515fb0taer8ltn6rk8hCq5T
Fhp9gXmyfeaaJ0XoLY2n0dXsSGUsRd9zZPayhMFWrJdi4KdmVUw+k24NQkFLsrNTYs/rhv2LBzE1
CPzOT5kUMu7cw8xukjtKzhvWIJMH0zvjlhMnHgvbvXBpI1mWRcMOcoQJHLFs0IYB9fyBrC6kvJUv
S8SPNf/LRKDI/vh+vPAu5tF0PuFM8TdQEdojl8j2fm4fUjk8ofFYVbv9W4+BMcLA76d/ki3zJnDM
2RmSXzd913cyk4Xa9R2SzapmN9m4ydnCU285JS6RVFJrWmv8+0rTriWjfOLeB8Bsj71Lj/s2Wq0S
g+QOkRB8ISfgRGqeee3m++cgKu9ht2t7J+I6bX0GrYpIv3OHQBw67eJ9cBfBjvuReIkLe2Nerv6r
i1pakOgRYaoUmPaamqijh2aEbW3C7smLOpc/qGArSPoPFPKqJw8GeOEC0tzWCfdy70xAg5UgGOz0
gnHbOSVWaOUCmeROLEbXEiXrmXIt23a7C3NctI/k8dNISHBNk4d5CnX58iwFnyBzTythrxai4NcE
A7XSz7tDdg2GBSt0l1f450AY8EgVTCTK5yvVO10242ib8yVAF1EOukiHhTcvR+nKPV+rFBibgk+P
1qxdCyhqxy/2KQU/Z2q7KYzOkfn3BkT0IY7LBhibslhTpjqxOZD8ygbyvbYXni2Iz9KmIag/0i/e
RAaNBPR1WZqtS8OW1q1AnYj0RIAkjWqsRrKK1NbuzGGaQ1F9WfCXjOxngke+5CKM2p5tJRFSKDF7
522iiPaywJ24H/sb1Omx/cPJ9fmtaRqdPtyg/TcnVRRz9jIK40AJ297t5nyCrpB8tmFe674Uy2tx
gbk5fYIe5KarUJr69VyIC2v93+hyUAAsVupQ8wAOfWw7wHGiR0N7FaqSPPkzAvlJ3t3Q7zje4xlG
0is31juT0Z8LbWHu6MAHzApmThyTYzkOdmC75pl7IiPSxNIfVOiCnSn5pFC2pQZ9/XkMG/ccCKHQ
KAiHaA5T17QGBFt6ulEeppXSJJg9OBIXizt8lXtnUec0spEgzE1HQ3TqxeM8+iR8ua4PmZ+JOvxG
4JO/Oop4bxCcJu2HbybtghEVwO1qKLgWcEPOQn6yHz2mGKCOMZbwvPSm2QlKnL8KAf5PYy7ozpRv
QUcRqLMHaDpOLkx5r0xpQR6S/5lwndzV1gniXOvNCR64JKkvYwMtSsERCOH4TOKMInFu5rf0gHpH
L2KuIxVrUk/wO41X6IDz8BF1k0NYKGXcs7j4F8vTCRxDF6/tB85UsvXGiH05rFxh5Ot24YVxdwh3
yxFE4voWwNknEEm1oBxHGRBNFgUfqsdlhRrnjYMWDPQndzDV9bFjMGLbjrRYGSV8WRDvnd2WlXav
jfAPPkGxDua91YtC6urHNrkRVDGzO5zCPvc7L4K59BpLnyKsDvWw3yp+X20ZKmGjIk6aoAf8igch
RLQkWPv/Lzno/ewyHozGB0Dhxc57JTqFDBJqPLQ9aWz20QTdZNCMRwH0bjrE5daJecwaam8mdCVe
DbjN1g9GZUjY07nGhWYMZM0BRy1P5zPJqXTmhYDgQtArFaDQC/22KbuKg6eXC5kGqtYy+f9qLaGi
eGMJiYE2YmQ9WHC7Vj2JvDtWengCZrpuekxUkvNflMldvfxh2xNUwe6Pktb0vkv1/txz5afaSN+Q
qnCBaLr8Gdd5i3Hjr+7Q2vkBs6PDeyrYKshqe7wfJ71eOl9ceRbCF6VxDUHaJLUZhb1NnT/9XhEX
qdIkywGblQwjbpFUNj5MNZjAbLaK0RZJEUd3K/83Mvgcx6ZT9Cluy+5KbRUaFaQQZH/9036A7jeR
EqYhY2JkMxoGbeDy72TwPvzpviMzEwaDlzyLLspVFzxeYYkzo32xOtQEdDYdQFAHzQCM0c5Y5Uir
SyrsIIdHknPBAn7zKZarYKizMT8+15E1Poj8XuXj0Q+wOdwAKRZEIs27EDiaAsSBnA9ayat4LgyM
pEhOknBrSQPQha2apSAfsYuB9VOvFCoyNr5i9LbhQMyDFdRQrcAC0AUzP8UMXOVeAqKiof2oBOgh
YAV0n+n1vYAI0yAjgoKpngPrXoTFGyzabAogSAVyeyC4yZbJez97xxp+xOHVMPGrdVlAjdSukm4m
Qd6gKvdVTaYfOoKtLMF3Flqr8VM2Q3EyQ+KY2YGPwOUSqrSZDfAEFRUnNhxztcMN0nHmYUnm1D37
YFz4sqvPPN9xUcQO/i5A41zblyugqe3EbODJHcZytvJziDPQQdwO4JrhQBS5VrgNxCjDivpyhpUW
0cUzpmJk2n/gE53HyXX17q4tETCik8/3O2eQ13wCCG+o5TckRAUfXjqd4ML17hwuWWPKjqnlwBqZ
eRmlGV56ArmmELzQ9jLZk/8W2cEKB7dRP1LE6+gl8724jJ80psA5lWkrhT8HdTwhHoBytjTGE+/y
alaVJMJnEI1NwWN77Xoc0g1swPpZHLvERzyA7HBSW+Eau/gFn83NsJ44NDLWf0Xep/lLSYN9Rejv
4+T6jfKk4tkw/RGk2YbU+nZEVP3YvrL1T/a7B6eYL+xjOlnreT9YFgyyyuOeOXdqmbc8pAYenBfN
wr9lHlQZ8u4YbpyurvqfV+UG3/YdTbndFZJUZ89+stats3o6xkQptLRs9ufbv3aDHlxqFTyB5UxY
iDqdWmbGcN81bphW+EP+/BdVAOQNTSHoCgsEAb7xwprCsteNR3JxorNrId95VlUjUISQfcT7EDrp
BbDLih8cI/nJi4XDI/B93KHX9pij5jj6776Tfry6wc5nep0FyNlibec4XflIAYp0YwJUP/Gh/WEZ
06NhfJg051RVSWYofHpMEc6qdSVHGlL48HTHjkiH5UX2vophSIow6ti/rmJgNwF1AyLB6roun25X
4oVuRxEDU61/QvBir/DrAR2Ah7PffsV7Dou1nqgiS/1dV45Tt2P07rq6+nvPV/bHgW94fpztPMBI
G1JDFskSaGcSsbDlrORIFKMN9ottQ4+0YYrL/0yw1kRqOP5e5cEC05c0F69vQ2uzoSrERArBlRgq
TsXiimC6vDPzRodvs6THPnNte/Af7NX3z/x28XhtYd9JaHV2KkIS6tPh0lP5uPEvzkcoA5OP388P
I3ezCKttKKD0kCJYZ2x42P4Jdb7c2uP7X7U/nmP/eRvcgI3bR2BZNu4Dh+R0rZToswpi7sbosCx9
J5zMwSwDwedTYELNCvz2EmIEpQKd36grnANdW0+YWT86ynMF7l22WE5IToPTumACwqfDLM8EmgBt
3kMXmFLgFUnYZQ931FQvs6WUzgoCOaygRtew0o78SQUpq+BqE4B2BqQDWu5yOdyQsTH6srd+CUyo
txk5r+dOVYki6z+yXklQ7U//65DbVC3YtDBofN6Bheg6VfUcNYzKEiP2VTFInW5SKHxpjd6lngCw
QE9ZqugCNwznqSTBfucWbepQu5LZZTG2RBeqAaJIKqHNtvR9+hUspFrt/lW4wQhZO4Y6WJdls1Cq
mcu07oa1QKigXN3jawsKsfzjmUyOc8jhumwkd4IXg+2s2EnIluzXrvGuA0qtNiCocgWmy3JQkdlp
j19yW28hi13yEqpycj4QkjQnr57U8TEMTrKdFNyifqyc5QhSeJi2eYvuNCELaJ5cL85bbPxmvzxh
k8g6U9MNwoWoZOTek72tb02NuQY0x9DTK269xESMt4soHLsl17OtX80r6ibx/za3hEG8VLT16gUJ
SeUNW6OSP/YMxV3Azfae8ChundKF99//sNEhnaloHUZcJ4TvfXMDbnuoJRG9DIjkGrB8ZJ5xDvZZ
YwTZiXBxenDxi4iKNzzh2IoBvPdAI60oHIUvvWdtXghx+K6eUrJhKC9FRdSyS0x+MCiF/cJ9jeSz
RgKoGF7uZsXhzv/aQynfojKCutbPCcEockpxhkWDGd3s67DmQFoQiRen3JRqNy6d5Io5ZBjHiO8M
caTQl/bbiOlyF6MRy0dTMlUnQNvGA0KwWMdB+ab0k+Z6w9q6dn+jioECOayszhL7YxgexxgVUDR0
CF4wjnn2EkvlvC/RIqYV4rR67Wj/KEVl/P5TK1Vel+j6QXcZdNgTuS59cnVAd1VQVU7BOcmhNZyC
O3wPi1N+CISVR9zqhCcRwX5w90bEbylgWN2bSXIzOdy/iPKfWZahJv2FQBX8uUEuNERxK/cuOeul
c8piY6okZeh4mS0dzJ3tnUBBmI58R7jiAzSx3y4JctCYUrxKalZeGKRG2Rm9w1G3m7PnzwyCnbY1
SiIlcoWyndzJuTdPCmIUjjjnRwNpGFkUj++cplHXLLmK24O0lSpl7eJ+wOTMkYYYWW/pl5wvLRIq
BHI4cyf3UhIZq7dPkakSH04iH5WwD+r/3W8/fU3f/2YDcYl2fApo5jTDxvoi3BGW3Totmpte+HFC
aGdHZ1eezoaxXbF7f2zhCQ8oiuAmUlIWYcmNzTIWUYefOqvteEwtH8uGdTMKnGHAZKlmxYMc8opw
8I5Cmp6JCC30JrlmGfCnhxQK5uaCsknnqDmg0duGHHkag5JgO/onmzotWNJmh5JazRebWn2P8Mjm
n1MMdtXo4EdkbMuRKWiZz8Mj3LarzNGY5eCZvXy6EBKWM7omFmmFhiZvHr/Etdx3e5veoZ8YWVUb
5ver8HDtZV/LT7V4m+8qLowtlTBBLImxG8P0GQQ7beWJnU/i/kaYwrACsdyp8jdilZ7ABtErh71v
tN7EPkwgJT4Os6znYoro0/oxfAcSWNrSrEytylzmK/mAPS73yKAeE+eB0q3HPZgt3drE+ASe4Md5
KGlFK+pT7kfjOe9nNf5+PwMtLfvpUbVOWkS4/oSxv7noeaK8wxcWAaUczMSu34QYF7BFfIgJxc8T
gCcIylPSN3TSBo/M168gAva8jWjx+Z7TyFwcRMl3xWvqk8QDol6nwO8LL1zJKcmZ7KfUWPsQTuvk
FFTVoWd8iJkjhzV5mI7758aplmq+cTWFh6rOd2Ugl4g7qF6cZ9gJkAnXmSSias+V8eJCDiBvf6pK
ohANe5/K0OChC+GVmalbGEW4WXJnpYbfLvUjscfDfJPY5q4nhdgKp+xxY5F4b8ZoONGGATCj30bI
VDOgGK4cpLeffy5vcxhmpwcDA1EfNgwXlfCADamQihzCHarmd+3Ob40Trl6ee0S0gB8nK2hByWYF
5OphxtBrY0NtVjAQ+bOLwNThIaEu+euW22rjBqqAdZGh3CYIu77j7L0SfAYmadZmmW+aR2hsWcGZ
canW5DByoqskB9MX7MyicnNF+cpoQoai6PM/+P5GjYGe9G0ROLZQuRvrlD+8/hR8EcWK8kzZUp4b
o+VOIze4cPIcWtgLAfdcs70TL9wFM5hhnuS5mCqA7l1th731AWGKCYZ6cCDnrGHJTCy9VtMRl9GI
XuU07RXkvX6vqhrXPKtVfcqFrtC5s7etCNFREZqsuZgNj+fxdnk+FX+0lDJ6GlrNBZ1wuGO/BOyE
PQ4YyqOZRffWT+QOg1HgWx67lMvteXhgk3h8wCUTeVO2KEJQRwD6yCncLpXXsxnljYjEO+dZbPRb
3QBkNJt0UI1UnsSHuT/2gLY0BQ3yKZJHUujvopR0y17p/dCSclTDqzpSxZZtStPLPjaj1ZE9jDlu
oQ0bLU0FpuK4xpoVhJcQ/7PlV2HfvjHxvpVoPcffamKLvImsZtBcVrFYr/KvyWufMa5Z8pxJazhp
DQC7fMCNWhfmHEVIxIfD04lBbhkQTsOJ4wawHQ2zC3TA38+KlFrWIA6MpbcZBtFWpapjJYBIy0tR
MNZuUnaB8wy4G/zLQgYjkn399WZkaGAsGL0UqXb79AUP7UGjrd7pooJ0ELdBgGfF5/v/0GUOrPWK
u9cWb6jfTkTv6LUlqn1HV05ckWkZ5VX3Rm54CS0924zFLkWeY28LROSWNf8ghR2N6HhwBy9MN79X
iEcQCfU2m+L5qq1eu+xBkZ14o9+Ccf+Tw2t/zCGWfUg3v5KVp87u2IlYm5/5l3LbghFNVUIi41w1
2NwfsuiVhsnnJj/2lJBwX4CySZR2J5aRpxKrsj2crmSxzFNJ+3wsTwwZ02kue72CyKMEUuwTlnvX
OswHBBSY5gZUq2Ak5bRVJn23gwlf7CCUInyp4qZqlzt2yjccOUNv7NDNzexVCZlUOTCH3yhiU63w
H2Um2VFn0m54y5uRordYK4tmxJ0bggiBEYIocNn/im968PtBoskIPqK6cuxMfpmFNnaaFKok7pet
OLCUXb9h8SbRM+CaLJHhS1do9el1pbTUvYr6J1cv5OGAobuuBFNv8txxaYTgbBjafpH7u5ZGUsZL
iQ682lUMgFV6WUVk/gwWVRqtrcPkTnYzd0qlp/aBzEjIz+MZKzdaKS0e0DCFXaCyt23ZR1xhUKDB
QS91e0uEpVE3FCkQmj0Smibsf/g7sPIWdtSmIMEy1KlzXZB3EptVOJnMpq9KuGW5AWQpdHI01Htn
8kM23oXtXrDNleIVvIdUUpKDO4iSye3UnLodBb+MyYROk5GBh2+5rbW/irjBfVCm7gOgaxF2ejjP
grl6o8Z3C/fytZe/ahWOaDq+3KJz+U8JZ1430ZLFhMTBSdQyRNpBwnEVSasSBTF1W/MFcatkrcMP
+eJgJGk3j2Ulqph0A/ar1bAEJW14IfP2DkYls454Hl6N5Pbxfr/bYG0kXuRbloUKgySITtuVQK0x
QAX5MEfWfhPx6jXcUn+fFSVExYzSCmEZx9U/DKN565stHBmulVR5Xgtt0b+Tsl46fmibys7aDU3D
lc8wjyHA+/VhwZayIlrB5p6t1P0aW7ydgOP26eph8BsYMJANTIXFgdLFKE6Iuw0o1hE2a5MZ+E5a
hpekNePWZ0hPkXTCuOoIhlpzngCOaAa1eny8CFPWtBb/SU9j3QByMvBMBmujmVk3bUz5KlPDovbx
HEV6K9cDRFhl0EF+R9uw8+4amnpdep6NXXfrw1giTWFYeTBClsiFJNXR2x0avQ2Z8fsEGkeK/7kq
2lbCFiRz6EIBfgUnhoT9dyHEA1fQsxzGoq9VfSjawkglTicqgzD59fNgkDhUm8tn30PR/WnedvD0
ONDcwar0QApxl7g1y2+q5weHlGgruDYOpqS375dJyN8aYiOshWux4YffttNZ0w+V2VzIho9mTFnj
17/3ofpvNadbjh0T8qC04x0EMEaSwxd2dIYnOqmmzUbi/xs1adQFcboPkTafPsvMelHhQ9BqLG7r
8OajwglqtHCjGZgJCEK8rIK1xojOHNrt2ZaMZJQyUyskPFzz/EL5wwKaDhCsvDSuGddZXigy60yi
ilBa3fJIjwu3s8AiP2ISyA1we5/qi9Dk2mybFnZo+9LnFWeqgjQiAz1+OFJkIGACBDSTS3RL+i/E
RfaCQI8af1eo0mitEuFR2mLavPvEdmQ4TMDfXLWr5Sgdh44i1Q0NUnw96Sa3QuNbYCNl9pHwS7Wj
bofXwGVgGx0FUuIz4JQBY/TAQJJecgN5pVyeySItQglVbAaftp+F/rylWy7g2AEXN+I9MMlYslRW
UIMPoFEIP/ghsksJg91EuDppEVTuKM2wXzU76jetd6HQYp7xCmcq1SRkSdMkoAqbihf5KurgGh4k
iyIk252mWBcZO960pQmYzML86g3X0wUoZqqOcl6+IY7BjORyiESzUOLyEzHw15SQSyJsc7IC2AHu
ehMQ4TESn9HImDb5NlOtJdkziSJWaFjq/OAbzGw1Kr0IssSpAb5IFYXd3f4rJxrDV4oDa7OZc0uQ
oP0C4dx2A5FCc80SSo5FVoI22+m2cPm+6VL9YPUsmeH+3fhHK63EriRECy7CLsnXGWJv5FrQLG1q
VthSna28bfXjOOyxsJ846x/lrKp7byT2+gUX3oPMH4l6jDZ7f08+KlNxmHafxokmilf2OMmkDOqw
uuLPiKRx2X4RrTTqkkXoiWW4fa9BnFiuYkF8Xhv48qGQTROd9K3lEXnxHhwsRTjdrifZPZy2hdny
Mq3qPD1r7OTH/uxvbIarAsgr29YXZ+GRNYECSM/8wxKrVF91UR6jXa2Wf3ULlF4O32hxNL3lFTxI
XBV4HFahp5pR/QRAYU5U/Yxkv+UZx6TkAjLGgAumF2IxybjPTPlAOC2NnuPgMehsv1WXiAjR1nir
0iPS4bLwaSYpdjGTw/yVm6qihQmcxJFcTqromlfDBu1j76DWi+WsS/St+Ez793mMX4mUu3Ux9MhS
wiMHZFqbORuVkSv6ZOd672rchQSNdTFZWoyt+Ra+Zze9L3gwKRWmvRmGiu/5HFyDZmq7C8YD1qlv
PNi7UJWxoEzXW+BOHvaGLnJk3BZ40Cc9BIAOjKH+wdlbQ0WpEF0Bjgp6c+dxC8AxHp5f9Q6eXSjK
4p6Y0Z4NvjE/z97ogcVYQHtHoXaF9lX88jIeYMo39DVPyIDs4qAN0vS/JYAsW9VBV/TpVkIKGFrh
nbueVkYu8ENHAioSkrLeOcjPqv4DJogwaajJv3msaRTn74VzJEiFgJlsWy52fsYyhKLcrj+HJX75
ltKsIyZvNk18O0nZ6Vp53bxLM99qV3yIRjJdTUt2v8C5U9uk4dWUnJh6/LjpellKYR/H40VJghK/
91EklWbhlGhd/28lO6jvFwsHjw5QmA2EnOzfkhSwKn9aZBAMzhziWKzj6am8uJxYs3PAzqIpTctI
LSPyAbeFXwBRrgQgcMftqKCF5q17K4ISDpqo0ZX1Ok+t4Shbze9HoghOR1W3lrclpf5tI1o2UxZu
m9AY0E1chPzZGuUV0WyTg3k5ql2Fl3MqYA38odsz3LTy3JCtgGN21fTW29avGbrstixy+ROBg4AW
/NVDEhSwjXp3MqIu9sa1mzhWWLTHAAOF0SWN+1mawDDGhnyImbWHvKsL+LTu56bEmHfj3dy5eIoG
goazcMcj0Yp62+UHVK+YecIkJ5R0qqe831sQ+gjCNiYJVad70wEuu+417NO0qbE08rEs1M6bdZL3
U914bOVhiK687Qh1cSmAjbcME0sYEDjspQo13BzWvQpIvr7vcGT3BR6Gvn3/3SFtfHuAd5J40IPu
J8GWS4HDJUfrH6vRD4nWzViP1z2IdVtFGhm0f6/+DQnZ6MkpdRKP1mFD6OksInV6dYTvIGlfvdjZ
NU3yovy+yUIVZsVHXYZfP56tW5fexBZjgcCEBAmUbK8pcZ8h+17tjV8WRy2yWNBVUUdVEXuKFTSl
6f+1Hedt3PPyIO50jShd1R56era+6Xgtr4UTYEGUc1vnSefXh423fF5RPMFeVVrrQZrm5aEgH20t
L5rUBu5t392pZS5J/IxQ9qjEVHm7jdUD/VoJqPMEWEetCnHNdubjU8CVWeVQR/QeSgWFyH3lzk3W
uyO6Q2mRnvPCc3vWsSRWfORko6XdgrHKpZ5cvZ3wjgg/KgqaCmZWgQtLoCdqVAlwKDVWmmXsy7sp
6pB+Bb85o2w4mDek8WtOGxTplbsCenjZaza/YECr7TmIS+xSPA0k7/Uo8jKyagp8jj7Tx3Hk1+n/
UppAoXgsXmEN6gKnu/l7jRpQUgih/MCL7xprJt1Re4Fwb1cl3G+OCEekmvgFv4OI28ORzkqo5l+R
IBHnttEdoXRN/Vv2QzxNFGEoauKqI/A9pBzAq9v8CIYWRDSDIPZK2GJZ1VZGFNaqSbvPHm/MEjXH
TBlwmok/uiDF5lOR/fEhqd7uHYAFgCubdLvbEJmv+SUDVyRFvp0gTwoCdKqXzsNteExo2HmpdKdU
TLee6uqBw84m5bWNKnM3uHuiTVtploLZzvWOgFLtmn0w9kn2Ga9sDugGEz9ndao2o+rRl20GZive
A+jgxltzz0fGTlpzmxRDm/gZhIWPiRSpbapDJdsRPOqBTuc/H2tdo3RMr4S6yql1SwP5AWic4XaR
Wc1wHxotKDka5Y+YlTpg3mbtQjiO3svDaytWjmpmCep+GDOsordRzokrGpMVeZTSaEgkmkcrpLf2
LbJfV/YTBbzSSg3JY78WT3KfjqkCjbIj4YjvBfbz9R7dzzX5fGML5dODPTKLBpDC8lETPTC7ovmq
reTUhWLhYPn0dTeRvCWpp3mukle2K0tkUMdNC5fmVQ7fFNypIfPaKj1FxtKlHv4qeH3KCIRG3Gi2
nUoquP5QekSO07LRYc8pFaVmLirpPYuST6fANCVhy02v/I/cGUm0wq6ftd9HAMaQcYhIVh9zX9Ob
XmJU1szwjUak9SWDAH0F8g5FP9xDlAj73wh1mkM195cuEAGWaVqhbdhOXbRJElhqdXp61G3Ublsl
7Of3xZ0RzC+LkD6gyVwF+Qt3GzIzs1Sd2pNrtJSXO+RtVyuG39e/fvGSmwY66XW+QgVpQGcrji8u
GQvAHJIcpl0CRDbVJ5JskQRWrVVaYC+i4MERP4ZkiVUdG9cAeIIr9BKOdR90JG2pDOTwjzaETllO
Jr9xV82gewlN6nNsNv4wieUNnw3kikDbYkvmj6zvQzRwVzhx71hNLmRCZo0/d8gZeWBtrMTTCbbJ
JqIRWHUO+0qLGF94gJDeMhpvY3Ox5Y4G//Eby+VSrERIh8aIUK2nDRbsUQGg+9rgYgfQOE76Hb5j
Tlz+jAfu9+P4kgK27E77vzDexoPEiY1y7jE99miBwutGdUV1W4x4QvP+aSX9oV2jWPP2771ZTnai
OrIrkXYCIEnFdJnCX7rFHAgp8cge4MfHzI3+tlkHE3xLeQ8jGV+5wXyCzXKm/pEwcfIoS4sKPktT
J+CAXKqjOpVo7GfBEQbOu6I7iQKK2fMMORdFplJ8Eghy2ginvRn6oyYHrTrc94H3dA6HR4/ReP0W
gEtot/5Dnox8D7PkCFHoBfpWhS3hJwcOfKRL1UpGdzRNAdzk+/GQS84hfspM2jHXEVro3QGzTQTX
yH9SOrtvU1k/qdafPuCED5yn6srOoFFVaxQxFCLA9JUISiDlAo0DtAinMzozyBWAUqdZQNVsUiNV
5+W8rl7YH7wWLkBqngRMVIHw+E/gCCofBzRSX1Q/9LLrOYL6AYVMVq9aTd3SqD/cA9DPs6EZ9P1R
BJhA69PdkGwmRQNCUUU/Bm31HzgTKrKdl1yNLXB/Uj7SiDInZMea7oW24956wHJXuhSf+cCkpaCG
r8+VuoMwWpCW2dKMr/5YVw5BGsPovfxfFaeuywYUFRV6XosqSIbIe4hUNZ6WcB9f+BiGsrW+f3vb
BEuAai+X5bmDnqC94b4HlLLNJBpBWp0x1H6C0FS3tEHgi5XPmXsnKI8i+tWnAZWwkj2v98Ata8i+
vbBqKsjAljd2FrLsREa3cq8nnWVRCFW9uD7JjdekTEsP57ks8EVMcVm7Bi1RDWkOn4s3mw67gOnE
KF+BPS3zjRTtS+Yi8TTUdFf9AGvtQX5D2iOvCY2xLr/zpkrmaQdSRiHkNJzkke7BZtNrPjDK/Dy/
UzFNdoIiHX9HwY0vn81d8a3lO6BA1NA5rPigBVuhNKrAUA2OOvrhLcLod4ln8gZT+yHqhdNLzJ24
3GwW7qXMmtHIMR2mWUYw1Hcxv6vlsLoZ0IG6sJp1WwKz32qDLyYfiTdrDBbtpVrl5wk+vCNgew8M
5t5eikPrzRJsYyG4QTmgg4zwHweC3o7EYPuj6ca3o9E9UzSVr2WEify4qLq5pqQJkNzp+LzhLt3X
qhd1O19Q7ZhrW/mmeNX/ALoIKpXULk2u+6qcYonh4IQeXMw8v4QhadgSNn5N+pd5ipZQ2EKi3Nx0
NB5eya+jPl4wn80lJ8i9LcTBYMAZHFd4HYMKhKVtVqmzSX89LrSuYCTAUEeVT6rbFIkMg3Vpn7Ac
vux9qW3rziChKsVU08PDcMr5JNjYuiOsot8ORLtJMqw7nhv3ODi5jhBx9KMdxhSgZxNNPCiohhFr
znUVARLvxyK210eKKY6/fint8lpCGHKkIxHtOmlVbpdvXR99r1W4SzXAHITNgnabUwZfQcIf8sQG
DuzX/28CBa3HD4qCut/TbShUvpvjPK+dDX+RxK1YVB0YS7D3AHgmHSmfc8hTSTpWOPaU/5P+Vkag
w4xr9nfyWUAwFq4sdsNGxWJ73vI9MhDW0dXB3H9Hps3EmmfNElQBqSxMDC2YuN3UsFqiF/+gn8cE
s1Qeq60LH/vQnn5yMxmR4oQEi5XmwDLRjDiGJfJPRB+MLKKrEWTUyXZPSbayVH5CCw5smTJRb0qP
HA977zBifOMRTWzvkVgAM52zUDL6PdTf7BAdT298o6MyN/A4pi9b3E9HlWcooGTklOVWEsv0vMua
qYX6EHkf78MIZvr30mPXXfghZXaEEhHM5tOqTbk5yBru4Hg8E+c4ZIs7CSXgZMoMnF6pV1h2K3Lx
ukjIztA3dw1ORw3MFRiYRbBQRovOfPLdX6ptlYvwT365lOCyV0TKuiq9tPazKXXUpBJCrsZKhYRE
A5xsYtiXNzm3YkLVHFPI4pGd4Mi/Ng440HUqBj/BZMmz339/UZ/0nzWl4DXppsqECOR2sb1F7eYv
LVGMZ2842GPStoSPQqvIAXJtRAzQVBq4puYBEaOqHThdTleURvtghX9UGc8EsWXm/D7I+j+cvQa6
bT8DUhnEt4/5V/VZeEncmuh3xqLL2bHDUJEL4DiOlhPPexCXaXyA7jnRgQaPgOVUcAZLAe2ihYWz
3hKUXuabVWc3CTFGamE4CC/tQmQc7XcejTTsm9gb7HTE3U4Hg0biq8qJsnJ4bpYWLA6NSMwixsSh
pFuYLflU7rbYoNa87IKm95+guq3UYTZpe+H/5kBg8ZOE9J4YnLs0PJwk94tI12tuIoiOG21/RCSr
2bkXkMYZINmCa/saGd0kxsoLU1Y6+nDtV5A8F4WXb8q+1ve4+tbSdpq1GyfiAtSW1Gv5Xp716GwI
amiWJGjCb3xWT4upXOJFgGk6JJLTc+J+QXtU00BcpHpbpP/fI3zEiy3MylyX6Xn0fCOz/JVGwpGy
vKKd/yCwUdhno/vuqDIRi58BztCV4cEeJjPLOfpoxpCGaSPWGbcFwx9HoX93k/K8uiTOV8jo8239
1X+iq9o2pMVGxrroTOgD0u8Uoi1V/RHX9TAvcyWWrRka0kcGXS9ZPejsx//aBsRTCDvXkuvgQIed
clobFiwXwH28lzHc9OjabRFxxeqW1VtN+yO+m42RlxaCd4goUSh3L/3sfMKX8CX6GuooKuIlIJAF
QyzFCqGfiyrjVPQsNYrnJXtJRLhddk7TMvi8rpPSDscor+4EYIRWrNoYT9JCyCUsflMOHCTUD5H5
xnQ21aHmMiPpp5XPp8/N1Um8WKqpH0rq4cdpStjZoH9sbCmyfJQCbgO87JMnVaqxQRu0ZQ0Au+iZ
bU24fHVh3vK1D65myb84cMYxXYNfrPxKb9vrjcH4Mg/FdomIfg+8iQ7kRGZgX6DaR1T85YNsCJNk
gahy4mQRZmCR9oiptRcJgYqiDdWACJ468cZYipC2a6J36Y+eNJ8ezcLA290cbPA5XVwuo6U18g4Q
p46/0vWKFnc0g/LwHIEVe/wgq0kdOdURKoOBd+HewjYNRpWYdr+q6w3dpQi16jA1CTl8gP4Ptc2X
8YfMtqRP7pnpemH8j75PRXoqYYQZTZpYxMrSsPPfdTt/TJWrGzfV/My6cVgfHzWbwaEb51TsWnb1
x0+fxn1mfJTPLPdIyuBUsp5p9KTH4cUOB7QOs+p99MWVWcR9hKsGlPuPLOFEPuGyuHD/JsFgmKhK
X8Ck8/O7Voe2HAe+LUo2tsA7jh7N+HT9zEjbUU6GzBpjK1C0dLoxybiEuCXYKBCjLhpjpqQvEBlO
OReiMg/4sGQ/2naK7Fpr6V1xcWZWZN3qMfIFT0m4877dKFCfqCQqaSkL5QgqRVR96KbMKCvLA6JQ
EQA2frb9nfMdszvV9ouIZX0xWHPMoGeXN8lJTc5XPLKOwdVdqMqfE5diZCJhK35+Lo99ZEX51QGi
8FLL22cd6r4gywegtUMWRxhcMI8zdGuzcZPQ5b1H+EkTEtBaGtifKQPff24MZQ+LdAZ5Z4uIfK/S
8icBk9EUjifL6WxaRDPXdXyxUS43PV5pwFuHBTh7IFPJz3akShy2YaI0I94O0xVMn3IVOLfT3loV
ETGmJODKK5O8DYFbQzK94S6AA3iwdFwB+6ftAbbYNlYB3/zcp7+0OIJ4gEKRxdXQ6pUkIZXV7amf
FgKO/fqz3g8rwxYlHiYuSbVrUc6qFxYhQcnyQE49C7idjG9ijmTIpEbEYxwLO4MgdEjXTssTGTWJ
XDhq4lbRsXSlQqccx1EVhnA4nq3TdrzBKICxskosnFR3YmJR4XNKQOMYE/wryzH8RNgTW8KD4iXd
c3cPIATb1qiuucE8lgDzL5sWoFUeBosGIhjtVGxL5OxWgLEyKy5Jeg9KIb21mUOtEXip21AzK/rc
UIzGVJDUWnuxt3CuyD3475+GH6WhLh2GBLdZIbFwf5Or529OWFD5PcM319V/Eh/rnW/ZfUX//DeA
EZKIzFU5AZqmOdqysI9H3JOR+ZQo3AXMql0eERdo10Qhm6ZNlxC3qgnbSwcEDMq8rCJ+qNuNEUGU
HO8liHzrvvE1ZF/2DnMhPUT2Kn2IxhWp39L7NQSlDzXpuTX/YxYAHJ08njm2okmg6XaiuRtIStS1
wfz4mMDSEIlN7bA4YAxWIXbgP2ZVbaYuzbzod7tEWb7joQXuPpRNicUGy/mLtgsXqOQPZhz5gtTP
D5pD+yNJIArN3t920pSROPOwOrWnvCzQ/vxnGgXRh4FxKN9l7PXwuoepc73y1OVfv0wFUWsLqe0z
vcNqlZGv/3L7Wcpa4ahbMkrPQLRdRn19wQL7MQpvdgM4+oFJUtkCCAbisxotgtUEHgB6XYqhwD/p
aaQlnlT29ItbuEYNMT35jlkL8oee+3T44lMh8cTvYhc8yGpD9ZNYDvNdVR5TcWebWZwdmLwt1fJY
RMuCpgQT/8MCmQhdYlCg8GxTLeaBwViz3Nthkuun3aA9pgw1DRG/27lh8xmNWU1IldL4iUwwczMq
oneLHXTCvxesRZDfCvZZM7iLU5ockutErQP/E2PfpwEmA1mVzZc4yiteHTZYu/Jie+HZof9CWGIz
lVaFwAWa57bqn3Oi2toLNRjXeFIefSuvjij/ghL/rO3I5k/3YuJjeNnG9Pg2bo+zWnZBZzx+zN7V
hsYVk0SS3QIq/P8QObI0wxEgqFIlPQ3ogxtvaBiP1rAAeq9+ctnn3/TN6dgpNDTsBYss0kBgBxPN
Dv+yt41P4Sgyz/5JM7jRDOG1BLQF+zTuc93SozZUrPxBJChXmb01Pc6ty8+cjLDW+g2ruQraPbsa
/hY7WeTrqUkfTS+7tc7ZLUJpkIzLj0CFo5N5nxd9MqRjRYqlGtI3bwNW3UyNgkUjajmOBu9wdn3v
5xDgK9YZPIZicI7Bau4vVV+2ap1sPnHxt6YdProweAXbfqITS/abQN+Q3Hl4JIqRC6iTKMX0jrQP
L017iQBwqJG8qzDrUE1icRCGapMTXq5VMb1cGLGwwPcPzWGchpQdKRcGwOG1aKY1JbZBtddjQNFH
dJJlMVlN+vP73iygCs9w9fVNGWHC+oSR5gaoX3GZigwpN6QD/bLZyv7Zdg5uT/FionD5imhG7wKi
OQkf1MplEopR8+2J0UmClsS6aDHSYRn57w3Hlx3V6IbHAbBvmzTzadpRF26yzCRlbZn9wZlosOeu
kQ8lMCm1eIqI0KoAdJ4oUaCncp1uHw+E4JpTl6MCwGINYpu2T/Owpm5plkVT2UIcD5tG/YsgWgfh
zZC5sp+KznZueGoMGnrFSU3ilNc0UsBAhzbXPGr7Vn0hjikDH3eUqg5+ZsMz6QMuqnBCE8BEIOHB
PzPKsbr3MCFJx1kdGEMpy6N7Ibg/SH6XiaqYuRl8UlP5TzunG5S+J/ntd4z4+dH4RQEqEMVy+zO2
zfTpkUgOXuYvRExYXVzc22WYvNKV1+kecUCLZhHoGYnXFltNtRfXedzbE3a96mawuikHvNsyFdSQ
SARJP2RhSbSHP8tWkWI5VN4NpODXPGhl/x1vZYPr28hJUsAvqXTxF7/YWQJe3A7iMECzAGaomVyR
Gfvsjm7s56V56dTUZHZQvAOwWIrun4Vdh2mNkK7se1prZDvtoJ0pgIFYKZC0jjF0LuRLcrbvvIUS
2GsyoPVKsxOQqQXwdCYCop+oxiJDRV7XgLDPROspOqJxshVq5wQxMrNJzkCMx1OYXim01xEKqAuU
VBzDfmjm36oAbIAezf2imfvW2yOZ4Pn7ovUuuJrng8myjB59JP5QvUsQBWnvMUf3z571YZvPDh26
ddBc30YlVFcXnaaB62IRL52l3V9dIVfiFjBc6+h3zIavADQUh/IroUBbjlII1EMRoza4SKGtEW31
fPL8eVULJFchktM/3zIcqP5eivHMlIFxnTsQvPIYDRT73YjYi7cZI3r17xGp/lJ9hiZTzF9l1evw
Z119/Y6XzlQqEdXrTFplTIsSfbKFrnrmaWXmmZIp9ELF+N4elXvZ7SzRWfIhEO/18GSLIRRaPiaZ
K1j71BtBsV8iwX2oF53nenNtLS1Dh8Ro3mJjxUzl0qsaq2OXlNx2juWEqkQot++ljzL0LMRR7Isi
XK5IkISPCNMSuLNvqBErNnqkerTJGd+03GOzYWXKFJFvLZaUVioiBphjU+IQj/1bRaOXN6IUQIoF
kim/NeVeWEwEBXuKkljq1sMjx81TSav2kgm5aX5sqVF0UnGrgrFbR6K3uRAf1MLZEP+cDnk29svx
b4kykvPySFNTr1It/NDMDPhie1xAbMwJSTIQrP+N6dchrqU1sZrsz/gf8/Gjv3CZ+RnxyfUyX/AE
0eWtCAgbWHRbqQReC5GfVvmr8OtQRHU0GrY/B+t/KGE4DppptO3wYksMJqPNh2UsuhlhWpyGj37a
Os6UdQeq/U2+W8ObJ0M+tGf0pQTmPRU0SpPfF4gfajENidV1743uLXicOXjJtGB4PLmWIPr4R1Yr
vW/zzwx0w7aZ4bHwLz5HUaNlwcBafL+Q0Kbiwdgh+B5bK2BDK7TsGs65HISV6c7IEOpKwcTxW1Mo
1SzqTK0Zyo1Sb7WTrGH1oYJ/fkHvQvGK7j8y0Ad3ZaWgudFkh73eEAAb720ncGkd61V/QxEZbPX6
3yVPU88tmCnNCI/H/VsGpE0ZKoUopSkia/iqGwSkUmzzFsygXfHvgXUkB/qtbAAIac0smoybtxlo
2Tbo8yTTNpGuROrheyd5g0lpzUp/BCikp89f6IqBMgoZNSIvU/+I3u4eGae/Ce5gzqecTFrnWBn9
Xj+zq75/fGm1Jn8WGJWevShGz8KSJNH8AlFomWlIQzg0+ewahycAQJAIKtlOCDR8dTeCV0s8t/3B
xueIQTEN5GELsm8lg2QzJWrLxtyDkQEPKeIWuGSdrB01prG+FY8nz9KiGkyyBPFrV9xjhjEgNOyz
TjTqbIGkXxwlOD8a7DNT9veiKpEXBz1GdMii66jZyNImyxETtFlcLSJjxZIn8pzSNDBFOExare9u
KxTBCQqmATVKDvhEu64Tm4EALKRavq6IJgdl/Zan+FQCiJKxwhK3vN3rHfFP4Dlrv+3vQ/aeIUQy
1mweUWEBI9/S1WbswMfZ2Yva45n8SPtO+EXZ//0PuLLZPzcZ1HsePLU9SAQUfmIMmGPj65I/W2P5
dKQXgHqJqbni+YIsM36d2GroAPkjElIBvu3sLRCGHSCgPgNVBWsSKXOheAV3J23K8GXHzfM/v/W7
3fLpDCxbdgnBrZjAoQKipFF+Sdc0KqE/TZVKId4HAYo9HX1WGufP+dNzp5R9ppFcyScGLIAeXE85
yd46GV7+wBUU6JL9Mh4ZM9Npi4KI41pdNAf98Qj8TSzUivFidVG43xwaHiBOeX0WBtsWGf4/b5v6
3cjz3bTI31GusWbugrEuLRe6u8DyZpNnG5h5KZdykjb0jqUqV4WjgrWpIj3fNWiypOTcG2TTk3KM
goixoJ7pgXFWjRjb+jFZvAIIcwgsYehDIMFsh4kp3BjevS4tn7y6DiCDN0x2szEuaU0Lds7dm6mh
GZE0C7Cg7lohkx4djyBdnNaSxwk/cOe6uCbvj7Xf0mJ1yIOyU+05GgwLN3xsZl0rN+6aBQ1UxiAy
t67qfCbOGZpafYAJHcU2vxox57Sk7+ZG28//4eriRp89pTdwgOqg16+7udfzrqzz1mUFGkKSR4+l
HhbXOnIi8bCyxhNSm01Kz/RWqIXmo2BXHktB/vrh0ZwgfRDxifzPAYzcsT8u7uFGZg00Od91zCdB
5zQt5Jx2ov93UIOiEnluMPhPuduqc84heVUXSXdspp6WMXUTrdvsBxBb63N80dfconH5UjbIjQAD
ky27DyCRBMUWPQqVdiPG2uKO23MscbCz/vqHGZ/Au7aVcCgJHAQSnIhBRqPOw9LrG9Z0VNl94JUp
DvDB++ZF5k/fNA+pCTnG0es9FtAprBnMQtGLhoFgSu5kAuQ8MD7Mrqn3KKYrBrXKgxk4NtA5aloG
/1I2dhk+WCyB8UxWGLbIG/k+LHYHejs9pb0aC+HZG22z+rjlwLWamDETR+F1vQ2gDpYBfITr2COX
mFwhvK+9ik6RngcxuarwfeYLe4v3/UWEe5KKrTSJc+5a7jcMVH+O3olZLYGb/o1HA8ghg3Jy1v6T
7ZUG82FicEUdm9Fm/Y/xAPzKJJyMgjMeyFhC9ZHgV/lYkuN31Hg1WN8rWETGb3WwC4/cVu1icGiH
8RfMssBvrOP0UrDDZGHxia+cVXF9i2WB3NdaZTQwqIANDtPGTEZxgpZt5/cPV+YV1QquU/FKHvyI
1aJ1dc0lVmq6tdpCUP8S/dezx4bR7sEQSAlEvoZWfwbXtujWaZSnx9AfC4DuYfDje17mhyrrUhT4
b4/NVqs8+dnKg4Je49JPADxMCKP8bybIBgxmXU3kl0SuFKng1RQZmUFb0smw+UGZx6l0JXdfmDuf
pPJUnd9UIfdM/zn+0Q0ao5MKceChbCqMsqEaX92KKh+bzGI1qLyYrKFw7aCyy7/12om8Y4vXtBLF
nvbbNiI/3IsrT0KDOxKyxRfR8ernnuKD08jqqZUKZ7c52Xb2TCY6wEQtNkBTpih3TZ8eBnFZhy6E
X5rV8CigeNa0OkPQEwyAWMw1WXk1SEzEgFbHJyJegOUNoY3dZRJoZoqHIe/DGG2sfzSf26g+lXrD
pOwURnTpQiAX6vjT/X47Hy8ofdrLxgvR0WiLVthpsOnNMfQ9cuxhNT3ncKeWvnxC+2xm1b8DAeh+
HbH9E60yZ8L3Fbo0aNPqWvtNC4hNZFOYH36pkztdy/Zl3uFvguEzJYfjbUykIx6yQYmmLUH0VUFP
Y2DPFXSyaD3gNK05YvjImaLpKvoagVF9MZRRtWUrYY/z18zW5ngOKvX0rWhuTLd0M8IFCLo0zI3t
28SbFmDHRsbljYW65kScaI7biqF4hktA34xHHu2VTqOuHIHQ/bfIsqAb3AGYjqrvhO8tcjcgCX4u
DAowZCEIP02GKi9k/3fnRByp4BdGWrhDiQ41f5ivK/NuTRxir6WJaJ65H9iJrEU+GyJ04plhV5fQ
VIGD4gA6rQEn/KF6h29Ra+ccIVxmqzGuKhodkb03ImuZOl1KSQQkUJpNbt+RWjW0oRh86c9Vorpx
VDvA0kTVILwRyk95G5K7L24Iy8ExsILo0uTuDbpsoO63yN+mNlndh3449UL14Ybvcpad1WeKlOGd
mtOYOO1rjDc8Q5oY9jQ3bYYE7RCaxkW4WO3u725mwTnw4wIjMeuyD41ixCJC/qm+7d+niIza0IlG
m8SHNHS8dYKhtA+YQxiqQb8mRE6xkx5AyHxFxpYvbe0DPzwUv2uiCl73TU50F0sFYEHrV2OVNrfc
nV80s5xzSuzka5/sR23efpR3eblaQRVzNcBPZBUsheZ/KknqC6nJAbWzsbUTOibAJzLVVpjeBpZA
RSGEdKCjovCNxdEoxOsNYaj9GctQyHnpdSMrDm8XA7gyqzyRPkS/mxdSxf+ZOztssmk+Py3hZakL
dPrR5f6O6Rs3y+u645Q13b3ukw/A6ri7hidmYejJVZsp3CgVIS+HpeCL1R4S+815sYkFgpuiq/9t
zS+JSVkBl+Hpb80BTMmqPDqWqnF4Bq9Hwl6e/mqaXqI6+v9YRtYRx92050BsdbgsKmSRmYli+Lh0
7tDHoSHL5CIfLOo3JI2wup0AquqfgPu2CNrwBnHfZIHCSv3gDARmiP6Z/08EdI9SHtZg7Ij4f7Eu
CM07jeFa1JR0oUlnaAMCHqtS9wzuj7nEGACvd8ZYgfWeYDvVUQMtkq7vbrBQbLe35bhej40cQssf
XCn5Mb1RmCWDQldI+mRSCmqRXV9ITwyqN2w4SSR/yYoYdzMtVg/1Lo7pud5A/FRUMxVz6HIfjzHh
Y5eq/t9so8xA/9iiDu2aU9U6bHAy4oKD9VJ92zih/6m5tWL7Xsits7e1amwlQKJSkhpKetyFJIJX
bpHo9V0ZhM/w1wEp28xIYzFyFKv+munk5C1PCtPmqiUlGFafqQ8Tck5ue038UlbseCLY+ob2plio
6l+yGfCAmnVQjYva0Oa2pfeVwzXTdaorauwdbtJko1uabel2WNlenGUyW5k2bmY+v4zLayw9gbjz
QbqLVOppZ8JQmJQI0Ih9Mj7o03tDDC1RiMwt1ApKSbHQRtzZ7mue+9oGjWk9NSTG6bUayX1GVh34
pogjaSlNGE71nKMl/Vb2cK7VK/YoFFZKZchJX2aPU+L4cWUxVM2nrMPdVxEjQEvimwNzwxTRmHJd
S1fEkBwP5eyN9pkpO5iweBKvBos9LjPChblmluAbXh0cwwZWsUa/TRJppfL3sR70nD0PlyzDgqqi
c/ypmE64r/bBk3BAPX08/jgBQYtXSRZ1Rqyb1PeYYaRl0ayDc7bAQJgp/6m2jlH3cnxvZ/ndJH6E
m5/zZ7oeXySuJVBpsYumba456vYifSDdThQRllckbflfqzOpX2UQiP63f+sD7zswTrkECll1EcuM
+rcyYJ8r/gzDRR/8j37riLrIg5ozxvu+eUJJlMg8xZmn/7kZuj6v1YB5FpnHAEiOMQVcccsliBo8
p6CCFIlfH71bPAlX3UNeYq7gcm4UnPgNERz8/jnPeZRn6+Lc6PSrZwqDicPCBA/xiBm5UhSIEx0X
sbUv5xtJZ3Bg6mhQHTJ3daGlpZl+MR+ZrjUMY2wNXaPZNdoyH2lr4UGOdiGaqAq97llnFMJMaMRp
ycJ9oyjx+hrYQUj2R/eLPn8TTJxPTGORFrj4+8/LMjw2WSGwFklf+sO9RF2QswEed2omJUUa27hv
tVxV4930Cp0z9zzYYdBwucOGz3jT/zcqLl18Qq78b/Pcz2E4oNGdUsX3vEKVM4oEWjbrhWO+gMsj
v03mxcXABNPd3EPzpmiCiaLcRXl7W1h7bO05VWFsItIVkx33Qr3nePphLXBZGzbnPQnkv7Pu0Wrb
/RW7bZ2UfY5JcpmTbwlOpzNoJhDI3idi3bNcp8jyxCHez+VXd2iw0fzJyaAQsW46gVNMSZDZiHmm
cxmJiH7ZSVGGw39E2TNXCPLmFpl21P2WSqwjs47Z9dBYXMUP3nGEERnC+I5WQrqwz/44PtHKrE/l
37QM01EwOrt8h90L4w7Vx/8ZoFJW812Q0hW3/rEXCjcvKXQfTEKQ0Tie8LGZre75cyeqSjPlPcsf
ur3KQKInSj8Tc/litVv+2qP2J5sirRUkq2HxxmHlVZHGD1eFHjxx9Z+0juiFmZDJwq7ou+6Rspv9
7D1OvxuR9itnKZgTONIIRBARLD/1PoKaQUkUJZszOmtlRalMa2FKhOTl6xkmLi1de1d/nowpR/Vm
LCJL3q7cCFoz7R8yphavWVvtFa6oJJiOuSSo3mJBk8KIaVE8LdVgZRhQ3VevekS7tXpG08KLWDYI
Gaglnsff8O0ddRSbYIjxD5n7QuqDFgbNA5bJ3O3Sbq7mj78CL451GbqLJGiAkfkoAbZvpLiVsokJ
rwlwNiPh2ggh/iXzxjgSP+hINQd3RQDpSA2+sV3GStCIvhTEY5EQVsl/KkYS7hN4l/wh9iz92dYI
lW9xYUZj/371h7WV/6zCFLju+IV3DqbWivaRDN/hUNu/g6AwiuagRThE3ASM32KMyRrtIpiiz2E/
gJGeD41VJN5OuSjuRks7u/jRNBtg6/tUkXlUaW0gcVqtgSPpXdpepNWIWV/F2eABQ7wc1Hi4+++Z
XXjclAgPWdTxHN0w9LvH9gCHjnOV2e/UAUk1XNoHQlPEc9WRJPiKCWeaxfTuXi/gkb1YnA8sihWo
RuCbBk2j6l6tkJh/Mu+KbUe05bYCoZsAqj/1bS4eRc62vz5aeGcMzwhKzUcqklvwyTtqNoFguRfc
bUYsR7K3s7EJiTbay7YmiZ9uPAWj6i0Z8gtVGACF6xwaoNNpXszlYGYyzRgqTbudFvfNvkgWf9Lq
Jxcr5gg8v4CCGPY1XhjfunLOl48PQPjDV+aWwfPyG7s/yet0KCD76lmaSs2KYb9ugPfx250DOqOy
fjEpDgCYfrDvVMUC4MulUM16cs8z3elYllmur1fQGX3mqDP8SpzpIgMX8epiWB7PL7m11QOqTCGb
9bsQYcfQrEYsz8hislZI72jQ01p8GIJD3jxIbwVKNQ176kHFUyhy4xRp9FhR6O+VD9fXyEEzMtzM
mJWiUZP8dCrNm+jr6BbwoxpFbBbvyY9cp6jwbUy19mhdWp2/c4pwS/7TO2AsB5mRYIrUW8IT6842
UzPO28Oi5LUNi6XHpDbtD5Z7paSJjgxZ2PGBHn/Y/vpZS1UpX3fNtM3U3gxIsqzpTW9gTPgAI8Xe
vJ+IIqMLQ4UuN1B8W7OzxxslOpTHwvxT6nNys9T1LqHRJhNDLrxtwnT/TmHkczS59CeFknId9Wh2
lVUVfCqPnFkkqCGjD4ujKyhAa/RxMoja6mDKNr87/bthxyGufdNB3PiE0bEjQgnwMktjs4+qfqdQ
5eH2HQ84Zc7LC8hxV/wjRDIK7qgPFS64eZ1NWPLjQP6CbwhprQtFj8YKFgYzfhJBKWZZdRv3ZHIc
5PtjyEzbGqYc37VhG73BNbmU99mf9x0aUuhFvgSZGffP/jjPUqt1pVEy5oa+4Wotg/CNcjKA2MWE
2qWiRt3cEhKRUZxiSBjLyt5EMO462cWzQP3b7TZPJCGW/2XtwODhSkOeX0tLdf8ZpvIujRhyeUUZ
IPEwov4YDk2sJSpVQSd1GoX5bqSHwKGavXDJs76TZ6tzouRdn2vOTPT18vQC3jOTaYWaYF4aYtF3
SFd2wADNtn7CYubfcfAHbYoqThCsRMh/ubq4MKuGOcaRbKumowSjaqGVMpeh0lCQm20N1ap9tr1A
INNjZQIbk+OOId78Np3yZSZEtAOmtwH0pzfc2OgNVVwyGoSNOqVQqZfIPmKYWYpxoCOP0HfHYPux
YFLbFzyElMA7FuShyk7Fcgn2fej/2/8Flw6RMYXzy/3G+rmkYac7JaOr9ydLAL0si3WDu8LEAiHx
Ba+r1iJrVUkkEz0lN1C2XRTalHp10E+t9XNJloUtB/2rwmvhOr4FkSv4TB5A2IZgrOwJPjAhZPC6
fgMYlyxEYrqWY4xNzOYxnOu5b9iZxoisl8fvaC/19b6sXd83w3vAm7Ik+glBy0SdzQHlcdqtxPvc
oZGU17z9OE69/Y6Knk2J2EiaRLBHFpPYTDDlqiPNsFYTwlz5Svn1Wa3ptHZl7ZN2Byzea9rpErQx
qy+SlDSKVRc0fkY5iUe+qxdGtjskniRRZ1M0eyaSx8Gw8fwnjhSMGjP6BvvuUe+GHGrZbeHvJkM8
D8cB+Ls7DM50nsIha/ZJMbbvcGNdUjeZzfntcadWZgOjXJoKOmbGlAaTfQaEpdUz+Nf4JRXS5WaQ
oWx2cD/4glMDiZKwf+uQz3ze6/ddl3u7KQchWXQ+06k98W0hWaZvKPuah+abutB3Jp0Sq+O0REnM
PPCPvIC/+kKDkpFS14Aqd9O9IeE33CrgTyY4hy+om0zFkl74Hm+jUQbl91GxEl6AwU8I7nDGaGGP
OcGVzDoZJqEYczeLt4k2y0OUco56NLe2yxmuEBJIBN8UewIHja9Vo77cMiVcACZGs2w6b01DVdo7
Zacovb/Gyiws42JDdnCSmigSoygR8Njms3rPLbd+TOkD2/teSCPtvMaEd0Y9GfvpP0H6b/c5mI7W
pjfOkXdEOO2fLs2IEKzQY7XcKMbVIgSSVNg4k/XEwkAooOczdFt1R6eVVYGY57lNpQzQY5EfMdSO
IQ+yiGkU9QsJFnPyWgwZA5tjQ7ipD4ICmYu6x5s+R+KNg5Ap1EG5ZBfxQdt+HrzDl1zzhanr+6cP
7TAaUzoIWmnJMP+SgAlw0ZFGKEvqxdds8tHSOpBsQceSPPhzi289FOs1SOo4CueQisIE70eaH0t6
xKY35DhVU5wafeIB/CUSQwxcbT4upwHOiqqPOYwqUQ2SMFj6TK0w6v5VOiFsGMV0zmFKXl421yjH
3Q02sqk8Btq9LRSGsnmLf2Qqcvi+xyJ1LFkWdDgRAu5m3chZdhxkrn0jECqvMv07j1l10lHMhscj
AnE7CvhtBAFehS1R9be5B0MMCU8VXiN9U32h9fXhSV0w69+SUMoU8s3Wmt8OP/h4GmKAYs0xlgkC
ia1KkU+FOeKOh+Lki3hdihB0FsQCxH7pUHIhK+aYReNHYTcQtekPK62VuAgHYSLgPEKJRe1q4ifI
sqn4yWcnQ7jsTIvGb5UTKBPnyOFr5Gzfuyi753o21q3PBfgax0R/ZkCoUmRbIIl381sgLHosCXct
xpAWz+Fz8UH+/2EC7hdssPL5OkD2LCAgnrfEqu+C/zDfp3YBTZNjM5G+7/CrVLRH3V5lqAEvIwLL
Y7JqTKI6RjJpFFpBdCsctx+VkJBmW/MtCCNNLXFj1T5Vd74KU9rZA0Usoq7Z1eoYEYx80DkkIdRD
zd5B8L5Xlbtew2iSXd2g8QLcKnAOKhn6Qod6JiLws0QJ0Gs8cI8fIsqaKWyyGKt1baSwSqOfyoAh
Mj9tMVeBn84fi6BGFoLE6FLDtNdMSWQBB6+QNK9jS7WFHxbxvb2xguXTY1rjkKiGBTUjmmi0uOsX
6AgeVnkSavfmJEIhhxRG8kuvqTz+G4zDvxvhPGckGsBftRY7IHCCBJycnrxRF3GjS8x8xXtymntt
ar1Ajwe1BdJwz+vuUsNy6ScEZuc2ZLYgc2qpPhL7UmImCYfxZRVuRtKg9S0nWgPYCYJj+3NclEpo
VANAy0KeTlP/64xTeQ6ASr7xo+Wiqo6xtWKIGMTFTDNCRI+OKl6P6yCgJAT4KVedyRbnYFGPZqTl
h0HgdnzzF077GiSbcW/VpJ1nFe/3oN4kso9KSvt7VHIctwYVqJWqn5ES71oC3+2UYKevfpE6L10X
Aj7M/3iN7eUkVUtIdwngByi19Ir7IFxIUK9hLupPBaUSMeEWKCkzHncUK0uXAfrJv0DO6P9g4A6p
7H0n6gsRZ5tDB470s6E1QfsQqPkngPxSJJEF2mzYpUnBlfcj4ujFG7fSIsz6Qoh0y6h8UZvsDl3f
2pJ9ShN7vwEZwTSfyG0Fm+QWDm+tYXliyASVh6cmaWVMs9v7JaJ9OBqzVAnZQdV309ZlYavEcJE3
GxWx5Yv7fRAnXBmI/oX1MjUv5eEs/XRm3tmS0av+2CGNw6S8fHWtVsJxeUY1ROhxLQYGWLZLW9A0
u3Xd827EAfLHDH/F0/Kt/BH6VsCp3tuKEoBnCn8dx+2he0H+utK2MU7rO8IUGxCNPw+MQt1hu+pr
uEIl3OsS7POQD+BTFZoMjJXOjmZJOFZfGF7k/b5pbtOZ/cTvniENOtyDm5N2B6NQQnVicADlL8ZW
dYHvmIpseQOkb8G9NKmVauLEWimwl/S3lMVJE+PTQfo45lveIOWkLo1alSc/j4wjqY1p3gw8HC6I
qZeA6aSLe50H5bO4kKdEzPXI0XHG9cewIxCR8Ew1T3uZRrLDISWXwTP8JdF58gjRKoX08zbYAsCU
GKM3uUM/VZ1C0KUEmyyseNgXJfVGgynFHzkcFoUe/TaXBsIfHJW00B/bS2qFPCnT5MUk3tBS7JWY
S3z0Xp2SRc9nF7bD/1iDyj7NCt0iUd/W6Q3RBNWEybuAFq2MYryO6OxUF9rEoqh1Yhix4fSbh6cL
/f6I6Y5ThecWVxUsjblFNlnRWTl552BUPbxX2GsACViEzuqJo7iaMt83rToiYtVDYWWZ6MbQ8wi7
F4DXuNifaG4vDMl+cv7Z7pZxPmlNQSnwznfDjTC7WGcZEd+C4vv2PBFhUlpNy9L2jPwYrsADgSug
2lrjvUS2QRRf5hRCZtVxT77Flun6au7GQGWmxnI5ULa06+yjyJseEzsbuNZxprj/PZnWgLAtr4Wt
8mdAA2szBE1HhkaLX93uNRxHOlF3ul6s8XtfNO7klhxhcMVNUi9EG/iD1YV2DyKrOlyZwIZgtnqN
zERPjWcv4XEt5XfgIt1T+bd8TzPZfZfOIgB3DJzyZQ0GFwBxt1g6S7zB870osckOh8tf4nX0O0zm
pbAQxWqXDXbZJtAOdNmGsxcdSSXefn47KXeM4lD8sr3QIyGzc2pWEPp+eSbBv2D+BC33oY4erJO2
dDEEL/7J4PRh3nayvl3yrA2esOMHgs9+rCX84WYhCzc039mqX+Wu5teVhWHwfFIk904QmUe3Sm1+
iyntgoo3psf1/deiWyz821n2ccVOTOTk4RCbuXoCJgg63hnAcDQ5UVg/uD483Oxp3PHoRBFJnR+9
foHVIiNu9733WB5OdTMO3/FgxKM2QqkndOz4l3nIbAjrHm69d7G/38Kjk/FwmdQ82adN/HoiKmfi
kFs4u5vP7e3M4LZDAdiqzNxUOpDPmJmmvnkET6uK4tN8eh7qu6vuq4fr1wpxkJ8MghQixA1m4aIP
tphilSRNg/1Dqmwkw8lw6O+58MfTbePJcT6dROO3/X0iphy9iI5OlvyRFki/O/+omNqH8pIMebRi
gIcDjIvFhRzAoADWfvYkhSKlTr0iFR+5FmOOvRuvaF/v+I6jOtFXa4Bfbm5CxqykcjXvaEtegVjx
kt7BRA1dvbrCw+bgETpQTZOPYqJLa3jrYsyKCQe4JI0hVohlKdvjKAYQqSpZysGbKKRWa5mPQ6/O
u1xNcmQ6SXE7CuRUH4b3xT0k8vM4riYo4exH8J9fDbwWJgT2D71RMfqDOhNXmZQSz9TDyv3fxmRQ
INgKhLdv5/zeiA7byOMVM27Z9N/kAEAZ+T68XzPqasPh6d5RZ5IBxy7qCHZ2ecNHrtinJ2MSDCar
UNHa+ncOZ688t0WgZKlrrCKvFoS2awqk1RnYEul00tS8cx/LqT5qNfLiURj9Grg1psdFzv3c1kW1
2Y4CpvVHD1BRHWag9mYdgtFvSlaAYHg4vRQkHyEpKtjSlxGZ1R2joGdytJJQ8DZiE9QWeW86nOqo
MWm0HG+0Boy5AIrOoLu4ylfj9pTfzMR3ywOtYhe2+7fcFfAbw3MjZmmNE4UI4TJ0NrOhPIhOzSkN
JfqHqXKq+zfinFM0ZXM8USww8aqcXklxQ4awywm/NvIfJxFy2w8IjqlqGCSU3eF5+ZtZdcEPlyyN
XlArv4tQ2ot6QZpZvGRGYrn/s7CPpPB9KLleXGHkMU2cmmCwOlNdnNs4ITA2+lDAa2pckAUnAfI3
5bjITcTmPH4AGd5wjIiypefepByaCKBsE1YJcCmLn5q7nZlZRJFpG2QDY4cpQ9zTun3JGZEW4LgP
AS5pMx8v9DPa7jOJItMwQRhlEPtGarZFH4UetCTVhqzoOSvWN65MsQuKd3VyShA/u9NcZn4yGKcV
9Lyi1BOcXqVl2BAx/dvSoqcGiPLxkdduQmF6lmfe1qQkY2xKbigjG8jWV2Nb7xM2YL7uWPYe6Pn+
4lLqIfhXYQhuRIwv31TCsWX40ukhSoCjJz46StK8n+3B888nWWylV66aXPo7wU/UzBYuf7v9gRa+
bpqsP4tK3xpprbrxctawryAp2s2tl7OWJ4W2RH9J7nxFQk/gqI5LAaoK+gZYeoBfIMN/ElgvlPcv
/x4dfJMudC+fqwMdsg960/H11dXKBqFre1O7Gdk+N7YjIWtlmDZO/OtbJ/j5XKY49FuOfDEL1Bxx
9RMdAwihyAqD5onQw+OTe0HB0k3R0LG+M91Dxyd3CpunKBGrKLNlW4rQ5ZOHrAQqE5q8ckXrZPDK
C9tn0mkFHK6rfPtshepRVNPrqOo1AFOygQ6e38lnMPDFfnnCOcvJ6z4G278ku3Qr9ehRXohTDQXs
VaPNRdWADw8qVF54n871emxgE5lz926La43cZNAd7QQoqbB3rzB89IcjP8miBBoXC3bFhCxSfiaH
tUGdDco9TchcU/QXXpSwUfKVyJUs9gSJi9VqMln40CistT0sOTPdpbfdstDsEMcw0ptMihSgoHn7
55XBzztAl1yZsTaCSU20JICfyx0bJtltuFEnt95HBHAwm1HGXOesd7nXES1nLqjTuIyJp5Sy2Qzp
1OsWHqzAsrIhb3EHvbgCZW6XpDE9RdNa8JY8GjeqdDyxK/qkQLqRfA5kI6N7a3kP78eU24KVj43f
JWbYtwdVo5vFDATKU52a0tWqYloF4Uan8xSyLhnGMkWvE/hEmUjgyPNRw3iqgbRYoLnST0RHGK/P
eM9//xNtpl0m8bRktgBmTep6o2IhooqjXHWlePSdgI5P45Wuy8zuZgbFL6DV7eQcQaeuM1YB4Mit
+prjllmNcEu1+/PNTP0Oe6QwiCBxiy+JPMSeQU8f519/fSBR6pulGLvnvzHgcQTwKBrruk90gDhz
gxJEFDsOui0dJyQQN5TseuUstJR7zf9kaY8qQjpqEfKr3LAKxv/W/GG5UG2h0ncVTXI+p1YvihnG
vPhxxpxdXBqvMkAyu4s1COwj01OVYZbdyVr4rSvnjgOF/sQHn/komyI/A81o12ODbhfSiJGFJ8Zk
AUn48xbYz1MuKYRBZYMgolCitqiDesCYLpRRswXJnvEcu5Sreyjth8jvTa8xBfp7YnrZ7TSw0U4+
8VaDDTlzcJNq1zBomf4Hn52JJXexcblFzqU/Fet4C7ddVLaMUgSs2goTufu3kYEdz5suu486MeMr
qimm66cBcWSntSCWf2cCFAOS1Bfx3S9KVIQ+wPT1RjQRc7db5iaEnkJkZSI2FL5vkfbHQHFFnuVm
5NjnBskqdlim+lbxfcQWt91BcoTFzaUt9vD/1UoNu8hHhK2ulgM5k4F7sAmtubt8ZB2yNHqb1nGz
tfaOO6SXnoBqL3MWRNuyVaPMbVWD9xfp8xgDvf+vq6FSY4jU4Qi5CnLZn/9ZBXUvxFUdh7GSrAzP
eapV+N12DuqtvV1u6nATsNcj4BcQ4A8itNxivAMVklVC/oI3+6TpFHu6k9Blqx+Jb7PLeW5jbNj8
Ruf1iVOhGsS9qJrpB/Tnu7/xy9jG9qQKQF+g2XVIn1h4JVGpQsF4pIvOIuJH/lYIIGUH+g6Pxfd/
9mZUymbLnxoAd3mZ94Glb3H9g7dufxkalPVJ4tUcq9n8dLvIHXz/2smsnqDFitnb1LlD6nFdxQsj
R9Xc2qOCv5rNyUlsHwes7+c0NCxywKjF9l6JXV0GNeFL9Zeq1F6hIb/clIU+s5EyuQmOvfM77L9x
Zx/il4QKpvWZaUNXKP9jUp3K0vdE7qkc3Z12S+ey9jVY0lWokHcxjKT4VX+qckN8HmgR8ceAvDWl
hC8rq+7MPGBWDPH8S1dnvK3WQGyck7R8XhgQGaysRXqnVFzJrGJAzLeOhBO4eMPAZbXhrg5XKIdY
SKCJYwgFWaMt6Pz+IBjDSMy+twSsMrxcWjaIXDgphqVqTq7pBcUvL51DzFbvlKhUtjsf7vRfX5KU
uhRWqlmtEzLnBRHJItHKV2f8qUVg0KJnArPQ1A6Lw53pQ58jmw79WJnoxX2BGulBE5jLfYgWHcwU
aaHRSqUECaoBF+AVtdIYPDASIp3nfhvvFXMfUmHe+KDAFyb0MBVgI7StL851mGikeSvjhm7Mooqn
sX74Xg2SFYzU8/51D41mVALrPsCdnsvAwyE7USnUOYaMljepdP0PWFbWOdMKqd9kHV3H2dbE7yG6
Z889x17RewiqAnD3t5yvJ+dvn9TnAJwnnR2ekJ09kxWdKFnoLcx1zJygk/kPxX8qo1v4YjHlJ+hI
/jPedy9v5TAVa5IYjoWDtRsgqfuz1kHeHaN1NtrYIq5C9SleseojwE4CfVb2VpPzC7uC6mwfksJw
77vwv8i9F74CSVyFIXMxXCqiLUDm35oBDTVtaO1HO9gzXn3LP8UKVo+e7n9pKcPqWLlIlJnS2trM
PxT1Y/hfBRjoBDbytV1gG/h/c+PuD2yJZnGnbi58vmAwDI922fpHGCrlMUn5l3X5PWlZKHA9TrmT
n/9KaVlEVyZb1P47c+jwzaOWgyOYINWY+/3z2B2Z91LIu54PQZZxujOI8PbCkMtDyxEHivKpF23H
1wvgQl8FD4cmACqItVjwLS2WY8WKZNepkPbILUhn7kSAGGUM+tjWHmx8PTqhfpVYN1pjE5cRASoG
TvG134qEROh5PjN3l0jABm7uMOlNtqtJAOFCLeuPW8WECDCPIlrkWOXXkJkbIEo77Ap+6YHNM5Mk
aqs1ZcCd0hEmgCl1jPEb1WQJ7AdHLb22VN9M2RrJkAnbiMePsuHc2ClqIJCWCqti5vHpIC95AaQC
Hi7SPpSRN4rvQlf0nrcAbzOUdAOA/StjMU+62weghW2QGNvqUhx/itJiepjRWzZpeqy/gcdv56fC
1KSIRhi52+13sSNiaZzdgUezS5HJu5z9RgRwLy3FOaoouHgq9BoOjyhN6RvezR/nn9Apdukkvvl9
JBVmFXYxohUiRGIQ8z12vm4C50DKw/ppcQ7Z23IPOmvzmv4pXh7nzgiXdStqsuynrx7gW+bomAI2
6NYHcNX95nYpAQTyU/38H23GNt7k0IS1puT38Vsz5jtLkN712cIqpPX6Ofi4rpmvuITSPSSoKPO5
5XF/t0Fg5n5LbNdqzUOcGjy+giCr+yrunR8bMKu4XezcNAUfHj2nxK3hKDKethHYmPP68IMPsJnd
aiGUIYFfVeuoH1aAO0sM1rdXdFG/f21nYKdWtbiYDenpQpwJIOu6XP1pke5n1cNJpyrgUkpLRiLH
xcPwnKafd/pfBX+Xe7pJJk1YQDgdRES7ICHwkrmHMJ+Q5Ts+anesgcblnZy4NmARgz7TjcR3srq1
K5MLE+IeDVoRGRNMof6/9WU1drT6H+i+6i1BPMfdlulghxjoDHA+5dZ+icFUbwya0W9rHq3hFrRE
sI7CIuDZJi/SnzchaXhi5Rqhgqa0Gw7CLCNG4NZChqo4aFHa//3phEFP8IOLnbQl2O+Ymqrsx+22
dGcRhuMqIHlRAk04QYcypLk0kXW+QhhAgfB7NBam2lXRq8Kg0ha3LxKRamw00T6vObmfjP12jILd
kVf7lf2ub7tt/eed0qtxNTeuXrIMg6Twjih8Xau/BSfqCQ10t5uKVAzuWoKOjjAgDc7nVleaTAXb
/gfX4Z9QrvSiDfbPjH4k3NYws09w3i13NIWBXS8xmb/+vQgEaX4Y9Ii7JCplZ+ppJ+lbbuVW4K2+
gBmEWxO7ZHM/H7fscCceXDtMdY5SNnkTyGqb5sl9NEmv1LCY3ozINf0PpZnQYTOVWOd5RAJDi+Zc
G/xAvWPtCgTNkYU/eZyFWcKdH8VsK8HFXReV091jnliIwjcw3z7vqdheddiPNPFBnJ2Q9n5F4nTD
ij3GCaaGWYzJskrOjwEi75Q+eubPYrQXlxfKyXwsG/fQjaAeJo1iGJyhI7sYpW1SL94mzaKLD4X6
d1UCygztTKk5ZvSWMvrftT2/eSrU6ApTRzYt1NmDb35BjAPC4+gZ0Mn5QJBAUWiDJDpwcoYS6MAT
whuho3+wy/GoTGyY5iIzeqGARMKeaL76bDFII22uLlzqeNjR/SN7uwNJQPpeTf0NSQ9UvbTwOU1n
Y2Ihtxs8DiC8KX4KhRyvk2+KYd2CSWsjBIGahCeU0Wi3bYfHQmPBSHrYJ3ivk4W2svqrNoLYFq4L
snAEO+LM1N9/H1/UsG6E+gzokpmroPNWNZa40eCk1m15Z65POso9Q4Dv1l41ePjA9C5ClFe2ws+B
Ps8JugtUgq/L2/uC19Cd0pqeRlIW0mAEK1zUb6N0lQl4wTfnetQRk6U0hrBpRe7+xQQFq6BxcpL6
YiTbYvgB5x2/pHONJM+dFbajQDSF8mSSlUbsXcQz7KFCcNZ1cMG6wcrJqv7xHYp6W+DE6nECcUbg
F+sPPgj28eCllODrUPFMYgA1ZjofIv1d0cvBz2AxI0ar+hN41lK+1U3n4s5KmB046QdeG/mwxXtQ
GOQRwmUJ5wMjb31qG0pj0Pjqn/GirHmNi1xVpBDG9Caed3Czup01FyeEeylL7v8uSD2+KcIYMqOW
5UV8UXJvMbodnBR4eMpHMA5Poczn0grs4BoRFX0MElhKnRqjPcjY4c54R/JzS/96J40gbA4ZrAkq
EqUl2lg1n6vAgji784mOPpv4vkXdn7zi4xSi1mlEklcQcu0NGYJ/esmQOFGv+5vaOZtNolNCfMob
E05BIqSIJLPZ2loyXl6haF2ieU/kgCe18CozVShyRgpd6t6WHDESS2EAh/tQZVb0YIm0UwC0Kmwx
UEG3v3SZUNtVYfvs/sPkrH10TfmHb0O+JQOyM8mElq/t64LE3Zqbz/IWjUUDEmjzXzXcaxC8ktr6
NIEZB9s+p7UG9dQMh7Fp+e07VkqZNY2pCxgnf3th6NwlemkXCaw8IQGEa0DONirABR4uq9bSW2ti
xaaa2fzroPFgUKFj0gWcewTdU1dTuirIgKCocT1EJXiUZcIlX9jE0DGjfYcFVL50UiwW27srtyiL
z0hs+A2ZYG4FoqW0CbmaJwx2BYDpQl/yB9sEM8r9dV1lzztigIg48OMiuKn6SXrP40IXYjhNfmEm
WN70a2JfTuUUwjiMgSTJmbox91gDnUcUuAJUBbSgOpxvXrA9dnvWKAwx/tL4jQzMB57CI03Lih8n
zQvqP6qsGhLXGwKBo5J2v3l31fQQJSf6xhMabJB15LperH8TcAz4VB5kWSXxUx8Af15EG61PRySW
Hv1XZQ1nYVxnge2eAdKLX0sZw8wR1+gk+AICJDCCRvsC3S1rA1D48CjireHQq2U6KZnWR1xFQdmg
MQXJfoMoz/UOsZfZVrwAV0onKEuALV6LXYbkCf8glaL8LT9JSCp/vQGcMB2ruIxamnoIZpSDfdiD
ibUFfzW9pxeNkzaMBKxZXzbk/L6Fq9VrlFH0ShhUjGBj7VIyAuTmjNnFkeW/qpt82n1qATwIVDjt
G5FBfmTffPQsozL9yTV0u9APTed9nc3rtnIu9dKVi8XzvFFAGSkfOftd/49ii6xxNKd56RhOOOlt
Ut8Udx/e5xOwYSykTwhQt+3xNJW/9HTlXn9766mR68ZxYMc+7Lb0Nm6x+0wMZBfTgJuAM+E8BJ6v
TDFVVsTqP34wjzUQSu0UcQ6cxR+YrLhoa2R0hAH5N+uQ6Ps0YJXo3PwtM0xXjS8P/f4YJkLlLmI2
RF7CXJtadnNOnn6n51QM+YwbGsSYo0Vu1KVurV8OdCywhGk6GexB4vFR/1gCTzevH7D59tK2bqip
MBWvZU4944Jz+FsDtbtlh/FOZAbqOeEjLk/EVxfDEtCbWAf1EkW16AZ8ot37yYggGWvyihI72OSu
P/n1x8Bdrq5HIPGewkTwRDVfLhEVICkBGpOF2g8NAAUSva5L8ETdJUmNutvbWeaU6CW3wcVzjbio
hsgFaggQaMQmDXgju0Qgw0pFuzBL7TysDpuRg40LWCaGaYouEsk9ePnVVd1QcLX7eUQiv10/+til
ygbtPap+eDEQ3SJ+wzBHH51rXs82bxtu6E6fUZgEM1KaCqVKIH4w5XRYKJG5QpqgG5EgPErFwKbk
HTTori/BVCM2mzFXo6R+LFstA9XIEqosV7u16G219O7dgeV76PpVLPbM00aLO/LR6NJJxSz/qpYx
cYdfdUCsnUAJdrVbzhWo9Dvr3b3SuR/AE1wDvVjJGM0lZeER725vcWpffYVyRqsr3KESmZRWlV30
T2Ez4DeEFmABpy6aCOKmb7reOxdyP47EL1CQRUbUQ24c/3m5JTlIJHYYu54xNVdi0AxS8RUe/JA8
1sc6zfG+mWxlAPEJgPHD/d9tHj8Jir0dRyThrvG9W/jMSczQ6K12i7+rh/9yA/QyfNHnQlRJebzZ
eFjPI3QipTrrj+iItjZJfh6GM8Yqu5FUGO6WJMGHD0S/WvbpEbx7SxpWoMPYxRXjb7nSHWpcx+jt
o1qMN2R5boJkd4jycxtXKgamL7jlJbPrgFs1/Oriaq2j9ycjlxQt659MVcgQ1dsVoJ6zcfimoh2a
REHPm2xf1GRmZyYA3Lwaunxs3EC8VGkl0yVyPFe3YmDe/7RN8+UuSGSuX4bOyDmfxIt25lwhI+hU
e70KsjP5gHAgFQCPI8GXzaNpKZoiHkLSWKa+LPJKTTEls6etXkBZGWutsKZ4vC8OFYvR1m4HS8pi
PTDbHgL89Uczj9H+31VwAGVJX5rtnBmoY5iPxF6UTywKdV7Ib6fU4Z906ezcj06WZYNwgWI+Qw1U
SsGKcZG52ue6sV3NdawhANvQJ0H/lImrWxVqiMkGtUgEu3KNgqRj4A/zBUI52UsJDmtQA6HwILkm
zHYR4aiT66kWyyuTcM6+mgdsbmE8rhTYMG6YuX18QWEu7tNZ90HvcDcP595Ddl2+Zf7OmTjnGsGc
wwWAnK46eAsHt9//Cxjpu5USLl5V9otDMeSAypUhxKCY2LP+SUzrRICgsn7zg4BOWz633aPdD6DZ
x8/p4+as7fOEtuVJuAl2+GXoSQXXc5YkOsYcMJJcAVDbrwyXlTwy1svQ7HPz7cRkNCYaCsLQmQ0N
XQ7pHBCbsBEuNbu3FcAiB9q5W8QkL8Irdsqv/l15LgVj6mgzJn+syZO97NH2WyRG/AfGPcKcNLRl
+TVEN0cnEthSD42oiLPKET9MwmuAUVo+QSJ9+Zlde++UnjqIixs4x4qVLm/zs0p1ngkhrNE1VAeX
VHFYV8L3MnEUbmEYr3VS/PAhvNMfC6rYMMOESh0wKpGLAXLrwJWRr0+1ZOyxjAEdYMnxvHU4yFV5
i0CNdwAcZXx0ovauRlvpzMwWBJsH5KJtAhWlqPapkV4fbpA7NflFJn9ctvJ7vaaHts/2EmEwEQHx
0syBjjq5AwMMztbbuuNlF6TJnzeUEx5pmF+YSDtrpzQt+S/D8hzwuQd2gdF6fbDF3FKIoWQmV37s
/sgc6otsSOQcplyt4N2r2Cgq9v9GQppjKcM21PqcICY/B6E1P0TEvvjQzezK9RssJY/mS6N8v+qR
ypxEWsc5RODidbPcDH3GmNyEFjkba2KogpOT+iZ3oXB2aq74fb+SdxGTR4Pqo0CIvW4LpxK2OUCo
5YvGuuvna1OcDjfKTtkIjjC3mxD926fv9iZnwgckA/53ITcoo3dd/2cLWAuz2a4kiORXeUETVECl
a00zTmg9F3ciOE5otHOweI7PecZRQCSDUy4uMkxWAmg8JPZtXOCHJGlaEHZcofNiYnbitOq654mb
hBfXV1LDCwGA+aLbofEPuy9gnEKs7Oz6H5kVzrZBGaidPz3Qj3uJ5RLvvcWAOgUlMo2wnDaVB78p
IfchHmgmIyaD8MWJ++Ng3+WA9v133J6V5mgxaLRLpT1xfs+Wr1Mo7SrcO7p+G/2gYQOsQHvxkevG
/GT3SmyHvPp7Fh1HBmtDJ9aQcPlvfvCqCfbZSRxMb1hoW+/yu2sMBpCGGBQi2fW6KbLp6ZSwOvqw
Ml+s3sGgsIzVSgPyUlqpScPGekoOLIUJ3F0ayFnQMU+Pr6WHooO9xg8fItlT3fuPR9SmUSpxwcPW
A0XLmemJIAEBppajs21Se1Bz5VIwb3V+X1ng+WeIOhZbjycFyRNYSVcpBtxMv+VF3dQVXA7OlgmC
vDMR+Z19xv47Ecd1j+KEGc0RKdvnul/km2bCr39m/uYotK2fnUOLnXGyZCkX8OHga/pyQBNygJ4F
nTGU2SXsTA0hQeGQOX3fI4F3tXvbZXv9crwkr05lEHDKG1i+xJuUrEhBerv+4DYfSHuQ6A93y/UA
AjUaFKwPDLomAHmOgewCGwr0A7skgTdjtbnh1vi8mMgDud0etj/El3L2z/bzSP8msy2BsAHSSXTC
b6+Ioyy1AYyTmOK1v4bor7PRnbaXAF00Vn06UE7mO5ImfgBXURmpPQi1iWptbTTPsqKPY8lg54G0
i9HQtS5HOU6HO9LQqPF9On7hGEME1JnqinBI7n2Mg7Thv7RJYVJIF/j2+/hkkXnkRZzerFbwvZvy
C3u59yBY6WoqeLywTUAHXpirSbHg9kiwz+3OPajvvtIxTsDZI5m68OijwA65p3MYI8UHbyKIxyNT
uSkjzXDW8ZT9OfkSqckzWmPvR79S1V+jWmJ1QDOhHfnJ8kUHOYw0zCqXqmSfY6ZLa8FI2jsxthPD
dHLOvrvUPKDQLn3HoF+bMi1CR68enqbit7ZGYRfRGe0ott4YXPlCWDnLfCUPdUitKcKEwS+zIH2G
UMQPBNvaFJpnY/4gUsVCOf/krYHI4E38fwzrIrnOV68dYZ3dqpUM0+oJbfw0EC9Xo1iJ/hkgjUK1
aJmH+7HBzOvdhjaqrZdXzYsTx0yc9nSiYNQtPuFgyk1hUxBlLcEHzRiN0MiISUeaiKV4nxz/7h/V
JcYxe5KWqIB1iHIUxQILERIXMJko+PEej+gg6QOmP9c0+UrEznY96B5xNW2U6VEh7tLPVNEMr6Mo
dUmvfRaJjFMkT0nALlXNOE8gyXIDUS/Pq96chtXUMWC7zGF7UTDNxvyFbUC4rJYCwiHTzQaXIahQ
5BJPtSzPvXaAQ82dAS8nldwgohb6Wrzv8u4BsYNpcky4xfLQXR7cyD41lnjLB+hBV74/f+VNO8lL
sCa4ko6smoKE98H5WJpxJGwomtIjxF/QDhKD5tLMHbtPZudGdRyr8Xl5+xqwGz8mOVwDrGG3XJpy
AsOWLQe9xFyRn2J7crewJBf2/t27t1LawVr0gWl2LMa9F3NFLIHS4cbtSG+DFx6sGTsw3awal0yr
htHY16/ebTOfDGaZkO/GXxkktXaTzgE2OT+sRsaYMdev6+agQyaCSTVAFGLUfi2ZCVEo1xfSuPur
kDpMIeKMWknoxsbziDowuzxAt47rL6dT3mOhHL3sqvUR+ApGBdAPUz2Qa2ngot3822dZTeXUgtzJ
tiwale56u+Pr6vkUYKZjIghxFvy7y9MAkI5UzwL12FOKlKoygwy78cjqcL+br9UAFQEW6tTz7A2R
G7nNoT+8RwBMUCQclZyhZTwUQP/U1Z4rd5G+uhckMgXeXgFC1J9KOiwRfSkoDVT5GIKzSj0dX9tk
kt1cWFZzC7a+h2djIg6FpubPBOwismkLk64mwwPnlzKLEvOm4XKyjQN+5W5B8eXcUORK7PuWaYWd
G2Kvlyq1BHUe06X7gwqA4EZiHAd51aXPNihuc9gfhIsckS2S2Ttpjf1Kh4LmFwS25ikZaM85fzKh
/pkQ7UFJxu6IV6DHvYRIsv+KI7IMyFHZzKiH5REHdQ/qCKW92IZdo5st8rW/PEgbm9hilJMDLoy5
wfMdULKDQ5nPoVlUkFXAXPag88ykILnNUsRbvHZKTEKQe2zB883Gq0mtkRjjxYwGmyRGGaMnxw+5
B9h5LRAdnXBDQ+vZuq8ABPqNZtg54Bb9yd0cRj1swuylGHJapp8VhhMj/HviOiI5OBvh6UkzRSLY
QV/JXHnjP5MFqFkxw3ZX5zkBf+QBBOpGDsQjJVHR/QubFrUyEG9iZM42lSTTJQLliDHRmSRhvWM8
MS/k8TIEICFHu95T/u+RX15TnGLkxb6bm055Tx8WE2vnH+HjBSkerHbutvULRMRoLMRSq3yuEMgt
QpooRugVlwTD0qeoLJFhW0cv1/cuPer9p7Nti4fUwQFKUXmDKUo9RGKhobqHaECOkXawsQrezimu
x7clktQPNVBqef99IIZb/t5SSVK0FyWZxqbFZjOpMpUGONLA4QeGBbKMk/js2u+TdKfwjWuJ2Zb5
ov/Z75x618fwWRXaFE7t00pGXPO4MQBm6MlDISdcpstlMjd92mqPgjXlVPoSjP/ZtpdNx0naiiJV
numW/2f/oa+R+L6q0tC5aY1Qf76zPYKUVGLg7tiEMQGXi1QXqvWX3j+PByZ1JByd7NLLP6pSh//d
WAgsTKpN5UoGGjesBhSVz0OLrVXGJtjPaSM8JN+ARvrYEDL/VerNSYXwV5Vg55weq1EzhEh8at1L
G+Vfo0iv4oyT/dOc5m2/ednbff7No6Q6UKVCZLIfsJS4QDV6urV4oiczwcCf9oQTCZusaPghI8I2
I0RVc0eZO9qhmcYlpnrQUXs2Gthb2eTFcX+bmyPT3dfwt3CTCtuoEIYdLBeZLMfH+NMHnapXOKtc
Bvx3pEh4ZDQtn8IXojRYQMgKxxk+/5Ll8emNR5vrdPkAMDvI4Uw/F+wmC+refv0twqvZ1Ib1MnLI
up6JKFDTvYaG92rBmGJku6JPi86LKgQVdMgP1Qw2oGSenw8ohbg3UoEbCz+kFMPo3Ykyw6ZPwIoF
9pdPZiMUMK0u3gFnR4xkylNrirmCWx/PId78Nh828f0Ks/hYyiMhiLC+DQE1v1FRQOy7PAu1UTuZ
G1qA+D5m4+cLetkrPsVxPbuJ0IYiJgV5mMTiY0eZCgR4xCnDdd0fBLWZ30dTyG2tygvQ+bZq9N6V
q6OyFOqaamVGYTp9PkgaYLGl+A6EaO8ooX2GSNGjbcHYMaW+ikn0jfzXqj9CHTw67bkiMvLyAdvL
JSLwxN+ASGlfNEQGBXUb0jd+rcWgQoHC6/oJXX+qugPj4NdcInX4vjLkIrb4Fu6ySjc7VlBONYaZ
D6Nu8gAwPe7KjUEKYCkJsGlY1OnEwTw/QusPwulScY1WYOts9T2WKSFTiry/ZE6xLxT3pW/FfnAK
JPBzLuRZQBqC/Dzdfp/4hZYrWBlVw4CSDZXHJR9goI6e6IulfnhsMNxs4fW8ODL6CSMKcxzOQsvC
bcn75W1bzqUt9SuewJtAJZa/xIGoxwZDG/qD/U4aVE1oCaGIhjripdCFtlUPfxf+TL6HYFZURmjw
3n+fvhMJPJIgKlN6ebqTGE4Ef3vSsMGxt+nIsW8itR+iSZGZ/rpVXk22yktqrirLVyAFc3+bM0ZI
r+AlkXiTDONRwWSbNBdlPPLaXhjPHElCHKkgTx6VDnWzDXPikeNAWY9aAFkbnUC9kkHF4TDqSFI2
QaBzFXGmhv5n8hDKfD0S/izlotkc6Uf+A6o4XmJYu4tjhoywsc3laHYF+2ZfPqU6Sv0bNyfyjt3Q
hG/8O2uD0E/vcZEKA/KIqpIfoH5yOpx53KzZOFUjXN0LJi3okqHmTIrsTfhI6Sq7ijVBle3LwiOs
vV2Q3CRon88/1YHCHnRAPOsSCHsQJueJDJN5anLtzolanSM/Ac7G2MVJ749JF7ZajHpoNOF9Ig+N
jjiaReWUpbP+vmn2/5tD5iyPE/5LnezUIVd969qAwFX3yySIxaa63L+M5sPtVmcANQbHLmITIlXy
D351kumH7HEJagnol4b3l5sMUzyi/hy1OtNx/7FVH/WhW4TSSRbKvXevkhchv4zevQF6Wf2DKqC3
qAIGLIzM+pe3YKMU+PU4ThCNgl9SNeFwdRRgdTAbtJkLR6Lz+6K3kVxIXxKQ1atU8WirT/wvyzwg
S7Nf+Kh517mL+z9UJdFks5KgBlnEq8QxR7K+ggauCn3t6qXTYrFbnt70nZydmEXjjxFI31EmAKnc
7u/0IUQghg0S79/grwnLGe/aRscW+zuY7dpeQ3oGG06GftJUVWEY0TGqsQnhGFrFhvSZf1F/mK8b
HPrAFeStxXKmJNX4ju6mq8aRB2fIxnCFSgwwAscvSy32E+mUksl1KlzpNSLrqWb2LSP+9yoCoTXx
NFd8AYs9tNuFEN2F68JkCRqxCMsI2co0HVaU3bVEdMDfdW4prK44oy7S+xPsPTJnu0CYwoHe34Yg
wECCJy8PqzPZx7SoLCG8Ad6vhPcWc3OxtBVYbWI93AFbB+HLe7EYcW7AFrm6TnUaoniIRfYa31e9
6EzilocVRbkquLrHdRyqhP3TBgnGhyEy9fdng268t6Dl2oMYWMzfPIA7r98f3dZXoudBUuFwhnD9
QIQbqR4UvO+L3V0+pWfKSqnOtQZwZ3fRXUa5hOv5CpTnwql+9SuBKZtYlwD99Rhf46D9X44g3rPk
RGnFsyfqK/G0w1YOv5ad8sgPbj19Ihkb+9SPPl9tcRxawLcFpTAclhrwf0bPGovK63qm4Gtc0XCN
+ZUpHiJ6chD5V3IQG4V9hrYi65dnqCNdrmYIGhCNUGQS8ZrAx0KSjn7eAtDr9DupCJmavYl+oG7V
uwoLCsuV8xWiVMO+pyCr8akqDDodSW9qavceOwiq4iVyvxjmuS4GoF9iypyLEtE3nZe9tgK3SBqr
KHP0C0MCbDFz2il5zcMISwBf8t+88uq7JP3sE7c78LGkbzkIZCgz/nAV4Sm1tfIOuwXAfAjG9ZpB
itrNpGwCabmD3i4IoZn1wLbjLQ0ROG4lApnf4JmXkgSN3cRLi7typ4P1HKLPDueexB+RmsZTp7o6
tXWJbh41CACJEts1KfYP2UHpsZJ39DGrQozHoMIwIRH+LZBOKn6HmUY2tyxgwfIBvvuV63XTE3Ak
3OSVckuZ7ImQWh4wkc9RBv8mtE8jhBeTIsy5q1AhZO8sG/lk55CzpTvPd9/qO9qBd3UpeQvpt0yV
n52QtnuxuXvY2j0cLNEzUChU01zYSjmgAB75p49gTKslaMrJt35E2G8y4L5Sd7z+Uk38UkHulRZ3
w/JpRIr5+4zrUFjyD0ZxvFZUxDUS9obZVLoADzfwCOBeNiHcQYUGPiFa3DP3gOTYt01AwPNx9SMe
BAWISxm0IgHWBnEisPllmUIhy4cQCnXw6At2IoaI3X4OYlQOjM35u+DZ+rxg7ZKeLoP4UYKKXwOd
e7q0MEeKBqG2wOWCDoceinKoOI4GaKDRNVyly1hVnWlSwGxK+YF6ljKpbTLN/edphFB5yTe2BLmb
Pqb/ED/ar4ytFHJj11HjVRzD1rq61EVqlLSAhvVV5cP3XwlVr6wPZV6u2vEoJTIQvGRfEpZbsR27
jEYRbjOqzhpER2AXUyiyk06TEcELgKwcT0/dMgLUDxcy1/TFmhSgvnzVy1OPMCrt/3To2nOSsrAQ
Y0FT6qD9/x4F88ouQ74249ZCHXSNocuEdUMuYI1Q9yDg2zUJSoukfn5QjhGcgrFGPXl/ZDchaS+U
RK0v44PXnX5xmCt1ob5jU03uD7M1gKBRwFkwn45J2pU27/YqKqsEr3qXQmPtxZ9zNlb0eHQhmTcT
UlvGGmWTaJSR6mbKKOOD4OakVIuqNlLdwYJF6Y8Xz5lV0CtQ2DJTwYEhfbVDb5Br3vwMEf6N4X9x
3qV4ghvM6QfvDZExmhrpA4EwdCqicEBd9i/ba4g/qbmNPKV5fQPEZmZILukqYJL5SDmlUKAbzC61
oK28ep2GY/OUyrRbW3Cr2FiyjnWlyT3lx5VfkvF7lpRXiKILlE8/hq0/5S2tn5MPTRkBdHct2APf
N7aVK25baJ3DVuUXK0rrmBK8ZRTh+s++4j6tyNX7NtbFeUqrZ3jv6rnVJhNmXCs89uL7ZQJbb4bo
4cBEDipQRc2NEGTKhI5cOVTRv/tOH1n8XzA3RPeGs7828DR6z3T60zDHh4EWiT+xB93Cu2S9wUF4
NPAvS4ghIqy7ydBBLcTS4p2nEspbvk9cZsEeTN4SM2tx5JTAcoT+IICPN8vLMR9LrtbuKY5ybDCo
4DvZT9O5d/FypwxtglKY0Z/V+tP82dtfqIK5o0tsvOcxRBJgYA6q/Fmf5ORBe41ShCcQwmbTOJTw
UNZB2t3Efj6EBC3qod6VmfI+9p3LduYSVoLZPwXURAWzV2LkAT6m1P25+VcySgdr8k7KU/H0+0Cv
Q1yisLfiLCAzln5lzI/JANniYBhITQauMs2GWd0EODNVMp9X2PRCIxzi+TUsxX+f77atfFvhlGFv
8LckiLZ6pdn336vysS11mB0plgX/IprHZE1phK6fvGGJ9QaCHjzMG1AfYYJOmbWE2W18Qd/AIrOj
TH/vYJ/Jdg51i5xJyjDFJ0Q0TzNT+Zzl3AvlrphFqytfBi+erLGGK90azZ4csYqdxfGrBOehxZXX
kkCAA4hMmpbVIbVkEy407fMRcXTOrBqzp/cvXURvv7iotwNrb4wDEzW97f37UGUL1rpQ1tglnLru
qJx6CGy/WLVCy58E65+kXBFR2z74l0UwmsswJ6i4AOtQ+P5LM8P2LDLhdAJ8EvPHLhHoiH5RP+jz
qqM0pQIanzk7HXRBov34wB/oyYaKM7F9XtFzRqb2D4ixkv/0O7ux8sltQQM+FCwQ+8xjQC25Of4m
j0xgwhybbwpdpdUa3mAnSTYrtKGRmkOuhqmS8x3vFzfSqL/kEtX2N75YA0O8hPmNzPSBxaLA06rN
w6GULfd+Xm/VLuhRE5QiGJN+sAXSXVqMe7w1UteLXHZVRMeWGPeMXbA/wY2RyX6p0VbFkfAa4AmD
Cnzljl+49cX/nmP3NTwJXSk3blMifnklIsumX3d0jKaiQyzTy02iLksZKjzDQsiflDwmiuVqfOLf
9KvS1E1VZUj4AsCpupYbO2BCnvgu2YLleJ+FKp8CUKYY7V4oSEQZNBTbauDPURT9UC7w9uY2l7X6
qWx0eNP1jSwuk0JTGpexfMHB/XcQ7rhAsZOkSPlERb/U1lA3+dguBZDs29018xXonEHTRbrTapEh
f21LBVsabTmzvFXBpW1tC3sFp4v+XRZCSAx3IDEmsaVovAigxc5w1z/UroyzCHJxTGSFbXLUK7bt
nuYEJRUBbpvAJEmJEh20ptIxYmKFjdhU5OTTT8IFdWR1mpe1ZryPiCuSOuHXMsZGb8E/QWYHfHRX
39piHETZOh0QfGZkAfcENKIiyf99efhw94YNTcbVLILV+PHN63QqwNaCr06mMNglj2nIkuRTbn88
mwN4d15dwEBYcFIhTai/qbWrIV9k9a12cl+KwJzjToU+6we/TG8SN6+NGzvGvAcsHbqSYplhTAr4
mK3Ps1TiDx0ASwaooIzd0opn63sWQjsz8aQrnRcMgmXlzrM6WR1hWbhgBN23Ljyx0qmJaAmjayYy
IgeYZMEFNqfRJy+ucPq97i/3R4GNp46qsef+G8pyzvpm98rm6AsTslcWb1cnQ4v64qFdNuoDOjtB
gS9SJV5APqOkIVJmbBnPBoxZ+obrY1UvAEgaq7L3uxU2SkJ1lnV+tgohylSfEpjwwW7bdZEb7iqR
uQ0oFWYx5P74kF/mbhsq64qMTuvh5UZoX4AozcUuHdYUIlBsUKJudneKPhbcQ+E6dlM+TC/hKDkD
wTBmwF20w9HFJ8rKoFW+GXSbS83r5yNqMSjxWOwQ52KWClpg+K00JeZzzgaAzSc4+kqSR6nbecrp
sYOLMMMM5Bqis4Cws5e+OYJbIYVek66NbkUb8fvxeaGrBe7CBJ6T4FVSQ1EJtwi6k5INEaMKwIK4
YxCen8YmvuJpY2J+zNJOen1o6kVNIeS2jG5fUj2xzVBtsSV5lS5FID+vAVa+gCYbb3Yp+pRa29BN
r9vcPNiutPZ16A99UD/eioMg+RtL/tL3Ett8d23WfN/JL6QkJALwYnV1mrLQFHwROagGSxL52e96
eC1Il0VskWFIAvTlFJcvdxQ4gRnBQlsZPSBu/h3atsiXWsRj8CDfYCqH4heyZyt7P65Ok/b5aazL
pfNB9hNL43lhHUlT+YDPU5uZO7fEJ6AXY139iJeSCSB7Nbht3V5W1KwCFGAOGJe2T/va5vWVb9Fd
ZwFfCuqYmiYIwduvK5a8sUXCBY2xi6RoxYWdEiN2jXJOZ/jmJfMutfHbyMKj3EVexy7t2l3eORsx
ySqMWyG5VXZzyrU9/HBkzrCa0T5pgw9ogrJzt31QMoeJYRgMuGtaQI0hQsRaLOsLbLNbr7Co7oo1
zWc860OUWr6BgXA/Lvk1Lw/+oN0RoUjDYrTRjiX+MkQ11IKtKT8X/S3+1qF/v1WCpEKMt0Gzncwq
eKNalhK3vBoy6hQh/+Vx86bw+z6lYyMS3oYBaTEwriiQji8/Yg6Pq7s31lP1O8Va2SMTF/rGnLoF
Ec8py3nS2+5Il8SYcFwn26OetmTl8pTnMg3ib8bvGQSfpa+YbYpNV4uBVe7HDFsg+Q7zvN8qiJIN
4ZOR5fCJ972rNxCWzgiOYcwo/OcmWuUX57RHXpQFOY6JN1jY9BzREyhbJ0NU/jMZYj641UP1uuaO
6ZTTjSVxU/ZBePO10GfFrfC/npevgiVYs+2lOHforJ1uObw9y1Lha4ZbWvrvKOQ3Qfko44utXYyS
7weJ9u0TstlVMZ+ntGIqb39TA/tE18nQusnqtAMn0MOozzLEzacwdYMJh5iIQb0/emJnxKo6w0hY
JbVgPGJTkHekATRN3lTBr5xk68QRBFAShVGyT1OzekLiDurVJTWt+dL29FstKsEa5v7CgFYcQJ9S
k7EDjI6h554o3xZ0z7jPeiYn3BEWXcb/ugQjbxihNoGdlo8mMPAHtmi75t5r/RBZUwZutPJUCA2e
IE3SudWzzLNuR1/3jwdLsVZ1AREKs61KMf2NJ21XCSNWobiXtsiGXZHvOxBgpzVyGfPOueehAH/G
cx6H24Dg/poUJRmqq3fTmDilbfwOEh76hhrVwkizZuj7slxc0ryaXb23WpvJDrtJ9ZIP1yFDaGGy
UjGPyh1BtuSB7cpLybwywCQtA0U/YWk74IPieT0LZXhJ3r29PNfki6ayclIKT7vt8PiYXQ7xXCoI
Fk7RYT+qIAY0E4hYjn/+nmUZJYxrTLYl39qw38JNUFrwh7SM18UOE5Uppt5HDtiW1/+CVpW9TJX3
dhunDA4iQEEZcYM2NMht6WZgxyxj8rNYOwFbxIasx/63igsfqnIyWhO4qh0pwvz9GlFcg9w1rawf
W8ivwlnqSdmurcipCtF8OuYl1aXk2spp98yPmG+9oKjfTO3UuttLrXCEO6CahaZWRYCYIFFJw7+Y
lAUIyJRyZ6qKb3XW0HplnfJazWcoTBXdWmZ8vYFH+MTG0o9/ZS5PcQ03+9C7HyIUb9dGktDLkIsR
0tbbFgKXd58A27v0/BUE43pYIQZudYdsPOZjdHfES9TUfHcpeejRfhROrnWLPFVCq7i140ruzaV7
OCkQ4BqhlpkP2QZk6yJBKhEu0gRtQLXZ1bzLafNYDGGAbPCQpLdQnO5s+wktk5jSYuD6QhUDetgO
+qcbXb4+0k0ah6/y+k8EX3V8KHTwwB5rK10rh3VaObQ+3kr3AMqarpVfTRFfDwSJkRgmpo1eD42W
7XmwjOjnaUqHSg7XUAA0ias/ETfB4LHZdkfDztrkiPPzOXEI1HJ18ig8A9PH1PWeNoU6V6x3nAUO
rH0wosdwSMdKEQvsdljXGKSF3j/2BbLSyzVdqa388rr25zBGkNdx7UhQx5Sfw3XX+BVVcJiv97qo
F1mPFxi2uGTzebWxcIluhn7B+OCjb92UbkN58r0PxZ1NZz5nNIqh484O0xm/Rx8+OzPole+XfcKQ
7oS+PM/5KjOHW+dTJR5UjSE+9ERXZfomIxpK6c3wq36yU3D0o82+BZDxKnN2VKb+/jS18bpLfdfV
aazy/mce9BiNWuQeo7Fff0UFCtpXQm+x8M7nyUpcSdOPf5MnstlPxXSetGRPmjO8wpAiAAnfOmpd
wdN9tiwKKLRHp+NVfq9EZhL8UgVxbLeJg/Y45r41tmxN1yp2kXHqyuzT45XVNhIaubU0a9bDOvCv
u0yppnMeXnQ/0FPvIQlVyU1wkSdowwkSCf6gEgCrePwxbPN8a1CVF/JtoNFs3jW4ZLoDgrImLJ+i
+B/XanzJx2WrheWy3fClTn+oaviLVU8LpQZLC5YOQDWEgQBuGDPfLZ6zGDsXNDqI2nEvkksrG3Ut
t+e5mhvV9iHqR7BDq01eF+nKKci4IztzBuHYRvtXt4F3ZBegwbluRIyPPr/nZX3zkTvyRQxSW1SX
q7pafNq+XiAo+h9bFs57UzgvS/kL8/jEfhD1qDxeLGe3ZTQueWfcC1SY//em18iho1OzcY0vW1BS
V1uxlXs1PyPLAYu3u2+lTQOtX2jS6NBPzcnGuqyd557BtfTikjmIydTdNE9NznT7aDAp6rK4n+Tv
MagMCzc+IEYPVpCJnFsVJhQMPqPOsIrWud5IhyqnEoY6G5k4JIFLlBs27IgTqKobA59lB6raiS4w
tQQU0DAozQHVxtpuy89qhfC9j+v8ULZuw6hcgKMAZ8G+UtmMl5HCyCcrd4dQ9qA7oREfqYVATMUP
fGkhw3lc5pmPK9MFVa3T1Btl0GhCVvxrLFTtWgmjgTI+CfsQrRWU4JBuwX9qhiRPiyURNuRUlO5Y
23xUjviITeBdYbNuBzMrQ2Ix0yBkYxRes+uf+FMkfoUuIHRe4z+5CRxRu5x4TTATJAjRv2Yt8trl
qlD1pqw4zDVaViqXvca55RR/DAugnHJG+k/d9kIBp0GPhPW5A/B4+dodFUET8HRMERfFX1YqN6FA
tXG2LmM5VrWdlyaiIlVzAleh6SaSMuYLGfwapHqr+IPmfy3yCWqpb9PFAVbRUstzCEXrHBiecNtg
L8A44BxGYYtWUR5/iiwIoIaao3j8Ns4vdWcqUSwNb333D07FEOAXlMCo2d07gbddI/P6YhlJUerD
bt7hE6pPfEIlqZ/F6YhvprsSykr97l+KLXSoHOT65umuCLHTVlOBGMsZ/oSwLmbiwTQYSydjHZlN
y99qBB33UNZlKRYdl6uwAnAC3QCRZG4pt9fM1J5vOzi+MOHh/0zkUAalL5WwRJ8DH4HVZKtxg/mz
XrzwOrJaM/ueg4aY1BDiaUv++CoRA+PfSU1fk5E2LNkT/GGQkv1r23nqv6v+y6/3ociN7cOVXMyJ
oKgM5EZNITas39P9A0w+FwhDmPHYKJpcfDdg/0U0bljdp2MO5N/65HNC+WtL02LeCzzToOvXNXi/
sVFxzM/rykCX8BpXq/kOCUQKCAlyUwm9DK6WVF53LLaHVmlRnbB1fi2f1w0XSU8geI3BQu6GRaFv
t+y/jICIVldGsr29e+O89DngiRYMaFDL4nmO/kd9J+kZs9eIowSTrRKMAZFmroTkpJ5bNtmpKEBa
5sb3Zom/Wzg8mHy0hYLbEo5ngykn6LJu5GjT46zTcV7p6esQNgzNRoNHQx0628k64uYPrNiIpgoy
DHv5j6kUQPpGMyvJaDobl0ySYoKmjqFszqWlK3u2WZWiHvelmTZU/U+2423U+4oewRZE7DqPGpbj
rL9U+bQ5feVSY+c91YeLbuGePJ0tk4XOt2gvEBmXpG4yWG08gumttohLQ4fVBp23rj6cBPoHzMBf
E/UUYEgrPj6T/qu101RVoCDZfUe+RgDlhnhxmuV35/JmeM/6mxFZ+uiyznbDLhOxtIlzW+exuA63
Vc5fKapx5d5zvkpt/dqHOzJRMBgFnZ/KkV9W/TdMxjiIOFUKmDNzVoeDDWx5VKRY1jc1jgIhqHlv
D/tY35YwSOE5x0PrkE9ndVH4apQfOw3UyVvoVgFBJPSsv9w6WJcB+w5stVMnEobRzp9fVOIwcUth
ifsEg/eDkIY0AvG/VxCj47KgWQWnFVzbDzm0QAUkgm4ZiYX13sz8cinz31FKqNY8Jh5KkSTByTxt
FWFC93ZCoCR8tH1amf1phwAyttjcOVpLwPJOmd746qqzccIrwDQzpFyw0lwD6jSLMDLLGBnN8Nqb
TFGTsFL/htN+YycfPTc5Qm4bcI/unkAmqn3GoeNyF0I0hcBzV1t179D+buYDVi2iITqe48MNbZC/
OzTPW4Nzol2fvTEETZUUVUqGf8AK3UKmxWMX+OQQ3aV3E/KwmY5c0elLcdWoSyKb4onM612eePfP
1XOMY+RKCHV8LOZn4O/MVDd+HgpHtl9LuplD8aEWzs/vRLRNgedxen20fxXpCC3TEbUSBpa2f8V6
21f5G+lMTOyZ600SreS0YjmYd6FGH0Tzy/D9lGWDRdoWtp+4Gt96Cnffph07L7EHOJ/lRMX/Q4bD
Md/YuE/dT2EbID264QpNJSe7hZOZvdE4kDY+Y89DMR3aLYzjp+uTSa+uKaU0Q3aLC9M5c/6EiwhW
WFPgDuPPHDxkmpklWp73VxTXS98fqWY+ox1NF8ew3X03Pn5D4YPVtG6flsE9wOHD3TiMxsRAk4QC
ucvBk7fdJq66dUG5lSmw5qm1zV+sYRxsKxFMik7iuMbiEvJVWsvsIoLXvUfNHJswVVXkBG8n2y7V
Fe7NMzp8PCRcTaUVZsCjX+KmaeDxFO+vfd8u0hUxAbr7g6Eysvzqa2IE9DjUPz5YQ0/nVioKmxyN
szPBAQnOBNGcBtZqwu25LDQC3D1OUuJbctNwE9O9pNjJ6cCBdPKiFn8N4W0RTuuXCmWgYt5RQtpN
Vm5fFWkpW7DihirTXs1vjHOGsT1MkvmFBFUzBlzJd6j4NAwS379EheqzQc3w6GjggRiHlT7gh8Hy
+UKxYUN6nrTXe/gHsRT9+LZJ7gsrrD9zWr+lWKOleLeedDXgQAYL/qdsUpjNZv3Xt97iHOSIGXPA
uuY8t76AK5omSnxKVQJT97BA+/nJYeGxaAkYvCgRg0KCVG9E59QMkobkHbkO8m673epNap3qTND4
DdS4CIFCW6GFJlMc2spZM8gK4M9gKWHdlh6legTLgOKgqI8ca044bChThAHlPRhLI5X4QAywDUk8
WqmFMN5GVbfnaLrSlH1j4CrmQM+eI6P8nTI5tLvPGl/gh7f2c4FQYhIPGUxKP4+/DfYg2TpAtd0i
16X2S9gxRyKj5La8mPcQs/xMYPFFC1H2XsD5DHbNvhHapgpgD0uyrsrDAg6h9Qj7QFPUQUVDBj8K
bW8VajPtw4/ndoTYLWG6Zt428BazzePGHpkX3J6yywpBQ82dnkD8sMKe7tPdhgwxVS5gqjPlqbSV
D0u9SU3nvTR4oX9eFvEeAaHR8IiUh8Lq9/flcy+lfSaKYwHlt+Hyn54ISKG0p1fztRP2v38B+L8M
S51h1qYJwgVMCssH5jY/3Pd/2pX1C8zKb6ouzzN3s9j9nyqym1a4NGW4PV40ir9ZSWQuPnHCKBzg
5TTwR2uTlJ+ssnS5BXjapZXJIQJ20mwvG8g1QIzWBOKMjNMt4Ps9Q8TP8Xuov4Zy3tCdfRmvAs4c
rvUmsXdAbuYP0vNFRCpyq8j+y0kp5YALcsXCKGXzKFXnutL4f1cmuadfrZfwTBAS3oMqW7sRAz+P
bPUQ70HAoXN6706HakYWL+XhMz8dNndueCwvUSc7lTMRCgmtjVd7JBaKZB01K7qGnNwzC34ft3xb
HdhieLVTQBPN+/o7K954DcqFBAMxjtu2gz6imDz+ePcTxTx3mDyHJTkq+wJfheYaMXXyahDtCS6P
ekyFinzyDH8XLCP6+UHBAF+Ad3j4pyHi/1Lpm88p4GkxbjytGa6/18bGxRrOxJJkdcFHCoIiWYcM
Qur9EXgGtb4C0tAWejXFBFjG1PK0FcmNmF2UUcvOu8CSIx8fkyJtAUY2WkQHlfUOb93zGGyma+pf
lhU17KM8l1ZzfcrVkfie4xpszM8IjSwpO1JwquwlbAzjcCpbrItwjZ9CUEYO6SUoXMhZJdFEFB4Y
NFYg4oaQf17uGvXhnSwqTr1ES11IwrG3I8LnadeYRIlThipSup2iH+ZbtTtPNHNTgCkYhUZLO72L
q7oZ9O3FELx2PnH42ePMp9XKlmU+wS4OSZIAvl1rdXQHtcaqVmQo52u6HHWYm38ehem9cz/y55Gi
m9uzES94KMjnrtCNeuY75P+CnilAqIbSUaLQ/36Cq/hDB2tlDHm2Hqd0aK9GQeT8oxX8zPNrVixC
YM5iQoc42HoJULTgzYFzDL8FwLtCWRvdAmtxY+O8g2d/h0bvc73gNgoF/Eu8eXECdiM9dn6b10w8
wset2TTsSBMUJMwH7oJdzejnjIUaKeNf+M3SCT2B2GqZmqU3WH9VgnVC5RkLNnWhhZKV0JjQqfFK
q1ci+WbzGFwst5z9TKo1jCeJ1ojCOihv/zvbceqFoqOz/yViIJRZIKCDHxIJ2rtnfhZNQ7YTIVKR
bPdS7WjlTh5jPF+waGf5Xs+5ltTuhsBSDyqO6Z3TTSTTiDFLRnK42YetaKXCafswVI0V+yP21qOR
2cc6ePVXbfZKz7Qw8/dd75w0CmnPmb+3JCVKxkjTRN8zBbdVQKYPTjSbnCNaLYzq94G7ByN1lRCf
pUxHHLLMpjwpRpBcn7ees0G1w0uky4Y1v4bqt2YCtXvTl3K8jdCDwNig1ZuFpBCAqOz3HmtWCbLs
cxDq8CsYi+b7P5ddkbSDE360RIUbB2puIfyrA7qvh7M+SRmZDapCXW8WIM5CNUFBBM9A8aSpFeWW
yEUG8BOYc65sQVXubQFGzLzAyYguN2wJYqg0Wpwd1LnEXgGQWIxVfedOJ8z5NwftQR+fdoMHDYkg
MstYl0DMeJxQEecTR37RRzKtDwYKyWob7uKSwMVCTn4SaPEdUxP6gtN3KGj9rFVmevZEHPFb50N6
CnRqhfDlKNVNpKdQyoSR0/2KHziEHCyyr7kz0Cvq0gNlHVH02S1N99kGwjjakLSTHHDX0Zk0c/DT
1ma92qNdI7eEIWtjMN3sIqMkubBSq18AqJ4sNphLtfKEDi+aNvdVr13Lr3EQnq7U2CYi0UmTXhgk
QHnGgI8YJ8n5wsk9yG/aXelKF0YDv2ZJsMlY+8TpoN6FM1BpYM3u4O/7KYyS7JWa3SK3Wx5/qMQR
ZJomFllvlxeULFqo7dfAUeA8V8+swJTVI4dr9EwVwXtI5u9+p7m1VhLCtuW20wvAixR3eboEOeg1
XGpwnbpVlZOuqaA2QsPbzmnu3buC33847xZR1PJw/3HJ9vo96AtgXJdg4r9hxIbvR40oowkngTiD
6g82dqXk/MEmEGbxeqb2MhFL5Ahw7mxFweybhTd1cSKGo1Yw/suKRiBJLnKIkv/ZJAxb4SIKaw4s
IVfcpYHLL3EgmQ4oBgeM6C3WqUfiqIshKHGACse92A4Dm6R3H7c7I1uBr++j3ci1t4k1julZxZrb
O5bRUAp/wLigApk025cS9f5oPixUU+d4JYk/Izlpu0WxEvQG63tKUBFU4vJYgv72PVvxdSEaXlds
GN0MZOQGv1nMrPTnUZzFURxzuqW0qISj1eGuXzXV8PumCrW5njFRSeeoLKeND7EEZQ8TldRDX3ck
nq4bSRrv93b290nj3Ed/MX8UOwbBYFdQiCQlVM2lWO1roS/+MJCPTsfXcYy0SREWL0fwSstz7QDi
e1inzdVsNuIKY6wTV7KCjKAa6S/Z4oebQZPAAhkPv4YB69j7zGOe0p8NJ8bjEuSzaz9suSyuy5hp
jNQmyf4eMMFCSBhirAHv10zo+mt6YjKWD72uFxUmO307DiEUtt3Hm3esjftMNGGqJJoD0FlDEnYb
cPyd1zcuS4iyv0xYGJUpn6DeArK47ORnGTA5aOwYoa9Z6HOqZ4lqnFhWpFG6xBzNr78uVUuHEwkc
5CT/vHPRP1YBDBkNZt4HIHPd1OflIqP6qpYtFx+N4ZLTaiouKCwBuskJxXRRSOTdCbSQufNYwB+m
Lz65lbMj/Il1NMxKuzQ6n9LfDn2B5jaMrIq1xVmhULbs7s27MSBhz6tuW9T1bSHIMfVlFx0xG0Wv
vZ4sMSy05FYep+sreoEC+v2RZKb9odn5nWDo2s7lno65+Dwn8Yfekjs2wrIRwmAKkcH4jsBsXhbz
s+vlAiV87LLhj/Rd3TwFwbBpF5aARtMuDiAUTSypad2tTMJ+qUjwfbs1tYEBAflxVYLRpMrOXnr7
0cCUBErOdCQkGxBEvHOCBzufHqv5Ja+HxavvdOq5Cz08HafWYH3HAAGUt0IZdmRQMV6K7RZMqprM
uxGPd/TjedoF1Zj6EfrXxUomdqbjxwgXOMDCBpiaD/g6po55TqBcQICJ8eygRFDHKxiTw+kPbXra
BD+N5n8QSQ9FlrPMM6H0eIth3BtvAhYbsvsgIhv9QcMlpJPNwCjWHm7Y2Y6jVRtVz/SKJ7m8r4zi
fuFe8Z6kAkp2iklLQlcyw8Sg8LxwRch6b7pO3EWaCXoeVZa32hBh24LHzs/orQPEZ9b1eIW9WFOR
XIZejrArYP+bGGPvkLTOvvaq9q1EMQX+RvvocqlEM60Uob1zYe9qPKLSX9F+NU1EFm/eo9eu3itI
ts/2/+dLiosfaxYJv7Mn2tQJkdYqwPdURN8qmTUfXx1F/6hJCKA0SjjPmZUavj+/x3O99NvXzD0W
ZOGUBReQLwZH/XOeWM39BG8p6u3Px3whHwLeVe/rFSEnW5Ho1lAp6+lHsym7s75WoBN/SvRNh4ug
Liii3+kHH3reVWX/ZTTmld9v9lA6G5kioIih4kVdAQ4CPLWva9P/UvFYwx4j/t4JsKbRr9zbfkOq
gAeNekuGCB4Y7NB6s+4W4GQz+nONcP3wB6A/dCZTXw7kVLMfrG7bo9ALSnYPeHicJUv8nvcFtz/9
osmVL7SQO1xruFDvGPIy13fQuR3tkfbpmNphXELkWcM1xLGCsQnZ0POdwcSwk7XkUsUJODy6F0br
iU35NSGLbrAZeaUpaeTxXB5fxPQpowWZv8VvI+uw52C3srbt2/kA2R4VVdwoea1BuSjWq6k24s07
+oZT9vAAiEC2IgOa/ZxjxG8380dPWwrSBUPY/bH+kIcJJkDpj0Fd0oHIwR38i75IJFTNDph8ZXLG
Pt240FwUXJjk+ewKx11O9gPNVPwu1QQTUg+YdBu6g3fssrgwVnP4Z1hVSOPFoI2nQKDGvpywjhFs
FoH2A3CvGSZCW0rvstRZmYtSwS8qbHR8zRfMsz+jDMnjrgSBpDrGPM2AnFJ6xrAxroLhJhzptXEw
tm0obX9kW5nBdLhYjUB3TY+fLougmrpFxbw9uxVEBEw8Iw3GqCi5kDsf6TsD+n0+QSkVX9dWVbd/
8974vBFmda80CGk/VC8W0VwvMyEvnAkPRYRwIxlWoV00WWXKnws4GHOQiTRLc7beJhgKUOw085uF
6AnCoKNqmiDLsMxEGxONZTWhA3DTTEgcKfmwPUWd5lP1RnG7Q6R54pqFPm1IiUDvjjHnfI4RyMMB
9VpxpMmt4coOgTQ5CBHpHookBmMPyzP4NYLJDD5SJ0t0jifmXgdRETtrczmLJx1+5n8GCLu17Nb8
F2QKtTws18DWmyPpeo98rxVF6CIqkYIblcwTBKPb7KTIxbqmI3u/M31Yy5vRjFDGMPYnzZsgdcFv
wwWFRrxiYjObiVrGf/unjJFteuF5wFsYw4TTxZ6G5qJvUl71XvD84Qg+vQjS7dfstT7ezwb9xawX
9b1AjuwGA1OYbwmfo98FMT9CcjySasgZjEB0R++B7z/uHSwufH9aKEwvJVdU/QA0yvx6URyQ4Wnk
84UttHFxN4rgbbA+MvPlY9ub6qAshqTucun7vlzj3pf4VkFMnCU8IGmcy6XAjTriMgmt0Qg0GwzK
hneonlBLuc3s9wXRx17XsuN8wFRsab+Xwa7k5xNifJs0dLUfBtD0q1sGuTBxnwTWXYcIUgdo442S
wqY5TLjqEDTesIvgEiT43TPNoGPNq9E5l9R+N4sBZuXro6Q+3eqIxvsmKMCvE/LwiwpvIJBlBEKA
nhpf/TZCBjlcChwe1oA1ritb6GHgmxo9LzJ7OBanxAauGzz4MgzaKsKhhyIqsIZX0J6iQCwlMOi8
JDMvekXgpf0WwOgdB61nDx8KtqFValyx0JiXC1ZiSQIPC9yt6FQrQzKrpUTNnHyl6cBmUX9uOKxd
t7t2TEGyb6rK1LRhPdFdt1jjDIr2i5WWsF6JqeJFmn8+RGac9Xkl7dxZlcuANfV/yjLAdRZprOFP
+EJHt6zy2dS1MOE+CPUg/njerEMwFiC8YzFVsUT48K7ABKaZP+1bfZ8zV1tQ/0r8Y253ZOGVA6sn
3VlpIGft5ZP6X+68R9tmJe2yRyUbozQ5fj/r0QqJoljKvQJir9rVMRaRmR6Dq7ubE7y0jQR2ZH5Z
2jH1ElilQHLt7OQAnWcyspFASU85x35oC8f1Di/5i3PKEPb4gD4iKGEtCa6erwBFCInCs5JyBAln
UHRIu6Gi/NVs1J1AI31qJNS4HVXm1JlVNNCxPCMGXcKPwRI59r8cX57wIAhqCOAoVN3u1VcLXa/4
ElBUw+8tssjPgPanOBa7s40B6E828Dt1guMipHv5sw4EZw7sYbbauG7ud9L/b+hNWHmrgcJOnTav
l6sUzjK8/EBmeiLVijBNqET5Ikl3i8SCKiI19NqEEK2vXVle0N4ETdEW0RtkeD3JXikOiOOg6CWP
MgxnYFRpDNw/hQyZavARDe3SK1GjNBTZnnz+5HMNdO3sqEU7eyFGe2uosSy5lYuNXjs1pFXpd9f4
OVsECJepYzoSzCuyp+F7+oXLImH3y8aYhaJs5Rr0BqY8W8v+NqcyVEKXjb+Q6UncY3CXdGv5kaSZ
UpPeRt/6eg3kiQlYURMTAIb/YHUh3Q/QrXtUQSAy5KuEx5G4B1H3CsQLumrXSY3X8aaZfDABWaPY
BDDHQ1PZYwrFQCF1i8wtV4nSSlbP641XUFBTw0qE6+gbqZYCleSHgOFvktd0wdJzqXpmSc+jRHeN
ScFk6mJmnzqhrneFcn8ry2q7g9i5kmjK8Hrky3WTTOscFelZezLA0Tp+8dFtolaGDzP+aIbTmK/d
7FDibyFRQx61J0ckKci3HA8cNLnbyni5x04t7+IlI24S62Lywj4jaN5ATT1n108OzIaEVwS+B6R+
bU5lV/yHgsgIes3fDUsresAZ5Y4+jD6eFNBL4chagS3786dsVM8UDviVEHtbrmcQrADbLkuaHG1Q
YB8PLrn2iZaqapX/utbVVBXCXFvwqGR1C2hwZY2r5msFRdzlz2iTqoQWxlumiGXB7zpAa+vEfWLB
4b4SGvQz4Nv1UFG/YedK8A/lNkHcSIyuFcIlBITyclIitOCW19QCkH1NcocwI6txoPIT9x0rX1Wx
tvzDNxBpo7QnpMmgs47flN6dm7UeX96uM3fXgrnY2gEFUCXnRI5LAbcmn2/Qsna7hMOJ7B65A54a
Jn29DuVtexRlZA2UQJrNuus+kclCUml5Hq/jQ/O8x5SbCHukGolBIS+gl1dpa40ipJx8RDKFuykN
+97+Znx+RRFp6lhkhxpEBo6SBC6ARxBlcz23afDGIUXZWvVxV4dCn7fnWb+COerUZRcPXltYFGNj
PTsUXe3uUS7DpTTAdYUQG2Z1oMmhPhiLXukVP/WbXtVHJds6ycWwAe1etVYArzluW6LiT280qQSI
i54g09H++OEh1KmzPwSmkQHy/T8XIYdyiAlRltQeDRzO4UVnTpuRVJS/yRlhGH1CqZ4GGdt/kyuP
JWHlV4TMSH+0J70e4e6Cj/4zJt8NErkPEywarRdAVN4PaLZyOZ8vc0BpEmjAZkEvUupx6hOuJl4h
/MULY1J8K6CYfaWciePOlew736uCP1cfRSz3XlJIqaVR2sgnc3DVHbWLsRvHcYcklgRSWUPe4vCx
Y42FLKDXF8Vu1qAVRBfS3mKkqOCKvqPZTlUDsr6O6wcOkSYbeZAAEC87N31XqxWSFb1RoOFeBp/5
E+IU/nDTDTucvyKcySO++H4G2RcVe7SYc/juwGBIrNtNA68+l1ELxjSaf4c0jR3N0H3qS+UpUwQ2
iNa4r/Jlgqtnv83a1yAqMLPhuuWxfKpWgE6775mR1tlIvMLHSPiBuCe0DrevQfRk9+Tmm/+/Kay3
vM9geGC+WH5uSt5AkoLX0XCXz+dHEFq11x9uIEyT4HXP4pK397/S0nfeo78AQ0DJ9CuuLUpKc9IE
ZY89uH7U2GwgR7ojXzGpiT87EN7kXuxIHVVM+EAZgz909jO4dSgHjHLCpxEY7eqrAfHTdF7ZxgYT
tR98lwIJqrROQXFseceUOzb14k4i7U2/b8/JJ6LFhoRw6kJM5aDthR/1fYn7R+Ki2gfYLWyUta0r
ST3vC4bNErzmD9x3bNr2HttJ7uWb/Tm8+prbtH7UMf0w2UUsGzwMaOmp7olC6D4J6M6AVJgOmQEl
AZ2BywOenp751UXlJIQSqRbqj2KfPCk6GfasZsOTSjxmGnkEmTL+8p0Nz39fPUgW+j5zotXiJ1gc
rOzSm5Z4MGL8vkFFQUIx2wIt2bF6uj73WHT4n2DiXBXWYGMK6xMu2hCj2woVEPzpqNi5wuPY6y2Q
Kt2GhcU2U/rpuasTfmBWiEu2Ya7v/AR11WOizBh1qRlDRd9i0E05fTGagmkXqrh4rgXyaI0rrCtF
Y4dLaj019IdQ8dMGvyY0rhSro1VQgDnvZu6TEhVQPilimqRSG2MogDIB34qFM6YZJovHepLJmqis
XZo4I3PxvvJqTSOhOenXXXSsw1N28/u+fcFMhXHlwHv0ELpiGDkbWMmQacqIHiUD+LOh5qw0mRJs
3VoXNwBtNCzpJpR2CuDllmea4aycKn/r1usez4v1G5xx3RUC4jTjnlh3unWwASYb0bZiEX9JG+XF
F0kZa6/LRy0Ub5iwRmy2QkgCPD/4M5F/NhkhKM6fyqeHmpHtdN8chBwAJ2kIRZ8bN4zJSJbr6bc1
eUSL1wpEyCufSAY0Mx33V4czrQm7cSVVDaOrppCmgzIIKYgK6tk9N0LrcIhRT5g5AzUBu4eb/Eou
C2X2dBTNdwr7KOdW7Ud3CEh5OARu7/sBcPOlq3ZBTzoiqiXId9yszojuf9tfoQ0fLMhFCu+bHDbd
yR7jm/MCG7A75oJsweGUy7LokCI0jkQlWhjmkA2YbiHKnFaAQBVs32wOlE6sqrGPAOpv5nAAbOh9
3Q3x3WhTjf5Mf/8FXLC2Zipmf8zxI2YMESUFHgTFyT8/WoOfHENrOsbb26XFvL/tW+JuTIu95AFR
z9DIaUaiClnonmJv2rjPa3XBvluOd7Fom1Tl+l02p+zPpvHYKD5CgqB+T0tJhQYN1WYeR8jQ3Z3w
6DrceXd2TUJG7RhugBdmYlZQFoUJ9YYzNnNr0M3fgVkS8OELSpVhH6AphvvM8+s1HIn5HJ2OH/70
rpLizn9XFbZMhpX92CVBFLW6zTjHG3zNfl45V9ek/hXYA5PmUMmvK2dgA+B0G+IbTJtdaMjvS3Hc
YgcyyPgi8dRh67qMc3waxX0768Le37XVSljKab2za7NPh+VdOBCJvZBNZk4LvuVUdslUY/U+t2/F
DJdCnaszMUKf0eFSnX9pGGznsyN5n6YiUq++VuPrk0ZS9bJ4V5+JUHKr0JOSjtXJNV0nSb6M3ikc
Bm/MmOnjFWNzf4WCyYb3c6tTpgf9DzN6YxHfmNQ2rJjGaNbbECxjsQNAX4pu0ZYb1aR/3hg9I1FR
I6cihThpkla8BYr5H0Y0Tr0ZD9f5DqAVZeYdjEW72yVV0W/ypcCLsnMDriCcgg9bimFuQqzsjfQs
7J65QeywqYn/+qPDWqEQVsA7p4uUWE9Epsz4R/4Y+H9lV8zt2haJG+fY8x+cuCy7b6F69IHD4hbl
ES4fAfikNh+vQOyqekbulQ/liZC59PqpemObFKeZ8QszNJ9zVhZz0OihTb89+RUbB9zlstBNzQAM
x2hT5fzL7PN8roQjdJr+p6KhDTNnV4rc/jAAZVn+hJRiFC+yHbk7Bjc2FNYroIncBHvoGXcIob8X
EQcQwX5UTlYcr82rK2LrjG6FdnV+zI2Sgsj8GxTz1cVnhl1DsPJ4QhAKPb7pghUaK3HYJqwriyZV
z2qvb4aMUcOPs7OFm7IN1Vhd88i/yqnolrAd9K9EAfVBnpEcDqyw5dCole9TVymRVx9InfNBGkk1
Nx80P24TlB+b+QI/+IWGd+iyXhrxVnWIExpt8696t3jj9XkzR57sMGAokdfeFBjZabSt+TkMYgEM
USCNE5KuIR0C0pVA8uyaZsHiqbzoN9BQ6zdz4+WNun/mdorKNxrdLIQSnqNBVCxQVGu8Azov8+Eq
ohjfgRwAsz4H/j8n3AlbgmVx+H3PsO0ITJp+lKdwJ5DZMUXUT1B6mc6xlS9YqoK0mwUnjQlsGkEa
UhS0IBwTYxlu9ltTljpDCzI6NqLEPLzS6hVoMl/E7P3gg/Mc3QFbG7uhVF4UisEB+Q3VfiQS99zj
DEaNTw1p/4+zEb3d6O4JC7q7gBg7UP8Ue+5dxMZUs9UJTX1ZrhCE7FGU751jK5UQQue4/IYehQ5H
2hZtX/kKmXZ7NTNJlCMPLYiXXvqZqWnJM6N8eNlf/7TemlJ4yI16K4aWyirFtnXoDOxh0c4QnkPd
5z2pO7AOsAND8d5I1LpdQIsvATvqMQ8GvnT+paIRX6Vs7DqZhVEaIWCVner4O6H65mD6iSFpwNqQ
1jV0+wjQ7FhvDevyROoxt2gkFGemi+byTLwFvV4y6lgEym3C58uVrESmdfOUOefScBVjvSELyXCl
gCzWK38p4CUbgCgSntbe8VOYcNNPcUSaiGB/hAmxZQZ684U2bvJ2SGeY9o7X7ujlG8H4jgJSnWti
DcFg6wvkY5GYuBnnNr9WBWtOgZo8MmhtgvjXv9pBSbJa11RO3RVuiUBp0NNclkXYUpEAmDa3Uykg
xvE7PF1zz0Cv4641Al2sAeGSX5FuydAygDs3ex7rnnUm+UbwRW+NFs/QGYQMPTFSwaa1chzapPwr
MCyrhvnGJhLMeCYf+Nfqy+Vk+zj/nN8plxHVrFfTDploid0gTBlMu7VLHP/TEfHLO6Fpx+g/LpW4
xeycW158KEo19QZ9r0xR8vJcOlwcKNDTJVKSAmewK1bZHGkWu7xZA5F+zK2GNX1YV4E3uza9tnDB
94wEEV4NQk3u0R1Ab27xzS/vsF8kVDVzfLhQbB49unnK/Dl5VZSL7i9pR+eK1T9VBoaQXZ3chs/b
ZOSGNzsNoV3gP6cRpL+hrLScst8Y6HyCei/4gsLKixseRciYBQWQ+qave8Q5SELdIARQHevBqPyb
efXd/0PF3mv0kMdOTTIflsdWAUVfRnetj+WRjRGvPVSvdx9Olcei7Y2VQtGKDd4h0sh8HjV3HirB
I/JaqY+UtUZoW8ZKwTbHYj3d202iWTTCsCWo9yVzOVHWchw3ujf/3apAf8ZojRE08kiGvnwNp7B7
jC7x9ELFXvXMr7gRIYwn6yd9dPeUzJV7YkZMSjfp/EkBjfE60cyftUIB9uJZ64GOGzcFOidlfuoD
YVdc85inAj5Uz/E+3dEo+xX8KdlZ7MhVMs0qOt+piPpP8Rs79d/9fDmGzpvkxrwiulFrbQf/Kk+q
vfWUTEjBcpkJglmHJK+8iqcGv9mU5qrigo4NsQrafSI7XVIqU2/OCuUFcMsnCtjJUiL0gXkQKpAY
gHTLqnz7xzKe9Qjl0RtoKuM8aZ9UW70ISxGK0OPEWZPrRA1VGpVafR/SFpHBDdxIzWz/RAxvkFpA
drKlIN2wdPmNnkbcBiTuoov5Ty+FgeRTx33qOznXiQoovGdIM7fkJQ37y2gR+ZTZ5M/ZUlPyWaBx
o75+ZZpTR6iCalxr3377f6hludItigWsYwgg2Bqoc/32H0lNBVa3wN5UrtnMQNQ32N6vmLIGhsTo
8MHdxVpuTVEFDK7bEKBnq1JxCy2abHk/PxFQ3/RW//OFGxCleF62Y7wOxUxmoK5vLj+F4YM26VuS
d7vJBtCtna7YnzpxKsVKiTp4Obp6FOMfysk2VQeEoGn2PUIDslKwvVz5m2PHHJAC81Fuqvf8fE+Q
JmImc182lMJDBZ2aQO8iWtnUbXvjWmS8JmYawvna4wOry28Eg29epYVsvp/EY7VVovvtkfFoTGj/
EdH9sSa5bw4hUTpevOE/CLpUBEcbUiPkP4yoKD9BHEzBX8pyUwiFAaZ5Jqc+bpSfYzqaxKN9Ric/
i3oN1dBMtvkDfl6CrhqSO1Y0SvZXn6N0n84k0M0LsiNChUp7zib63g2byGxeAZqMXD1wdFbZEX8b
ADJoJySsfe5K389UdN7zWaTUMeH7HEK+klk+ydG2XQc96whFyM8Q3YqGEotp2uGlszNqBCp6nyVN
QXAGQNiv5miot+tKWZG+p/OY4dAAebtMbHvPamr61uigb5GeqSqlM3wwI3ezvDbf64gHZidDrqfE
FBLcQIuK0fwCUWNDokZqgLStJbPSKdxJVI3wesnxpNyAFkVYLiFS2L/7TAMXAMzNPz7kugpeMcQt
AepMr7E4FIAa9I+S54e4SYCQveQ0aWBrkJJHsYfrgO71RA5y0PA3EZL2Y06wMf0SjWyF8AfJnUEM
i2e4MSZ8cW9lqG92+z553mTTTkGM39CsSSstZ2XhJkefxNaxQ+URuWSvsQmEx46c9av9fS+9JhI9
2FcwzSPeEHsYaduPXYiK44kU3GaG2iLjVgjwVai6buHiulurzZV1UYGyrI6Qy0gt0eEJf0IemWlC
NAaq5sEZxf61FNWOaOpQ/XTrmGmobn3qfLVgN+wxSY5LX9weaiOtEU/7aaTeUZQXR7bAbcSYQ71n
fEJoH8bjV0jRtyoF6EiBucPF9y7DhlOEAVuJ1EcNLaSKL/IsgTbbrwQ+OmmjNNb5SbHmR0k8DQqi
Xl8MT1PlDaOaVItMC9Jcmv/fF7EbjQIiDyRG69lazNY0gNZaUKjBVlh7lpyQGFIVvMDbiqmckf20
sJnUFsAZk2YwrPZRmvN8wLrC9LTE1KnO8YgGy5okVD0JLBsN/prxVWW6WuCrDaDRRagwKeAS0l8x
AmqNcecqwwB49zz4ZW/VtszhkO8dT2mlrpL6pYBIKS42CPaLqeYJH6VVBzE5oAc4Kd8HjZqZUTkC
ZRSIbBzLBWqilWIhUej/eyYa2avtD9bWrUeltJiAQrpF5u8Ibg6RwZuxPsc65F8LSEk7AG1wNLhX
jWWbxas46g88FPfrYWGRcaYE5TKXxLLCV8GlrvVzlw4l8GzhBPTkUsoAnBapsItxVX6tPLNlMV/d
gHEDNhv9LDH6k8I8O+PId+PRuf0JiYOpsSebFmg0L5Or3a4q6VJR11rB4tHv6kUlK91Mkr7YhK7F
eWnct5Y0cCpK7P3Ft5YrDBlU9RDqMuSWFGnw+B7mIMSmVOaZMJNsWUr4Pdw1etLmnRoX+Qz+oWXz
y9dlmosoPC4vM24V3qIHxSeBGwcNOgtJJ+VWHgO9KxLP61s/65dYp3iMD/xMKWmqi19VjOmQTw38
Xgn6HTOaltyntgdjOY9/47w0mJ1lraCtAqa8bjmxHhCsSkmxiYuHmWofDgGAo/oj0PIPoztqstBL
cczaLI+tb+VAZVF0AVNphQSgU8EgOvme/lcsj1XjXgnOUnXdJOErEprCwFspXFYvwdD6bJAHuu+c
RUwtB2MCXKIbIQEl8kYG2va96dwr5wpmWCX1hKtj3eytC8Uekoua2CX9OVpuyVfzjq3O7dTeyabh
Q0YqhjC6Db8NE07uRnuMGTqDjJywLz34YNnUsz5ji6gHIKlzwm6G1YsGaYqcC+eJC6sjzVXVqHST
zlIAjFfJat07pHRE3gTZl1QPclRYLGfQ9Fq9BeSBcOlqN82BJG8qx8FyDHQDBJBRs3U1futryj2h
Sn8BAXCP8wYPgh/MQ55T53ppvVD5sXSwRTwDRG0CJ5aDw0zanONMj4RBvfleuzyFuxnaNqgwv8sR
IsHWkzd2FhqQ2lXfyKKhooS04pGykOMckl2r2y15DeMrBxZVLUNxIqDs6Gp9x/0eDdICw9Yy22af
7TWy49LOH9b5IOsb6+NBgITc02JtOQRyjN68YEy2Qd71u1oIJmk4VsDcUtoLljxmwK979HAjx/oU
U8/WYrFGd3mlSb95mTkoJcLirFGjQ/BZlTYsNrUSN5q5BFQHgrHBbdE8cWtOxPhSvEiSwkUrSv8Y
lGml3u2cgrwiH/F0x8AGz/HUuCIrsr3Ng1HrUXsERJxwB7aIwSSCV9y2Y+c1+FFJulYY7WNxbK0T
HKTDW7eru59RWnVGrxZMveHGl2MfGU9KyRYBnVtaPKf5pf+J/wX25c01GcFjzi8l4kYGgLy3PnHd
hwJ722+VpITAn87fpZvtf6GORYi9sjxTtk52/M807P0z8dC7G1muTYQJJB1y27sjhRe7fRWoY78h
dav7q3jGTM+92uqZT7qevYhma3OBnDLQGYpUAJ4TLrAUHzY0F1SLVNmsPcmI5Lcr37f5OM87ZzoT
OMk2sFecaTt8cxRdYGnJ//pjo1TjADpW37cpfTJgxhjJj5yZmRUpzVnca9+Rx78WNPdXGELuQoi0
qe8lntrTzheHl654S+3jp0Ld1WRCJedbPIRqX//LBHljfl5wOKWBS9jzZQQGPyjlYvpf7E1tlaTD
fbaIwdQ7koisYSkg9JyTfFVsy1qNldrNyvxboFYm513b/ayRI6/Q/ucwGp/8NR+KFtS+WJNYVjhL
HU2KW3730WLDuxPdymH9fY05Qx5pvEId3keSmPXjXYoy2gsI/uIUgD4KJ1AVYmQ0NeXW8SK83HeC
CCf5Q2CIACorR+N36/Is4Ba/ZHATvN7EME65EmCdbdkaohkSJknNVcDU/Dou4iE9QYUoX6e3l574
0YR+5gCIVw+51tzPfWHw+TUaNdkkPFevVNwWcmxexLcLU+tSRe+0D59I5EGuBL49WxCwZVIm6jhM
qF400UAEnIwIwoxq07xgyhzWNazA9yZkNEmp+ifVFXpZrL0rKSTV7i3qT4J5DHhj7PfffeLJNHg0
Yh+eE9waB3HVUNQbQ+WloKZ8rJgRFRFjjMviGGx0u/Y73uzS1lAMOWbjVsN0bcTVKbcEwfMye/1K
fTC+OuCB1w5qsaSIbpw8rFwN14UQAQ7C5h5n09/bhqkFMuRHMV60f6N5pR0axZSDi9AYHIEipRJa
UIv0fehRXMsoHsXaJlNMZotgmQMmvMcBbUg6dEISL1csvXGFXFZEznSCBSzdCbq/t9iXDP46ydGD
OM3s2ZQQwQ8K/HEnu+bPtXOgxojKKwbQ5fh7XjgcMhoc488iDcraSBxaJ6na/WKdGPtS7069JtEE
jBL+Wkwvs6J5NLoSQs+O5k1OX8jChfoIF3U9zi/WgfocMlJStA+fLnj5xxZdRkT/CKwtMpNIePoz
yRrGBhEvJ5+uq+J9mxJqwrW0M1AXNj7cIxPCYFDIAn3Ai7dzq1tJo+H6lZN+EpawO7tBtpaGaYMY
wFkW7R6wgJYJ9aOoGsTfR3FpXAGDn7EJ7w203TT+lTFx4W/qrTkxuG2xQ3MacdMEPzZLDgH8coRp
nnoRsTbhcnpdrchfzvMdMCU35xgjRkBNfZnpPobFQSBh0z/+auMHgJL96mBrVVKygW0ONWiXMKPm
TOO0n9FZ+NN5DgpvyM9oSEKpOUtGGw1SRHOzhYuL6182XeQy+VNg17sCgqOzpU/WzGUZISqiiJEQ
1sbnqFUPP5RC0TrqnKBEr5zefxTChR/D6JUcQiHAMaFpvP6i/xFHU2lJK3ErEmn8/zr6l3h4CIBw
0i1tUZL5SjBJ3M3yo1i01W0FjLKuHzwZcnZFMYQHyTgOYZZCakGfGjDoUCCLCojNDjucGUubJE96
nm1ojERlX4tR3HvlSzv/E/5gJExsIDqlVHxHkHFS7cPYJ8ehYX778hoc+qG682aTc884S5o/cn7d
IQlymNjK/XlaI8KLSyQVx4TvIb3/tLbjfC6rfFRqvU9p3xl4f7tSQ0Bsu0AzEj4rT0peyHz/iI7a
8ZlDdILapTJlQzEOMTyBSrac43OltdxyikRqs++9ihUMxHJjqwch8PkrIEH0RoqQJaLCJGPk3cCt
3twzwLJR0w0nnqPimxKVhkc9tLQRKuxxo1vCIc9Vvif09BDwRZAqxMti0XJX/9vi6fUrPZgs6Ywy
S+180hnXSXI8YnN7ewLk536fX+7PVDUmnM2bMG51MnRO3J5KJ355giAlpo7yNjxgOTR4jZ9mLixj
xhelACsI5jaeggG2a50+AMFjHisz6maEp0ddvjqwQvkW3Eaexon+JNeQiseQ1FlgB/cnmoIB8hoQ
Zh6B3rDmZuT6dKG69NE+A7PMDgQgxluvRlu4qNQ0hn5keucGo1BukZISZ8a5cIOxjApA2e+nKkfw
efyfyI+FGPRSGwc+oSUlYJgM3taxDKZwhRc7ryjoP07bcNV9vdBzOklZoOpdMdXk/2x8bwLkHaWT
V+wFTZJRlqXWCsMvH/06mujwdS99xUbZ7CXkfzfcb2pnICghC6xy895gg9l17lMzVcFn+R+/nvji
fEJqtb3pr+BjJwDI9bvjaVPB6K3IsremiG8zqlcgOtHiVMw7JKPnSDUSBMPl6u0zFk4CpkqucUvB
dZEqXYAMpMwoekbHXB1T3euSYfgdP2ln7zR3GpxmatfVuX5mTqbCBs7PCCr3Ap8ulj06xgmf2/B2
U2mKoopu15O+Ae3zqsek0Zbqd4OoEyjhPVRyfa9C35gu3r0qJoL75aUAuuw9IyLGl+JaLok1+KTz
I0BlL87jfgr59/iiISU0XXcV5C/hFX8Yld/Nko8eD2iPtscJwMLJneDekHaVobYNycb4fpU2l3xs
ycuaAAY+pPNJSQJcUWp4vivzq2YmHZBdbSeMzNYiCJY1WmK2khnqF+LIYqAlDSJNCPWiPESyy2Cj
LdU5R1TdoITRr90OnRHU/LbpP7cjPyo/2NmzrwqYsDo5H+u+kfbgE4Q/0DUdDqP2cOAwEExiI8Ac
H35Wk4qHKrHUCyxd5/owJiIK30/vaPaBezoEVUuRZ/PS0/MSo54PNsONpGCnvPrCiTOzndtvW778
bbu80SKoiCt72hDClE4rNkANAeHcwFQ4dRGS039cGh22kDTzqeGBcGYwi9cuvJcS9gTHrOHAfMEW
wAh/puupFmPCvVSQS/bGW78OZNf2nzrerQvDMwXoqddBiB7LqysGLAlouYg/VkETvsc0wjxGap1n
ynqD8kQIMweHo4f5DMos7dCTpfpXRAWaF2kL2OCcO3lMPqvw98aBaf9uNcG87RWy25S+oqa3ldEJ
MnAxPjof1VVAp1kEzY1NGIJV5t7apil2tGFwTy/bQ/Wsn4wxMYpqsx22XlZbmZcC0oHlxWezwY8A
81l2ro6RI8povSeXNSNnCkirSuxBvfOKogggyeXrSr0JL5jHeeL2sEx8VbTltvqfKwWkzIxRrf1d
ljYz0zDxlztp61a/uWOfB1vMky1cpkWmJFNvG1/cYIj93kZ7PMYutbDVJkLbhNXrVPCpcD1p41xe
6TUnQKsZ88d/FgVP0f9YyUslQl9NmHYd4DEOCdVEBtjVgd7bt2uDqagJjOXBr12k5nkgxQY97M8b
7ic1QKXLRpe7I+BucAjkgD0Ew/3gS0SDNjDa48eZ+wPsY3kORN86Qfuy9SSKEki+iDBez2UXOrDD
kYiCrzlsZwTZ5IiYx80ATgih5svlhaQgE5obNi5+kJA7j4MieIAtt5OLXyyOW5Dzx0Q6B6wn5pEr
3vuzZEA3eNvrKqYULl1Nj6WUDLmu6FN/z8blGCjQWtgNQajIFkADHQWwOmNYbOaL7LE/fBPyNlr3
xG6wqT8D4GGFmofgV5Yw1cX8qBoQcU8JJDdpJPZhC/FkmdP+tAZUI2sSmoDJ02Fng9y0eBVtothw
6jRKS5KPxbnNpMeoyNn3jC5fr1W83ywEmviE+G7GmUQVo5/nwG2ypaaUifSGaEpW7DJ+1Xj/b29d
V2do8CIVN0jPsZCUabXOMG7qx3NbEIG7O8f7yXAL9+DZ5hLClQNyhROZaQ3Xfe4sn83bj3IziF8W
EPwVDQMoD1z41Gq4wsB+jshgAGkyG3EgJrOGe2J23b7waMo9gLHtv+hjghmv+cPptfWTyt5YlkkJ
L978anx7kovAnxrSEAhRr2zy7af+0HP9ZYlMfqvaL00XKV+QPqPlS74EGpEKkfCSiK76TiCrbiYN
3iiCfgHtfMgPdOeYMUVH9od42st0ZK+6+C6F8E0ndnCTLS+xfiVNGg33SM1Na4MOQXJH8u7DHbzb
m/Y6nBHt6pL0/2ykK5Orf2qUjHc+mBWaskh/AQYF3UthrikzGt0XxQUaLcEsfPXzSpqXSbprwa/e
ymccY/vPSsriDy/4cbxZ2NvGYQS339JiJYgzmbQVM3AFP9IIcfwr9QvkdKzLFXmQS/Ze+DP8iiWV
ujv+8Bp5kU/cWnhBgsiDW87hlZGLgy5LKUgqZ28Zai6mfCdnFlKMu95Wze+Bxhnah5Do0KMOtkGV
x97cp98ClsosI+1krI4RZCkl74UDVhvUIY48d6r+THlS7ke/4k5kKCYYxbwYWpLL3nJhRtu5ee/1
wk/fhC0NAlb8kbvFpHkq57IYWWMKFQj2orXovAfD4FrUx3GTkMobOdo4zD6IXydYxRHzNlGQVDLl
cd/JISDYM/gT2zvq1G5YZa/9fVqHfz1lIElLlKR67ywLbDDmZPE+6f59KM+tmSzrJNciy5428G3M
2MNbNPkRDrZHburm85iWYLfbpIQt69uy4p/A8yoS2rjOYAv+puDZQqgqIVeg4swJjD+JB7XkYJ6q
BIbnenom7sZ4ID/e0r48WPbMK8TF5T/OfwCbPOWEEUAX8VqeWNa+GuSTMxAM3NkhEGSy2xa8yQGW
TFmkTM+pERAy4yThOP4ymdN3i9leuL5cPsS/f7EF0SCDM6Tl65UoCO62DyFwR/VGP10mdienAtEY
X56u6oAMDAVxnWN9u9KZn1yOs1r4vm/C5wPjqEPt/+mLu8I4qi1+iHC1c/JKAoCRUHQQxTHa2oX1
aQBGEQEezq28qjcxTiR8Nk4nR1xaCBaMbxX7Q3krFw1Xmn05Q9BjkHJGnPLMN5qJar4fycqC5607
/9DtNsrVBosvTpTfEtQiGIY3mpp/brrD0DFNU1ZjSxZy7gkvKzTvUqDLiouBylVQPWjq+U5batCr
Drg3nlchppScy3Tv149NeoaS6ZQFNZUFMPRHuwjcuDOOIEsbZ+xnH/qTGZEl7TqVb+jBRXbRncUJ
GyIfU5ukTH7reDtHMs585fRPjsKoHHCe5Nve3X6VKdgeCfqOg6BYeHkzBqUyX49WhEkjSWQD4acQ
al8g59Mr3xkK8Q/cFft6IGfH9dxbp6JJYlegeHupa3rgco3eLJi1D5jUQSWogLbb0uc1Ob9hbpzu
ZxO5x+izQV/dC/06Ema0RrD07XQ3sWwr4GEMUUgUQAUVuyzmPGkQbuPFvAK2VXYNab7CmrhyCo0i
P84X7s3tFIRdnrP8rCCENEwTiQ8CeYOyzhhUZXBixzqZUTlz0twsOZg4EK+7i21Pzzd8UXrEyESI
8wF7NTFT54Z0iTKBMp+IrpXxUGO4mH6yTVC5T5QT8lK4XWvCuFw2FfxjDukPozVEh4UzDNMxjNfQ
9IKU1VATltTDrH+VZAlKZL4bdutXQD/FwAkI0nd7iGjEYPMA6DLyCNFLNcLN9GEikx95cxmVHDbd
c6hWvYHyTVnVh/ojQ+j06yL9aN/13P+fWCaSAnSRyXeIK4ZCdNArLC/515Yrx/TorGCqwDkhKfqa
Bxv4mOa0hjayz7YvnTWYatxeDVuanv2PmLZjmAMs0SiLN/QNkUTYPCR8QxvjdsbOMu67HgYYfXbj
gliw7pc3/C8ki7XdHRvclCDQEW+DzhdtufW2wo2AVqcKiYE+l0Cp47nwGii8Vnf1gfuLmBfc8mNT
cxZR46RvPjWn4ZuuVdbJghLWQL7gvD8HfBzdxHBx29iQ3ieQSBQNjmKENf/ZSWDM3Fs9afjfUfHK
ZtdHyvnR5VE9GXf+yRqEbQDf5wjYLDu0yPvLdkZrqSYxQ7iiII4ozu1X2B/aV0tDrEd1bR9p9dht
a1c5IMe28uG0iGUKj3riDjUGWWhvPZkyLKHT5gSKe3jVvXcAHjhAFnHn6fxJEq1YJbB+ep/w+4tC
Qc4n/lSnXP3mFmzqCb4+v0kiGH9oS1DZpknebvuo+dcwX8FK5msIcq/qVmlMKaLffJYGwVDHOzct
A9+d080AmX41wU2aeKnie5Lp/u0QviQDM4Bz+iGhVOYaYHw0Rl3uLINFAvFyryVC9gVZrC5grGYv
KOacBkAE3EiaAgxpvxB5is/CzSfLgY09ycYDr6U08HjHsVoAk+UC0VrLC+dUImmZgJitEbXc14q7
tWOMKxQj1cfgzkvKnMwqHQWd+XXAZBH+q+PKgHFwwD0gpkz6HBPrv4/V+2ic3Ufd80zetO2wdbiI
IQWB4bEmREsbXX8ygzsstei03MK6W+lg4QLLoaTdLcYDkEve9PFbs9io9JEvY8pqzdnZrj/xLmog
rKS+Xiy1D42OfZbw/kIqHe4MDC3Hq/2A5AHM7+Ugoh4gUn0tPsfSUamLPW3ZP0oUbHFRvyALUj9c
1nAjUK4pQGaSrkxBpdeBnUoMPF7gT7ZrJC3/mqgiiEUtV5S4whL7Rw4E23PyUFb0vz331SEs0eVI
uwidVRxugh0zAbqS3bi+Bx/in8eFIRlskzpA2OqvrzbruD5nClpPQju1AP9dNW2fu7wqqGwAXLNg
QN9ehyuxwgK+4R0O2IoSJ3oIzaRQ0UNhr+InsZwrAOSNHmskNa/D9a8jfmpSsvr4+G0gUEHN5pFu
1EhW6b4UT8LtBuDTbl7Sh4ov+bCMRD8O+ZCzcRdyQG+6uKKlcqx7jvkFnEvjQLvTnaSetlJYD9Mq
bP2t6BWJAXfttbML1bWEk7M9UwhxunVIzQjfvBQBeHIP5NmQi6Df03AFTxlAAljTVnHRDs1PgR7e
9MN83LIBFLBBDgsZ32OvhrIdYhSTPO9r4vA/1DHTpFSwo8Rx1oabYKwF4d/r0ncNI4Lr+XA1LjOq
1J3bBcxP5pmAgvSqHA2H7D9XD+bFS++OmAvi5U0Y+7huPgcN98njKa3KibpSq5stdKA/7nPL36zh
CUDjlLKJlSN9lXAGEdZjBaS9uhlZ/xtvshspUsBwhYtvIAiDhNaA/qchvBwmQVnTaphkM9HDMMtk
lnPOISq18lmqCEH6rmPNbDN9zwSOn+tKhOkD0p4AInFiGlPCO91a94LDxp+k0BCigeEUueCF55dF
JsUNHQhDQAf4u9Glcae+l8FcvgR0Akrxcr71O/rIyxAxG4V+HTI8f7pKcM9g6gjracPko5f5L9Kh
5IOD8E7Cf5m/V0gB+JZWWsiaLsLSB/bqtrNu8lw29e0q8HUbDvoMkHhegaeAR+vhYFBmlWJtWMj0
4ws3WFzXDEZV5jEC/jN3twXS+ZFdX+s+nUAA9Hrf2u7MvsGog72rGz+IZJ+2GprWNtk43RzhXdmw
+bKdebMYgR/RFuyK7hHz1d2LLVfd6HoRq9lUN3IFVk1ojLmk4kD25iLX9uHFlYbOVeLZIPp6RftB
MnpUWKv8aWfp236ouI8HjxjHLlxy9li4zb9zvxtQXfE75cd2XyndsHgTMfIBCzDlN/Jr8N+QkEF6
qDHYqJmwssQ0LE/Pi023CElFbjB7j9vn1PszhKLLjgkRjXHly7l0+1HBa1kpUEcoO0U3BUL0D1/B
vL5XUXp6fcUgaeTHvFZFpbwjtUHSbOIzv9OABRBaD+92MNSg0RKMPK5CwBVIWil9957MULbyN1p9
/DknjnHPcPKLEHSowCitSQAsHDLXkjf95rxf76YdCsIE8/ufkjLhibzhNNRA9JTI9Y/tIfmJdvBx
RdvZBh1lsf6xmwmN+4Z9cI1ODdleWot/e92cSWaKL8Fs2J+p7LzAaeSQfikVCRVGJc4/HcHEiA4z
SfUeY2KRDMihV66DS7Uaf1RgKE99jji9oh84sPVyZxH2nt17fQ/vt/60qxrgSAevHPA2eqlU64cF
YHQAde2lZkUU0AfXutZXjWJN/53WlQYfhAUFOKB/o914xGaudM+n2b6CuaC2AG3aws0SPCiyLwi4
OQH34Kew40UrxMVCfA2PUqAGN1RJRYxdVRSZwpCS6rW7ONdQb7VPTPfccdp7YgZqRJXFw7YiEUE4
KLDbv46HwLNrymDNNuxR6WVw5caPfYHSVUHBs2t6An6X38n+m4XljQtpPZzKIH04mBuYJawGUBPz
aQ+t+4KL4crL/E9/6qj4uuGwQBXvhB3yYjzkV9uoblxsLaW2hPhmAmc0Valtp7xT+BFF95i8jnrG
jxt97qgveGZjtB12iVrNPqSGCmnypnIkniSnjgKGT1S2LQRLDKVdChwjxxsLsqGc6DHL+fmHqFXY
6GE5hoFcnz9GKwSNOwslfdE5NQVVWdp7ypLQCELLmg2RtNAGMfacyhWjx19H4AyoJxR6EHeJ7xOF
58tqYcNygk9rOrcz6iPtrEXX9ZFujDfWRNw0S3KfN+eM1K9sFOu4NcoebpiXHV1uMFqis0Fb9+hA
InR8hQZUNx0iwvzhbokPuFz/i1BhQ7qoXK/X+8B0xB9O1pHSExkpeztN4E7vC4lvho1DHJ5T1Tdv
USuXDyBkDvb3lj6oBDT45o0Q2wslXcHCa5mz3F2MtzDyz4aaJP3xTzViyqYAjDti3gCi2nfkQjKl
q88htIUfHfnsemem09BBgpB0MrxxPSnHGJMvEI/0KXQ9+Gar3/6z2l4othAzWfnCn2o8QSGehBiT
+IWJFO732Xm16fYsI2BycKb4zilz+SBZvCO70P4YKhV1idejLTU6vSO1QteTQwh7e17uft1OIl45
pJF1VDTbvYZaMEPz6OTVt7kIAtCT3FqFwP83LYY5h/ieLDN9yXlRb7AwrQq8IGO/kcMEvPWnWfAn
ZolZs3JOsWF/Xe3hUFKWv9cmGNa9067qGqCfspKUXie0JV9g1LU/TeZThMj77Ijd81OxHUl7M3gp
yqXyVaiZ3FODKTex9cCukvsLcshDHYQXTzjyNzcdRZ7aICgFv3/sY1XcQn94dCSuv6YSAgednDNq
Oi4PP9FlBXJLVdEWN+WVvWfYubWfHuP51Aiik8DLlCvfQwEB233VbaYoblXUhohKKe8oSP/eeC0k
05yeKsE3B6T/dvtVX1nXYmten0eBfG7SwczOatA+3vm0bg1H4WliKS1/TUJakkpYqJEKXZrlZghM
OfJ2D81aEKMsmy9hIxwBH2qwK7zceld4SO1/JBaQzKL5Bv67kcdpQWTNEiDamk+lF6VPZP6CUnZ9
5Rm4QgaKCdlA7qEnrvt4opdXXnS8NNu26zWjw7vbEJvDoJocwHrM0LxexFc3BuZFR+nW8tZtinyR
nm+SzlmagW/IYlbh6aTaf+NpUXv2AVWfA2mzjL4BN8PEAFVh1hjm2JvxJDFZ1hWRHnLTabQICdxI
JcIyMMJH8m+hBP3sBrpjrGzfjySX5p+gYHNaEu645Yi59KtHrKKNJbAN0wg/JSSA55+OyQ8UM3my
q6Q4qztgZFBJbtTRG7O+HF4AyMS8gk3b9rhr3SWcQZyApg++JemzAuv4FML9GLQycseHTABFewRB
MxLDHnYvchZQ4PtfRDTNiqT0OxQhvFY/9pHhQmAIBohI1BRAxWLH2GerK9Ijt5ggq+iuE845GNxU
4EZMSJaTaZahvCMZqITcIhZGPvRFJWw8XNQZGrr58SjIudPScwIdmMWcUx3CBMd4DNeWXwxt44vd
1jqT9T9dtYbzTDHVFqIseCEGGKsuwpEJnd4WH0AE6B4jEg/mPYz85dUimuQnxVLsF6kl5vgW1ouc
Dm/YVJWH+3dz+aB4GmCh5iRpl0XGjhh9NKzNapXE3AaqqAmy1o9YebCQahB+8OuvucCnoEjxHJU1
kRiyY943BAnFzsgpuOH19WoXehtzpVfwG33tcNm1YOIre/Bcn+2Ud673oe4o7wDXtBmK/xMfj5KF
il81NdUuIC31JGnuo31I8BcO/8VeGCB8BnKWtyLCsMgNLXRo+XZ5hsfL0iUIileOgEJPbg3LYxgb
m0IVf+el9tBU4HqCt3Qn4UFhBb710YG+JrsS25k2iSd2JqJ3Qv+yIUk9IHYl9+gEJ3ReTH6OwIeB
DJ7UjOTNo6zyeMsTUUy3Rpc7lOtgGTI/jcaNxtdCTKC1gbxfmXDWpbAAuIpGNZxzrq5a+8UsOvuo
G7W8cO9y/JBHFzHQ2Z1hsjrABsGTs5ltAlOgs4SdUkdslrd18smaZKt75LY0bn4+N4caDhZV5xHz
734lCQW3Q5PvYrldSG1DO3cEUQ8J5E4soxNSfI3FWYnO+oE94/QGDcEBvGDJMKaqFP3V3IiwDH1k
2rL0zpysNI2SnxXmQpSod34dsR7BtnxFyxaFAmddRHlBHkHLozGTw5htFXKtdbGUXNnDAYeSBwKz
Y1UP5IgEm6zhwtp9lmN4x88cV05p48D5swqw/YzzxygJombX26UYB3PxpV/wjj/9/l4sO0gnzrUA
Cj2dRD+zvX1mXHYZKYdxYsbEc90zdLeODTventK452JnVgL8b22aEmMXSLB85STLnxIJNP/Brs7d
dq4AttkBn0JFPBNwOjMD8ybNwbcP6ZlUrHl984iViokwphKl8bdOUUTRnGIoMCJKM2qWAHRWcPLL
OcufifXHozTQNPfTod8FNsr49EBbohB7kRgEmP9Br96g37hoKy85BZePEKJJw8LUGdWSz+V5iAAH
m4s3NmtlOpizzw2nuzY3z6pFrFqQx4Ayh3p0RpF26kOdVfmQtXgvBkiSeC80ENmNF2x3tfQ1gYJk
Nq5XeJ5KseepEG3lvbUggppTBXKLYUW6c08CQQ9HKMgdHiwI+NuX+rM3FXU0niYZjPl5aLwvnzAk
NIJOCMXyzFEs0ksR8c9P2Iesfx5DTMzW1nCFWcJZWH9vH4MrcFZkA1ODFPnQUz4fBUPw7uRO5cqQ
ApHMQlMEf4crE6E/GrI514lsLC07o4v3T/TNLFyeJ+5+2HTlHquUzdTIvB5PeshjMYuX3Gft2bSL
jV7ciTqO/qG/R1DU7KsZjW52XS9RCmCqkM6ougFwgLet/lu3K5gJUUVOS2kUAc8Qb6r+Uf6XAgW/
IE/L9+HDCG0lhEeFPjfLy7WX5JNkUIwL5ukVeXEizUkBD6TWh+kDYrQFeEu4+fdu17JvWDXXL4ql
czV5PWlWWISYaKQQGVAgomZM9e9TdIcmpzwuMbt2yCbWpM2W9/gv/uPglklRR6HPA6ndfpEm0wmz
/63EfyADi4ocD0kCpnHPeMoRPNRDP/SnR/HbZAyM+r+HOCGnh0/FwuhzNW0PzrHm5Dhqk12UMJkm
RNkd13KphFWsWhqwSuB5ITvXdfC1DSc2+8SjMU17lYSWaE7oD+XHT1n6WkosOT6fftbapRGm38WY
H0NV5FAr36o1J9Dw7OafZg4ePp6JKudybF+Yd5QuII/p7TbqfKe6kzjKXfE95iZkRhVEAOswTfQY
AfJfoFOEfbMzogyg5cNEigXd8Itg5/ShcO5JTEs14leM72eju0W0OYhfY9iSJiDR/QWQpxdZofGM
Qfr1ca2y/GJu7dAAUpvUyGAN4L73SQNltLaBR9ZvX2Km9PqRNOCI6pyGZqwq+eevnxORYvPDi8hf
aTN5FVTaqPxYhCzz7cbvHzwwAM0xwbMj7QMZg4osAZzakHODKnf5RA3sYWsE3ksgsJTamgD5w72I
wylyvWBz1yhrpqh2O89xdD2L98WocMddcgoE3Gl81AdMjHKFSX6bEWXt3BtyI9YGSs6daaY/ZSsn
chp8C827eQC8TlSqJjiAS3vLYsL8pDk8PC56HK0fVNJV8v9AzoUeJ3GAmptxLM80zqmQ6gjd/FXy
NI5BdB8Qap2C5kxtnAu62m7Kr/A/T7263EKDeFdR8nF8xVudH5GgllKA5K9YpgaSrCl6PCZwVqfK
4q4PgX8XfChPBwXEBBEET79fOUUnthPD6T4wsLL9QjqXdgPQJDAw7ynOsIeOLoGvGVZ4rZ1aMQih
g/gK1OFN9Fnz3gkwBqakWiGkkYT9kaAhjNtnepTICnzjCv/vUoSE5Qa6o4vZndLrsGTIqfogcDi/
FWFDSeajHgZ4HvPZsNtX7clYJRgB+kbLbiF95gGN4ndAf8QvJHLNU4jBm+rONyYICK5IEV2baRU3
IZtPQ/IdodW78nP/Es/6B4pipd6/J8u4NAOKUt3UxhAWkU/V+LJzZtvGDkpMDL0ul+UGuEWXQ0Ry
0OVZi9ycA1ebvw7TYv7Csk4Re1cI6S6zIWD2KIKz4rHdS/XNoOIUt01Mt0uLu7dldNoSYjBXbsRs
A5+UybUFxiNtNWdpMcz36DnenCuBhhU0xfztZz+1TZEm+Z21qu6ngJLuQ9beKShT1S1BIr/VkwFt
zQ+lQPkfJxpC28XI9Ho5CvdjmKVNnGjktES8cB4hZutkVsqLOcIrPE6XAjlxwYt1ggO9E+SwgDK+
Z83pWbNh/WzB6+Q/kjG6xptOjSb6IYrfZfHn9R4sHCbyzAO2EXV5RFRy8HBFIGJ7sSO7pLelaML/
F8i4OyB8UTuV1vxr9ITzgR0W9E16iMxoF1xgOVMPkHJ1QsvwyA6nr50jb8/EJqo0RUDXwYbRI0Gv
OVDlZqsKEpOh8QrGu0bUjIF8yKG9eZoqE4M9KEK3jeHT4LkqvnMor0VHAiWDh534hDZ9g13U1eI4
XZvB8bChAypMb3A2JvwtcPDYU/POw1JOfiCM6Q78foF8q0wO9DSPUiuIx+qMu46wy+YU1luq0uR9
VQf1WZ2czdCgMD5dmlK/gtrU1tmPNY2ruEHda31iMw37rAPeaxKoNwpWJfWH/4H83pjaBG9eKaGz
Lnab/63qMzIgFnqXBX0EuOmTKb3q1YQY0I4zMB/yUR1NW9pOR1FSJ8VeA25Tvl2sud/ZJpqlO79v
sUm2yvtn+NiKQ/6gJHe9vvOu6+HpBiR4VNeMVK9z0UJ36SKAuMH7UHml3mGy3Uyvb7qc9/MK4H2T
WkC3n3JJkOTFibLO8/r/sERcHzj4OVBXpj5YqRgzVMyX8szVmvTwiI3FF1OjkxW7P5BXGSOZMweP
E0lHgnItFbpBdF7V/om/DCTyWtKRqGx6grc6qxtZgNbVzaTzsCXRcTIJRU2yCl5SWQTtrsjGB+8U
fpNb8H2UUosaw+KOOkPdbcqO6nKdlo3Mt+3UUd05vCxEjoAHlXnx3325S0vzhOl53gT1CqRjTXZv
EGgFoqDHDLHMx08hWvaudhXfcnbsTOXSRuTQTdP+HYRc68SDPACQrEny7rmsG+AqY+tvLjxRrL+c
rhdkazM+z8MZxWpaP+Ynvp/dPxQp9dUzRlKVEVwDgw9XfIsgxCMqGAPlde9+XQgwu8/LNW4xKrKL
fl9/GNk41ATz7jx14JUCi7908rt6QAKyR4sll0J7KqkSyl7rcYS1bpxwQShddtHYxR582HSygX4a
rHoKz1S8D9qsSBik9NHV3di3vxv2iJ4ZRR7yxeyTxrqYOdPGTQECmL5F1fcdU9yIDLm5bpApNEXJ
vQzA8R6Fg0AmOXtjUrl2Ja8gfV7kDC2XqjPxc30sM6PxRtMqn/5g//8BYIyovb5bJyo+8Sgur3MB
FhU4jPqDxGqYpB3SWbtSe2DxKey5XYT7pQ7p3291yu5LL452yOk1G/OhroZvUMPbBjL8BJFME7g8
d2l2dl1uvYLPjXxWJJtKBSjaLMTul9lWvP1VYoxbLqfTPCp8oOI888h0PnSvdem8k2gNHrXusSZR
1ACrlnFxbsgj7kCLZ1rRvWtpkEr8xTpXUzvSQFtbVv34ITyHQAlC08ugL1GBk+V3LZTL4FZd0g9O
SomHLotzgw4w4tpSVGXMzSrWFko1iDxSle7Q2uraZeP4lTv2kEiyiIwqiNeIGluHjeBIy9cgil6N
+pACbRgiutuueQiiaY/UoUVPY3lnyEf/JdT8QFDx+seEmkB080zh+acANgFNWqqLiIKeV+eUw4MN
xeajPHe9NrLxmhdzvlEXFTApyoKj/dNdu+hTEJTZjniKKhS6YWWXI87A0Pw22hswba6/ldvGi+uA
QA3yoBIHl8HTgT6M04jYWKUyy9I8FmktmMeiQGp/2/JC8ms2zIZLxBX0TGzJJf9bec0V5Ndq4KIi
A3e99yjcVqH6UX8XkMBSpHPvHmiNgbS/M7zCCY2/MRJ11cNYkvTyaV0O5JPQPF+xbzmYiSr7ybBy
P0H2IXfbk641S9cWC//SeIAh6oTPOEbEiHmSU82exej5CuHGmo/49f1Qc7N3OAQ1bPRTS/73OODh
NmGY0nfNEwGCm0KZP8nA+kzx3R2uUHMKdbcjHtbtogse8pAEgdrOvoJQOZcMZ8PYFxKXK3AMRjvW
AeiWQ4hYrj3VSMsuuLprYdb3xp2jOFqY+nD3lauNGWU2zTm5gsHjBrydI5YuBytLjYM++AVne8KD
Fhd0n0eKA7zhtx9zqBfd5aSdVVN3rEjhgqB/icgIdSur306shYQimIJ/eYwMzcRb+phoJP2DE9/B
jaI11mnMYgoW+nRwiE238beU4wokaP77j+8cW0xOGxdLdGiuZKpHpeiEtvx1JZg6Nkl6aNlxVxm4
Cf8veWMmvDNhHUUKIXPE9nONSpXEjkHWJJxOUWuO3DswTNwtHvJMEa+owgRDQa9uIsIykNVcaKG+
fYP2K5+3lM6jVqBDC5hIey+6Sbm3He9PyMLtIg6rG5OkdkCHBC0jhdNS+mX0oAJQYzdxWKJqARvs
uPWgRpme0/v8UO6SRpTz7AmpyaBVbXwyiCNaKb0EsWNpcZhIde/kpoj64SCg2Pn9P/q/cSXRJLSY
Pw4/BIfjJXCOD4gWw5+NkkrtdPAUfg2Iv73/Mmm5JpJKgrIWdpBIVA79bjKrRraodzgv6mMbnnoy
vcSeGVdIfgmy/pkGZRPkRxOd56d6P7+STYRWFrgAVJwTEdyLE6ORHA9JWqVg1jHFgehRG9d7PUsK
6AnoNBtObX11E8GueiAJLBWA7mJcVqUGSwJIVDKb3jMcKK4dICY4CBnYvpLU59iYRqGlGHPx55/X
rgNwvY4X+s7QALPNI9cEhLfoty5PMDE7m2gGdW9Iv4EP/tz6ZDnFYMX5XHFnUAPmW/d/5C68l0re
wCt+yrpPrklYlIp6sINLhMmxMkrlncKiWiNxIVhn6HlgIVpEX640eLTR6M2C4sijClqZ/nUcPySL
7KJ5dF5aB+VkXIi2kM1zakh1mV6Z4L43rYdwAw1PD7Ohb7A2gSRg0deD+Awh5w8viDgwN7sCCwqn
ZZQQzJoojUlJiMTSAioMACMFPlZQ6Zru69cyp11TmKY22v4LnckL61W4pTJrh9uP7HUbHqMGaieC
zwy9TmyJTgJQh2F+n3rNXPdGitArnFiTPPQ9JTyOuAj74/aYIf8iKBLxQHGlweD+rlhaeLIB4js9
1Cp3xZ0CvMddUQNCMn5+nZEjynwUOdmwofSZbsfDenllhLueJTXHwqRJRTU/E4wAPYK5dHKpOIPj
65ltAVnNeEW70pcohlE5aiHPv5U2CBvRvHOz3SLBV1QLmEvaut3JlXMZgGVBO+c26ToqV//jzhgu
GKT5bys1cjb5XXYfqZfMvxO6G0B/8hI2h6uVQOdz5e/TH7WPdrmWTs2VoRUTY5ZK12Vi4OH3jvWK
bJzFC50QP45BGvNsZ+hrUfOJ574JBVX6JhQ6NkJzA7JST5fqA5bIJ6hLt55XnVtCT8nd6LKSqgnp
cJ7RB58VYQ/jyEjB3VLtZxLJQu2MmFvEleXe9iZLCpqTg41Ww3Hno9/FIHCaPZCq1atTWezxXGaj
0fFJ/xVqJnz7CDC0uzVBEgij6ox8C0qLXWmeTBpkAFZOBFRp50fdJnyfz1UHiUgQL64FLKlHSIG7
KQ3tse1bzRfTX3KQ+vaLYZVLl1xRB3mAnbtCsGQHIR3G0efNg8PTVbPYj82nPTVvLqT1wtSvlDcY
0bFQLyzHIr5MbPQrVdW8fT7NzkB3PoPIpRS+lTFEmJgQNavDaZHqgTbhHqO6S+Y/8N0NX63Y3IL+
5ng9NVxegFafuVqjNrTOQz2Yjz7+BXxbESH12fp5fjO22pVd8Tl/sxn5P4BV1zPhpMqKxDSMQAII
oP505G0hj/+g+iy5w5J27L+C2qdzlXO1L8ltyRWcPp4NA/1cfhSpmACXH8aiQrlHQWgf8p0eVBf1
5dG6x9hb0Q4WfIMPeKt82CCId3gfve85LQTzg9P7sqprARVayb4+BZxs6nGyiO/03xXIhHNyTcuh
71tv7324KQekGvtYpnSSM+4ctJVtqnGOpWr2ItnNVkMAMPIO6yqt8apOEdIvzpZOCagUDtKxx/qI
NhIO8n7eOGRLoVvZ6XJAGePQJXKqi3WsFxsnYgnpnMLL45GXXdqauYmysh1mg+sqewQ2iFo4ZSOu
/5Tez+5Dk4ShyuPHnDm9QqSf1P9KaPRujsxok+BZ2R9IwNDVp7TixEi3d8aVqgk5AsYc3w9P232y
iE48nIMpHrXOoe6RnoC9dDxLLvWfhj+VukUEsiXVP0q5ulxthiGneIK3edh7W+igRhHg7zvhbVHF
4lNy13z4G0RrLMwlVPcxJ92OS72BuyFo+Tct5L1q0v8JqgW42j1NP5W7oGTk+wOiwkKgiv+QqAmP
xnv67egngD4KLIF/aDge/ZI4IpzXw6ZRIKAuUg7q8Y1KTJSB4APcYA/OyURb/8frggmqERpDTwU7
/5GH/qPAZ7OXTM7pAbki7uRaP2lgC+pDPu7CxX9eDOUsh0pTwi+9AG9VlvrZl4ozCdn/QfRBz9ao
bWCzgpS0pYg0kaysaXMXgoroXi59YK0ngSgkqc0OlRybrOEWNIYJhshaaPu1BxZsHprlvehXXj/m
HSjBcabN1KaWE3FePZSkUU4hk2FZzhVQ2ab8nH+5xF8xRZi3CTmgXyVyRr55fcCaucpdnxJvid0J
zFzeO9BepIUf2p/6FAu9RvpY7MY3YUS5aD7lOotHv3qRzzMJ5FC7Kq2Pk/I8TcJeslB6h8m4aq74
TH2H7L6A2g9UnWpcRmnC9lMuwPOvBEAnMxDaYBfSor+u6fG9ZAEokjEcr2Zsa4gsZeRFMHshvK/+
Q5vLpoWMIpEMNiZVZCCc3pQLM/8sR5q4Mztw8XGJnO+cmJlI3GuPW6sK7Je2ZfyTKq9BxrgZfV1B
+Xd1imflGReOoODyjT1HcRs+58RII88cH99LlU0tARtBbYiaVtpjIk3SmcGS37FWQkICnH3F9gr1
Fc4Boma5uWOUlXQK8/GCUIXizH132SYG5gplbLQ/vAxXVE1KbqLGV5H3r5zWGUfHG/Oiq2F12Zce
PO3+X1rTALwoAVRMMg5ASafFnJIasc3aIBdwPXQiGVES8mxLUoO3I11YsZ4zCZ9qx2ZtiY0nbgjL
mmL3YRcKzaETClUpm19g5PbHwGbOHUFElUiyM2DrufxzxykLrZk1yp1S8rbMy42H1LT50lbEIBDF
vjOurBWFmb92ANA1qOYNLWxSKrxDt+wxk9LLn3gbLLA1vHbsmU0IKARGG+XKhEN9kYSrVQ6Yas0i
HzE91GDOwQlfXKyh+VyaiUj7KYABGR+ByYgrg8ms4ucI0qWSjzQv+RCjFoNkm4PSXni6dqSXvhJg
DCKDIfrToBH+/ROwFThTeC16/ZZi43R9aa1yWVlq2e6GhKEUDu9uTebP52TfyCXZTOK7vcZuaDSZ
kiYd06eILux0Iwd5NU8qyDM5D/pj6yVdVm1kQNWsV6k1aFc4OpjbMZl3TpWyyxK+wkq5m41EGxBU
b2qjzta7osHYGt7NE5FT6Amf859riDMW9UT3Nn0NdKC68vogm1d/A29N1qUncZjGHY7Rvu0mk5W6
mR+7e3PLr1ySOwmkQKZJrz1A8+MoVGIIGPeRbQS3tFnDM4HUbuMK+q5cctEwmsxhKjyI/IZLTl23
5Lsdec+0mBJ8qaaaQ2coUKVnko6DJkni0m38rD9bGpaNfBb9szcxbkn0XxPEd3zDqfgpWgpi16eH
SkNludOsX65JNxSVtBD82pF/Tqziate0BUcllUozmGvvOMU92GH8fX3NzqJtJi6xqKSvTCChe0Sq
1cw3xJ0De1E6y/jLTm2z/u9K+zFfK8Q6NCQQw4+DdzZ8t1EaqnBQbmURfKQuyrDgJ6tjCtTp2RH9
j5dRkqYa39vE6m76dKiSy4jDO8SHMKi6DFAuvIHvWO/PBgr/qC4K3vVLEZZhxDxj+qczFYuPQYfS
pCLaZVTPfTiRYBorTSMV3m+0yyORRTR2yQeZjLY0egzFJFYPuIHyeM6vP70GzGZPRzO9c1saYwCS
o7bJamv+IjX9c9IsHV4+0wgH+YBn5Du02HknKwmjfXaCJ6wtYwdPRnlW3CCC15+XRbnAp1iIPL/O
qgrTMFz4xHRGM3lTw20BJ9kCyQ6ha48gB5vKwrwXhoEzSjNgygm9R+LUPHGSEcCXAomCfZn7sOzS
+ozu1kINZUmGsRpWNZJAPjXAjSsQAR3sA0ZUM9tX8fHUBCpEpRCwIVshdCsfxYBYbysXscQ0wAkk
FBvpKMprA9s0DK6FMCUPxsiO7Zc3+AbQaqnPDLVucBbYFriFnNsSM6ov+6idSZmXMqw/cgBe2/mH
aaKl4g319XjUAkRCHVrgvsDVNzvbDVwg0uWpGjiHGyPZnFXE89in4UZS3AQnEcQdPiJg3MOjpRdQ
IxLWiFBTEV0Hu6T8LX403URcSpsF+AsbJsQY5ui6GU/JoI40rhK/RPNzkQR5DqYwGn7vmNTOlnTr
HSfcvICHCReRFI5GYlyU6/A3G7bd5lQ7oaR+LzwCv8ljEjsWQrITZIccBji7OFCQxq8Ec8iJDnVt
jnteKL7vu7lifFc+8eS2SGbqN7viL5GHa72UP26YLVIJFbnQmh/os4iFrYesvXazkMrEZBDjLXdc
KWNSWSkVUVEpG3QonhvIqZajN82n2lH4OmU7gA5jLzGoX8cb7FGkZt6feuZodveDtzy4+SRgGc/a
R2yf2cQ23U/kPpCVlo0/pbJPQQi6Be1jR83fg3J81Nve5iuhQuReXwFDIxXEogxvXeqxZI62Gpie
LyVLw7ou4qPtOAqINR53o80kZjJN5TJB1x0h+JAgCXXaIR2L669GQQ4DMFSiTnv/FrVxkgP7wn9i
hR3sQeNHM788f/H5KBqRmEcYewCk8VeUIFl1/mZE/2F+Q3WPeMBmnP/FKtusJSQKKR4p7Gf/4wDc
wxdd56ZuIz9VeJx0eHchazoiCpEz4NNrtH1oqgxt0o24xHbkeLsG5io1JtmOokzWGhfJy4D5Sc9+
u19HjOjgE+xP8KzQYaAvVgdtnJTQiAq2iN2jR9MXAChaOOFE0n96V4QrCf4/I0mgT/btWKISToyB
Lrz+1gpusBw6gYc+md5oyr2/hrD5Ub9y+JFqdPD9vMoLMJqVdpJSUWPESYrygLkR/N9w3mzB+SEA
jBc9CpmWKBfdvhimFV8una6vrICRTt32lAedT+A+4jMLvlXfllsrO9FGH0nEbplYAcL6tHbU2Hbl
N1ir8PdpktdI5KEMeYkOYkTBus/J6sX5wtSDhg/PFMN4gNEaz52cMz24De/cvPW97PSCDSTO0wLf
UEp8A1zmRpjhAiI5zcGvutmRCj5ty4tyrLcugop01wZfnvWW8MDEBXWWc0bRy076hPYms3Dwq4IG
Mlitui7rVoyGdZTENo0atll76s0DZ6FXlaFXkgKv3aaFuE2rtWo4afXA33p6KagjIyL0UTf3bR8t
uIbvXF7NtPQho4wAC3SXoxUxzhCCdDrJ3sjUnhrVKORQtj11sfBOJkQYmsbQ11xdjP1X385v1LtU
Lz/kPkQDGGbJr2NEp2fFcw/YwI+NxTXuO6wu0pXYXC1ZSVKDPkR0yR1yv9iS8k211k7ROxuLz40v
0YagI3az4Bxj2Ro1ZPDFdiLmGxoF8qpEhW+BgH4+h3csBNCUlMj4rt9aA1KubWl6DfRddNzL4UpB
wnKXOKIyAQDSAnPZsDYiG2zKOOp2X4vaFdUPE6Cf383AxSpuPlN9RsWz8cTEWtzlUI1fjmlOqXT3
uP0600HJMg/mmN3HrPcsdc0Mvh1yxqwr8s4/09Jy2Y1OXwe4BH1NHgElw/BJ85HDwfe2+7FFDGPD
dQTfAs+spbR40CACecmKOhDAMCc0BNBPhkScZr0yhLIG4BzqmnUtDQ2RR3PHqq2Y7D6mcanUAVMx
EWtXcEbKy3ChhW3d17JmGDzi0WV9vw2hzgBwDLQd0xwgldJ8vod4a97XTke9+IEm+lsZmQmawHPI
20j7ABwAvU7wMEFT1PDTJ4oRK2/kgAET7zMwqHBDefz4V1biacwNh2ykMhHtgIXMp7hu74nASH5f
bKYrBk9jpp/KdM2hu/5xOJI2+TrwQsXhUj3zfYVqc60J6BHTLIMlLDbA9SKFTE/HXRGWF3f7Zorl
UWg8egZGyPrC6eU4qIkJeQPU34RFG/MmHc9E6tSiE1othDMgIIduFd1QJ1zAk7OD5Yi4bS/2hhz+
rBwb3x4FvrqQIsV8k5iQFaBMUZyWOh7J4zz2CoRDIOxO2hKsgtlxeECc/HyZrQ5E1yKAGfews+Te
Uztr423kk65Va723r42QLoC/kl4ZnjLnu6UsoyaUpp/xtB69TMzz5ee6lapoQpqJD6uWVo9xj9ac
YVp51DDz1U+EZzqm/5q4q8vpO2juyAPsJfZ5KY3LNMChq1wRquGA3BauDWtY3fwB0bg6B1i24YrV
+0eZ4rlBZdGCD7tyneOgYrRABPv/e16shCGTqiSu7UbBWS3+uuL9uoaOfKqLjxxJaAfJMUMXoRbJ
f7avMi8lAjciS+N5AbrbrG3w8NjYyWHYFerA8GmwQjOBgkHmIqQN4o6LL8gFZ6nzR4W8nmeDJEFs
ZVYEu0vg/0kMDacVwT3j3NNnQcP62iLKNskotve4H5lo8GmNkzkvrXYu+1fn62ezYBJBrDALifQN
nly19fODHeI5SWcX7nCz1pzV5lppL7rSw4OtMmLKNPEEX27h9JQDNnQoPKZA60OWX5Tqiu5gUzvw
c6Yv0ozgopvL7xHt8ng7VjR2tEOWEmo9dV5oVKJPyzKAEnvHYvgDYa7cM9WpJOP1NMSquMraI4R/
HVc4Jn8mE5Yq22rnofDKh6ZiDwXnp+65xj4QX3r4bZpdfYEHl55U/oz3805SEKxlwUVyzXrEqiQc
ZblwXfGqYMsRYdrSBH9mYDzaPvmIU4Buw0LcAmE7q9CtJL9irwrnHdYuA/QIekt9hc0bZvHxRvBj
bvmdFUxoCqwAv3i7ZRWcf3SGhJHHlh2L9elxjeK1Y+imSa8dd0ItY3OJHX1SchK8ckf2lYMYZWYT
2MQdIXBvYtIUhQV37ND4KcF7DHi6IjBJ42YuhFT4R88EGqoZ9XZ+WR8ZRrzuCzlugHU1H8MYbWeu
tLd9vpu0F1mz0ESGcsqvK39aPzK6cWXAqi6WMUyd+5rT//6zkneiDAN+5yHCzPlOHl0t5b89DJq7
OnhW6fliWz6qlqxkbeHzTBvD6LaN4cmyyTSCXgIE6YvThDT0kJ30NqWGJslJ8JWEzNVKrSiC4ydk
Tg7cfTnPOV+A2SrLh9lLvXjYGTFnogN91Xu5gG1N9jOxf7sxmA1ll62qF4jdCzSfrK2zNs0+gnm3
byvg0ryn1W6Imkw3EbHXMvtHzRdtjcm41OhPM6F9u6bycQlWdg7Bg+nb7bR3BYG2bnONTeNmt0qv
L8nX4Dct/pGrlqCYrECGpCZCLOQowyY5f8ensdrvCp5qc21Ly0pZwbDw96RmFRbug8YdvD2QKnij
3gvbUiwH0nJmJw/zi+WnBArCXMInAEiJkhddsI80jc4h705RqEoraunB0ffjmFc70MIERjdII7w8
pgS3zcGiQC8vmE3rVnvAXO/nlSk2MWRYJ9nXzg1W9qhNEKmF3+Ppe4o79FdQi8er23EziTbWC8Su
X7OJtb0w1CrZSVnA8l18XdD+gMVMQwBuEKPUs9motIfd6fTS3NiLxi6PUzcMutY37TE8YojOddgn
W5/0TrnGKp0leKk7COd0nw/mG71oiIRm3hXOV04ONzZ4kCrsbX/+Wj3bdBEXgvFC5TT2fuQ/eDH8
fgsM2vx0NMPHUWLjIg4Mb3/9bIsdMUoJ1utAvm6rMlHaxbrc9/OdcH9HnHGklom//p44976iOSA1
k1slA08lcVlrVqqaqZzPQon80HsM9MoK8Dios0C+ma29Qv6pDQQz62ZuVES7o79NC7+OKOr2z2bD
rKol0Oq/6h7UNpvtJ9lFdp/Yxg/l6t5geM6X4ibkqq9oVOguMjd8/UjX+3QYQj0+uMpFEg2oC/bP
ZXAuZsUIu/MBPgUM9tIhzD3/7yQP35OZzrNrOa50A10DQRsxbaB9s0EQUUgNBnUQR1Yfr/ZewRK/
d0xW2Rhx5tC00AkUnXXeQ8NxX94vT5kAbKZsUNVJryk/cQgH60nqxC30TZ3pTe7h/KgsnM/1jC8g
pMoNWH8INz6JyXVXSJGjKS4hoG1gRZbLDjk8FEDvR3OI8+oM5Z4Hre7q1mk8cKWdNyK1MiS/46v5
+311tfMeIMiUG5wFTiIZAAf/Hk4hp//3z5gdeSI9PUPHJnFElMkTdNhhEsopR7AbQvHf08y7gKe1
VgoEU66XbP3KKchrii6Y8E15+U+GD9SRV//f2M3iuxAFxN9z7DgJI3d1y2/HCtpcKbCci8RaXCJP
WHZnJZDpoof6oYNWL2TIVcwf/nELE9VxpQiF13Qubiyh34i8W+nP5/xHTpFTY1RzFAdW/Le4p9Cw
R1/GoQOnQ5fX9GG0uQ9d1RaQq4ajhvelCwkKDE5+DRVxlPdWVLnUUy+pER5S2O2tqnyIpnZsy+xf
fo6Kb3oMY4OIMdX0THc/jhIzGnB7NL2Rj8TOB8AIxHlBfq+3CCwPPCmlMgUVZx5/mBRPEVqqeaQA
9f1TrfdEZBbFwRXsnL60dmlA/lVOvVg5mzAZpa5JPAohQEV46lbz4rMZtXvZWPavWA4hZLmfVWlP
bFZyyrx/AWfjVXOEgwU+7PKvFaduF4lfPNJqaNu2PiKKLzdVrjHiXun3UIwr7Qtq+76XRczoI3X/
kB+l2+H5uGubB/5Q+NScF6I/J3MVMenCsVlpzqdxyNpSHrd0cfZ8tqtK0Xgu6gz8akFiq7wQEgoj
Bjv7087EQ1V4eIzQo604FV9vynWUUH3EJs4Afrd+WfLct075shCLy9irPkecnwX/vMqEHMW7IUMc
P/isA3/anBB0vNyAiy16U2z29ZDL4hGrS/gL1QHXiO76mfQsqsBSGDWYLbMGFt3CoGz2HbMag9XA
uVxBh3iXsKFVRsoF3DOy318QlxKjRUzrXakO+cdRoXWPVif7xA3czpNdiRnNQwXxqSdTsQQk/VtW
VNrMFeL4TItSBoKphtd3fy71aETCtrrv3WXajPbzuRRucLXDgEzd+Q8YLU0ZqvADHaesDIm5afC0
o3i9XTrDd5fjRFOYSqKCMO5ND6JV+Lj5gh+IqY1JxckpJ2knC3N96Zm3ulV7zgNmpP805/9pyNGZ
NvjPyRvRNQR6P3Epcr9ankAM13vFz93ZjVQ+v9KBgY+HmMBy+CFZidd/Nzuc9RlOTxrpTIj9mHZ4
pW4DkZDBX9L7HlVMxrxGhaHwnMUBCRLcGsB3AcxHUTDT3a07KeO3pmLNiTqKVaoTO5oUHWUvQnuD
usy4Uj7tQGIP2dGFM4uNoIbG9OaHNq9OtIAK4JYcRBXIh12bsRZ+XVvU/Sk9t/jUTedwcmcnAV0I
0AzGrsB1SDfO+AwjuMiDFEdWaPy9V+gTDEnNw+EXLjyhibY/Wf+leBtr8Wvanjm9wHA+Aptz6czf
dyNPZPuXP11ivexSN2ykVxC/tTaiTCEqxD3LDmEDh0m2D5T5EmsZNMcjZY5iE0NY1v0tWUNYNsLo
sEF7Xzx7rZhoS5pFBh36vswMCk8FNXa06DonM3jQsKKv6uuWs5Wrb1fsBFsjM6MucqHXnp1vVcPs
DM/4xX1I4mCriaXdL+U7eqb4g/cr7VDTDIRX0RuUqvbkVb4fVYtqRFvq2KOX8+rq59kzFNq0i7L9
7RIPL3IsebJWTX0Zb61q5rjb3D9O4LjkI38bnquipJErBLDbDJh/zhK+HOs/zXJVGC3kCKzdEAT6
jzYjqkCIV/LM4ehlhlpeOjIFINLuchCCdlS/edb/4JWWthwjhoT0QOoA/xIuQ1TUB/3gbvogJyO2
kzSa1nI8jbtBRXE2ZTrUkn9J6YMF/aZCRDhPiv8z1/imeVyAHmCH5js689IfjsIuE8wwdgIXVtRi
lNjDhEXTHQW4me8St2wNPaOrsGw7R9USgr9e5UuCm5zeILUiFwyoLMw6/QqPzDUUGqmOw66gn7mb
OYzVFG0Jxu1TIOzwhoMSB52OSjaS29Myqu0uHdGF6FpHo2pI9qImazrmCSvyMYIIFys8nIVvNwEx
l+U4QABI/eeaD9pkU6NSgus5LdGhy5qzjsBQsb3rh6FQHBrmqM2Tmly+rORUw3OVwGWhXmJOqlKI
VLyn8jdHUFUQ1+hsKabaygEJ6uQLC5jlYiVdRUBvuge0LHit93t6ZyeocNhiKHvOMy8IDVYxsAko
EcRcqH2WXxOLE3Rf2z0MKw1TvQVq4swbjfYLpEmgs9/HFEAUu+7CgXwnpI4R1DtAqpePzReiVGuI
fqpqClwwm3q2ak+tVLD/q/5B5i5+mVj9GwoHPv7VbVfT6+3NlKv4vAFRm/roV8Ef3L+U0S1zLOfZ
OqNYj/XNVwREZsC+C35dAarQ43kEsoLqpSID3pqhFXLzwKEzsN3zPhT9R6RCruzIj9qsG+sRUK3q
G2RBwTHpWM6IUhe9woTvE4veqCsOfy0oEfFQhHyKrZL583GLbNcbPAH9YAvk1C6D+NA5/ASYOaIl
1CDQk0LMKZCchSdH3g0zGP5+rEapL9HaHPTyUTItPXjCa9Eeb3+jnhbNerO5vKfjxZfea13stPkt
kAySHTLsDVjRg+YOVzO64y9Qt0Bcv8T6KdaiOXTLbvaE6OxP93WzlUTLKxv+HKTbVJuWFC6Mk9wq
J7GtvkYsSDOV7szy8Nh7/OP8I799gM7fZ0Qx48I7ppyOc07smE/Y6kbWf4wryyN9t3AyvWzxu1iy
ujdrVgZczVFbP+saF8vbq1jIPnq9Lbovt6oBi0fFNA3bUwpeEGJHuM/vcDCxK6iPD0VGYWVif2V1
oQArSWvBgf1gOvLB+qCROc75jOKtJH2w/4YyOP1SDc4NYV4X132hDUt19WJGQlguvisN2HECkPHR
aGlPjIYTR0HVocLrGG5c6zlSKqBzdk7DPnUNpIKieKBEuAAzrvLkXvnxHPeDPy6pZf/+jPLFMzn9
siFdVyrr1EOXoi1bl4agqyshXRBUC5GNfJ02n1b+atQe9ntp3rb1UVwWYyrDKAO4gXNoDHhHLp9J
N+n28vEcD05YWNFwxEGdUGvo5v/KdftkPdCg3ZPrkIHrdgqeShd982kw7MqjHWEC35r9TRx4d5Qk
pD+NWg3O4J9nqNiot7LorGVcYKgnNppEExcCCBy+n/2Z+7SVK3OmgqlhR2o34boj0NqxkOMnSPsI
xg5lqt5NaFCk9vylfI8WICJ7mxRIwfzTig72qh/yjiVYLG2R3gyw8ZvFJp9BDuPkUj3Mnec9gEVC
0txT1oMTrvYghEnS6OmzTAUXsAciGPN35MoD6vG2W82hzii2TziuUusm1eKFIieeGo1cHxZTpr42
8w5DO8CgsNDjw3o/3OP3gI5DGtkyCw6kcDO/YvtoQQ85bGWKUU8trYO+gB/mQnzNvIpgBLJdLTX6
or3bCgNl2bkBb2cAOl4S+K3mvCxjm4NUS8SxgUZIG2MqOhDvn2uqfinE96ZB5x5QZWLV8NjWFOGX
tYQe1gpn29nFjn71gCPlrggnGX/kAKz03OBe6q/zBRDIYWSkceWtQXAkdkMqbNndkeSGXlUxNX+7
IdS+jyAQ4GU32lTAFkfKc0yfU8sC2N7daNRb7CzXtvEjKQknlGGM1J4RC6UbJK2eJksJ2RvEY0JY
XpxS1YconZ9jZwBHOeEdHyVx/yJyfiqGAKf+sy2+FVDej5+CWeSvFDcTcoF9c4gMMm1tA+HE4Qm5
snG+rEEoE4Qa0XJ+k3GQKHOLaRVGbznTZyCBoiv7obZfeDZOuN/lTWBR1w/bG22KvF63Yxlmv2jP
OB0+4Oxk0IGbdDpR2dvZ6hEb1vi5mz+tfN2J+HlWEZMx65M1dPMmCSezk4PDEa5yuJPTvgk6k9ki
glw/pd3L9UatgTTL+WsO4bCrDwJSAIm8wxMPr5/x1GG1+xh04/hXli8jVlX9T2TKvwXG6qGQXZIL
7gB31G2t+iI6nj+aBL4vh9SJ4DAkL8sWr2z1BNN+1MnecJutpYTC0auInp7Doo4pnKPl0WQYfWJ9
LC+Da69hGxPdKR3d9M4dj3ZqGXa9m7llQ2oHkpgxV/ONAXto13RL8NJ4vd8s/27gUR/YxhdEsUcT
+GPpW4PHKlcp80O8udpyUbx2pfNelrWj3oQJo9cJl6LvEWPxlEnmV3z5fUU1c6Cq15nhAzT3hp2T
KFvDBs19XQ2qTy2oA9kNhXGZ6BwI97j7XqKGLM4ovo3KdtZj+2J2TWNbuhv5Itb9V9fS1hEp4akA
sM7UfBML+rHpC0UMTOHUqseS9XYkK+CFRvnZtWyMykbh0wEa+6SryX15HYX21IjX8mVwYvIY3VRQ
YbOV1I+xGp0mUpg2WKZmwadpD7Os6vTSQxMtkLgXoasWOJxVfUd7jcPof970YtR/t37YxwCpkLo+
xXWMZQmK60rx1SVthjAlpJyDOjYq9kRHDnpc3Czb4XaM2TnxqfEosw6z39qNwavCV7Va3NXDXy+h
8H+o+WM4rXxrHxMg/eNwQ3Jkft5ByURn89ok5Zn6K4Jfp7AVTdXi4ixcGPjaqeXd5sUog58vutjd
RoGdnqPhk6LDgRS48TDjSW53IX7El0barxsSZPaiVihQUIPekXU3gZBFy8KEEAkdbDpJoNzsCbc/
RAv5Osqi5dqzIbcQK+4D0WRDTYpM5kudnbMnc+kQHHwBUoBeUc6ptW7U0hpKeDQeX5SLsz8R+DUs
ckZOQLOK04ThhvOCfCEJFWhImJdZi+BjEfVAjEuZRgYNT2AFdmT6q2C9bA02M9eACW8jNQxDuWKh
oJu88MW2I+uJkn0DMjAj5ELYvN6sIxEQbctZGR3GqAAUQwyQtOEIQyR60rApHK+fpaFpG/MzV125
y1Gtkv87XtUF7yeqtXPkQovr42Xqa/c0QIxHLLPvdEY0lGqUBONNvpKAGQ28gaEZc0QzSSRjDE64
6OY2n9c4om3VIDwxdFSIl3lDwKCi4xXc3RLP+cXz9dhO1DfULdlOUvNzaI8B2gxKAOxuLSjNhU60
Dhg+9v6EC/JWugQAJzgESCsHorb1i+BkK9saFqBg63ST/KKjvAKe+H1gjZoDCyBpeX+YfBIP9PuD
EgGjzMLhOyi+OyK92spCM14hNANt/MZzYvknCHAWDrJRFKD9YVfzyBEryXzYoG7/HIv6g/0ZhioW
d+eU+vLNhBOylc1rqSf0wt/RBieAMlsmxoQJWX8pzbnb/BMI5r6tgJlzzMHhA19SZFFYUg/JJKwf
EypxEJbhOubhbmBScYzadW/JCVI4BY+INYbH3rg1nUXjiyZqI5MCTJieOo1gO0+xqMz2Vj2W+aFj
wpG8mM2ZmPGPWBc/zEa8A1FtkclrqBeiM1GyAMvqumocgz4qKvRJ6vP15nLIRojaOI1sOLmeu/V9
CCAh/hJuVCNYq60sye7pd1S99C9hDka/i7nq8cAvqg8YHbLzrqDlxie9kVUtwRAn3jSN9hRXNt6l
+1h/u/PALDCyjGvuHaEgMQ2OkebNREwwteevlaO46XYtF/Z2gRS675EVJ7yhYmKvZx5WHhrqHvtZ
oOjkDv120iBdX1+n0aksP6Ro+NjH3x+SMSH/5a+QXqi4adeajrRJVoRBMylSQ9G3SxFp9oGVVKvw
vahFQcIe2APgv0rxGBY6PznFFXpMZl2zDfJMMMn8sK+B1llyQ0QVT6QTud8Z8kkoC363MYm7Uipx
s0tucBpf7duasvYnx1uBdEn7CTSseDoVsTOCnC5F5Q8XP5kxr6Lh9/ZA4j2KQFuHcyzh/61rIStE
4/m0voZoaiS+0GeiSsIlyKQBDVG/+CBLLcw9GkMTAed1WQym6Ia9FnoIL7cpg1qO0XTwBYlj6xxH
jBXMyGq0aIJqCaoRlcC/9ix2+0bMGQRyBg7FthGvYz4YlJpFCV7vplb7acHLJPnj3ktiS2LxFwtg
EE3moxyYBao/D8cYp7IhbpVnPH9lI0t0wWuIxbtVbeTZE1xMv+HfEw6iJYXGlJYWFeSkQ6b77ok/
tHUr5l5vG9oef6SGqK4s0vs56UNaYgOWXHtZWgZbi6KPPrMJDpi4y2HriNoYAl97U6XsH54GAGD2
xrzVQlKkyis1E/5GVbc6ndv+VuZmVetlvPDxD9HUled6m6c6PIVyeTpoDPzuK+AbveJCF05vf6/O
NrKEtrtGJUeHk97JcQ54d54r0XZgIffqHXZ4/Kcy7V/3Vz339S9ojK90I1EwThqwypeeBuB2njQx
eqBztcE57/XxN9CL+5/EA/Nf12/8p+pMESu2RT+AgfnCRrq2Ue1g6Z2vCLU1IMxk6bbmMviTycA3
vTq9u5nnOdoq+L83RXmb3PpDNfPnRAfpjT2lD9DVtgxvJ+7wFg/gs+u9kzoexdscUgnX2a6jYexz
g/nrtl2upJf3qs+9CWh3ZuCwXdMBCXgHFTMKCv2tgscmQR0gi4frnyfwXptzevfkGbiW0CNFl9oN
Ad0IBMRLZy7+0nbtQ7h//zURM9f5Edb2y0PpXvf7oE99w73ELMkjmorBq5UNQcSHjhuAVGzHX02G
DQ7ERkrFpEHe7tXaFGoki95iOg/UaJr4FbkVHLF3QFGZfAOZtPVuIfGqKjwKaPtmdg100HVpA/mD
/+ux9cLva+zVgE2/HKISzvQgRvgLCsQJJ2ttDIQ/L2zEnyFiA7LRmJskGAwrJcR8lFE2dfyVSn9N
JFHXDlSbaHu08Rg5ZAUrvOtKM141+4kYQVzYhQZHd1quCBT6YOJahyARzQP5Mm+pj3UQGnHn+i4d
qy7GDwkQrw+Xkmz4sF0EbFCwyqrkOWnNVNxWCFAZGhbY8WCyOGoy5vc2u6Wh+lXrsipBM3332E9i
Rq6WCyCogqbuk6nWdqpEvQpVF/WWwwWOTdabFrM9PYmrqEYmAyMTEv/Vac4Q7y6+xDTLuHl4awMD
ZIMvbfn1iP/y9Gyvho0sWeKO2qtZkp8VfO+D7OAJatYwtLWeEyISO4tYh9hNiP4eCjOE1ksKYEYU
XXJYescVeM5fiEXhtrM2PLUmHWHw9mpbEFXczaITAlDrArUxD+n+yGgaPqYANTycdbSh2K6/Ajey
lGid5O+vQbKSLj3j0FQaDMMhvmAAL1W3A7dxJoOD6g4ox0mMjvbNFeA/V0lIvrHgvyxq5pBiMpz3
oL5k9Ab3XV9wghze0+Oe1YZe+WBnIedkUKyR8njzRs7YDv+btryCdItTNbVEzSi3XMXk342cikwG
snY25bWmIiYthnXzPzXZ541H3Y9P9dDrDZgwya/StTWLwPL+ogpIoxQUnfUqd6WAxfQaoSKdH14k
zskku0vHG/YxE3ckSfz/MVFq3EjywpcQCntW7JFKGhAPA12SDm7BjjH2ZX5hoKFTdw0At4D9Aj2K
4bAYgXkBl9OipSVihhdRcdfgpYi6xbv48MPgd+5QaDgTVe9jMeJgX5cDxr8BVZCRff0AJ4AXc1O9
NnqhE32u6+pWYGX+/vU8ftWslnsPPZ/q2ifQk76pVYoDfzW5hVFP4XddlyAII8zdcowAlFI+JNCm
bsBY2PvA0WkO6doc5h9QxQZgX500/onlvRJugtvJedGQwgME1I9QgBVUa3d/0lGwdIfHwOscYLAL
vZ5LNLbRZocfNIjgOa+GMEvCHYr4U8+eWk7V89vwfZRly4crW4bMC6nTSwhnHn3jB/hEE9fmHKFu
Gr5jIQc7xR6S0IV4lBdLoXQxgeLOyg0iPttclaMVI0kUHIAMlXTsg3eilDr++nD5GWUf35iA0G6E
vLyXyltuMKjXjJnxI28dYYItP5dBOWEWsibLSqVfat8X72uOiXacb4w/YNVZHt7+G+Rz2LZGyx6n
R2A6njlIgGuDKldTX5S3Ce54+UDKbUxkwjHaJi7zynsWwA5RZ7GYVhqIxBLfhGJMf1lw4ZW5BGFn
MeYLtygALxuu7uzEVY1s6UdevlPNdiyTZI7/JsIeAz3IVPJqvHT9PUN0bfQffl0XYcdMVVw2Rmik
XQ+VSWa2w1WZnMk0M2OuCnEyLD75K3fIt/wrBdSAEqcKdJxDvNmy3fJjFWQvC6f4gQhK2YmA8yXi
kjGbMD0CLmpIAtIUof6hROpKfy63Vf/HwGNGUxZ98HTH7r9DoigdhY57xJHZI9EBMy2a2Ptl+/MO
hfnYk+uDJI6tKQkpeYkRz37ZH8V+iGMW4pVBtlr274ATEM75CG2i9rvlQRqwV99oVQa2ONG3mgRq
frBFNl56x6rVsbFTpo+rAI2BAYbZGPSPychWh0iXKOsuQJ+wCcRurdrLH2yvjfafiUusyZzXxdz+
pVZkzq4dQufXQihg94ZZHTaV7mfZr4NPhPzNJVodzI6kS6E5NEBly9o+ZStKZp79yNhH+K8z8Iz3
lZkSCGxzdKKw/beBIjQdcPYA2jUIkd/iwYPsxQm73O+74jiF8Ej0utrNIJlTp/+d3iGpHYqQ4Mso
wivy8sjVOtRCwQU1b3LvmItisZOprVnDduMwyi8dhwczj1zR2YuXarOSC2POsb8dKYKw45IycC+v
vLOBb54+PRgxzTbjXdH6YaHcJmqw1oYwTOIJdKgBaYjNdgjm6R2M/5klnI21lbyU24XW//0Kp7Ea
Wa9inWnMmly/DCCmaPikPgua9fxok8KsrkjZDYthcCH35le5uzRwpTLigCy1NOtA5i0VXvZoMp7G
j1NNIqD5btQVbk9692Bb5UdPdLIa8j2pdn8P2mxeWyN9p4gH+AHQAgKEUA90YFI52EXoQ+q7Mgcc
tMsQ8v/0/nWOjQe99g3X6OZvJImQKFyiPITqLc/rargmVVxFNjoCMJtc83PCwgdgw+GsKPJO6P1e
kHpKwC1tOR+KJqihhyeI8n8QAKekOD+1RawCBFdYIF+X+qH809FdMO8ueQLXLXmz70A3VIvwxuM7
UII2xHwz9h6LpzcAgAx7zvN81/EM2xnTFz3NslQ0/8o1elhujIxeK5Mbu1tqphY5z9XRIUohdAeN
Uv3jsKJhIQGC9hDCW8gowmk0Sy9x4/q0xJFcdr4l7/ZGlMHNhQIkgZXW4TrbB27gIdZUWZeeYVXp
RwR/WAhSS0KV+Tbu0ck2Lk4qf5+fYdUuwwBNRB5tk/XETaU9H1rOwwQp3GzVn0HCu0htiAo7LXri
HyH42Wkimgzz0CnsV4Q9dRjZb8u78FXcCIAILgzl1ZuxuQhPBjd5ivZKwZPYGuG75ASE8IH4WRR+
8r5/jdDsU8q8sbqr4EOG7ka6mHU47xDd7woxnIE69XrDxp7Hq3bhwF9Gw5ptRkiu+f8d89EF/1MH
Q6U+d1xn9l0o51UmClpxUM/aKNDOH5twgMYTMDCuhwY0giennH5dLyLDkYV+FTq84hL0/WZ2DP4m
/lJpeI7j0Y1+VUd5ktMF6tjBU/fpniJXaYZoUXn8VmVszZUSUxzdbWEMPEGuZlHeMNUSa1HyFdNs
kU5QbsFtgesjMQz8icB9yNtsJFTPvE3Oa+AYQ8jHzQRjZ9xn4V1fxpXIUMKtBVlo+7JLHSMohv0R
6KzV0ULLgwQM1Wa1oaQrzVxGanJg0XMnJ1lqnpU9hLngXX89wXrKLfmixT2y56eFcSiM93YsPqHg
J9vXk9vdsgoneu2Wnzy/1PKQFWcvehcwhpGqR/7D+AsxH2JTbHOQpDKosb2iRZQdOEnbW+hEJxcz
dnd3NyD4FQ5YjzFq9KVRt2Czi5xULqZRCGdanT4rmS5Q8vXoUkZY+YtPN3m8dRQD8wJSfBiTpP9i
Z3AOpJQN9vDGpTx3kiNRZBsYEjK1hFR3tAGMqDhj72kO7S2YNBd78ak04lVxru4wjd7ILWGUF6nP
iHubaYTSET4NEA7yAW2gRAAzys6o5PovF0+tSO4sQ+2Rf8C+O/SbAxhfawYvMS10lkm/QH+iAEJ8
5GwweZnxlPkEMVuDlwihM4wDCgEbyNAWTePLDz2t5VBVB3eYFb8doXuMr3ynJ661t1n1iTDh+sn5
BT7lRDNKj+zq4O9JIoW4ax6nKEkkTAGHxMQqQNETpACo2Hd7pxu3KJ9fHoABuhh3/yCd6NBGpGxB
CFJrn6XHuX12fPq/XiGBJIGMw+vYKp3rTbJxh/wVt2VgZljwEkQDhDzTekNoSXKa4XoyXHZBYGw4
XRSbfHjzHYKSPtE9g3Szg/UOtayPUQ3317rHn9YarNNVXwnq/wZ/CnHj7RGt3plCIk5cEyVbyoYA
Fj5rBsjgLvfT2dl9tcNiqoJH52NRHogfrq7kau+lEc4+UBx9KvGCJhjEzAsYkTPDx33FcZ18whU/
z3Ju1v5/3yxjy0DcT6K2n+Uno3cDo7ltkdN8iK8KBZGAx2VewvDDbPDumRWJbhgOw99FNTVCqlzn
x/R7C9J2fEYaga5CMsSc7PhntGT9JYUFB/IPnexfgPD5xq4xCPSCy/UZ4mfh5uqctseiUAFZO2Hj
P+XjEdpcyNLFIPuJE+t7/+aZSkmEDO/ZIHkP9AwsUwxAocslVVSi8WpStQxJ9lsAKNGE4kudkwMT
eDQD04LJqwp6RUxiPm+eOZrcKgsfmQGPftNXtOLmFDF8LCXVJDp7kMGMcIxYODfWjZ9nDzgk4T/5
wpNA62aNZL40vqf3OsgPgobMZdy9GtTZzWhUZWGeOov/XDEhrwHHZgEJs5MF+zsLh+hoJq7suycr
qCjsUEiiEE84kfwWzRGgRgvI5wpa1fTqujwfgLynvUqmBibZwEftnSt3pqTQL2WC7JJkndf7lCB8
TjbIjYvGlkqtE83U2hvYs6wWBVm4p3nr0T32UYE8rkvAJ76q/FrEITnI5NXd3lV3CsWZRTiNwXnP
oyaQgyrwLsVhWpnDChEY6aYLswZgnfD33CCO+fk+cd6g4pHk3gQO2CaWA0VXaypOxyNdh8I5ez2c
gBkQTvvgN/8Xbie2yBS7bJc1qIaUvkGfGee51e6GdRbsxfg10qn9Ee8yglIPYyPZIVivDuu3cF9e
hkqdezK5Oxxb9Z3B+s0Jsi2NepfDOULhrZjXIrfns4sOpdYvDuNXwuLFCg3tSV0u5mCyakKW6g+g
0Lqwz9mCMUWAeyHEQ8MpaCId/+9Ak9SQ7LueZEXZ+EAzYWcgh11isIeQ4t6FTHYGmi+RFQ2mB3eM
2zRfFHEeL2KUXEYIIOPLfrXTGrm/ahblDZXqQFhd+WX6Cb64RQBWJONVPAXQ42GtqtplBuWgEMIp
HDgl1pbzzchGjRrmXnK3W/PqllvgHb78kyZuFbjGWuiqJ8FXFnWobIyPwSFW+maE/z7Ncfv5amU+
Jgxh+O6M7xul5rwd5kLxrt0tmjgAz4E4tN/Aox4HRejQCF0NdEwJNL1F/qRnUrgBkmASZbd68TET
pO1wd3G1WoAibp9l0QNfC5HhES/4qz3q7ucoIl8FZVqRem6pnjEEXRxeVFTkXLjdqYhBH/yIF9kw
DZ0CigzVMx+nMrCCUlp4hY+htRztq0nDS5t4UV2A1XZkP8tKHV5G3Mb2L894E5QqCAiNI0rpQ1c0
HW1LcbJeR+gAJffMxJ1Bc4UWe7JvfGsHAhQL89hsml+mwP3f800MD1mW5dpM2o7RgIJLgcsMcUto
DXZPg1ZHPUbSzhx4f9eqG3K2mZmqfbmUsgN21u5CRbpbHTM5vkez7Ra2GAPny1T6oolORT3Cbk+a
eRAWetDR/eCMV81+5psmj2sLYfZzPP8FA2+ABk17WP/5D2QA0NZW0Fsn98/aE3PImM7HjXDdLjDe
ggHlN8cTt7HdA1yU7/DUp12h6sb0npEdJzx7f1DmJqGVl+l9qSXzkfzn8mNXaB4FR66wdGBg719Y
BuLbmEL4mDwyIq8/kvvTPiF7SA8GFoNvrIY4QC4jWs0T5fQ1w4IoZkz32+yzltfc/bcF+IWoSCra
Iv/68s5JKJ+/3nrJr0UI1NQ3AeptWhW95Jf1qAwr4ito546BiNAOXRnrP2Vk5gNGaWYUbaf6jGGH
BV5fa41nD1geK7VCnu1r8lkRTqux8yHNdpB4JBTLvx7T0CCMDSFOkXDPlSRdhV/3QiSIQmOAf+nq
xBu31DoGSdOsrLULP6K5GHIcyuBl0F/JJ4uyYKMlFJ++pUlD4orTw3b1LNgPo1czT709+LmqaNJW
hbD365Wwf9MsdQL+QiILOHfGU38l9uJX0QCdfpQJ46s8kK6X/LVJ+mZY9WvblNFe1S99i4RVnmwG
VRbMv5paMThU4PKFu0rs7qYmS3DiI086CDV/nz/HNGF0b6VdZ89yk7Jo7uLyB8Gqh5EmwtP/iawJ
bV/jxntPCPoOwQZfVaSzhr3aFfCWyvLN5hxhFaIdb9uVsDqDCCmhNPgw9zQrzJzA7gxEbJCNN5KU
oMUVAakbmCEaM2zvPp55l/ADw8dtxt7wsYyKmZIrJcwiddu4kqbanp5xWpHaqgpSoRNg5zbPhhPi
X2jkBfZjj1ddTQz2VV9JmrRV+ZOzh1FAI4MRKQxjNEL6YBJC/OrO61csm3VEpGRNaZtdn3l28vNU
3faP/C0qckD+062uAhsLo2Rm+E4pihvUndhlr6S21e69UOfWuWAuLThqCvHKonBBlrof4iDwq/3w
v+rP0/E3ETbRVKKXZ1Cg49++Mys4yEz+wnjGmTx3wlCnJ5wUh5xYMybFxNsyxG8hlDXLhoZcxqXa
aDCQiS55gWb1CTCBiRx75dAcg/WeEv10beSNSCkMdVJ/r3HZuMgO/TDMeoT+aFyyN8h3T2loEn1N
oHsPoxd5MyS2UL/l2fIEhD2RxWId2Rvn3YJa9K0ykQVMfkpigDgEVj3sEx9BEFnE6qrAJPKBw3ji
cInh9mIgBoIGxdmTfbisO3muhOqsaJRdNoQ1vf0jj7D5qyvIIxnrt1UcGRZk7d8PnOBtMzA63yEk
xT/95cXG7cQrR81DQ711+iK7e8QuqfleeMxlnfwgnknoH1rnfPd6npJmaAqi1slexAa+lu/xtFgj
N/2Ly70ZRS7HVlvEfco7WO9CfkF1fsUsCCq/9FCeJ9YgqP+v3ZJIhTfc05WBaWATjqL8roou6f1P
/+o4W/Crr3mUtQdQc0EuWyLMmLio5v7m3vKvvg3BU0JZk1GIP+uKa4a0223GvoShF7sP5Y/59pvN
EIC841yPibuOfmMzjxNB0oF4P2Skyg/Q7BGRM1Fy5L2YHzX5IWcZ2ezIFA7KBFav2Oq1T5K191d0
Ty/RR/rj1oL5Z24cQmN5HVgLWURYKrrPmLT6b6V/4sqUNtYQLSkPb9OpHYXxzcJ6x5aku7S8iJzj
QZskj26GK2Xa3EAQIKc4OiJJSuitct6Y/CY8yjzSQ3gG/jG2KsGRn0hfVJsMmcY+Oce2Gp/gbv5q
ctsqttS2R+M5BArTDCceB9oFHGSejT1IJePXyNnvhYCZIBxY5SgUtTjGN0cuUNmmlBCyUrav8Vt3
YMkjUPlC/ED3gIWWLy71Dpe4v5m3DF9W5M+FPcQELmpiQ4WMqkh7BQZ2FxCtbb/0lnr8peunySzw
lhwXJBIuJ/NLsr9orRcB0hh2Eeu8eC/krGGXohQqZ8RZ9+plvB+L1d6vvNdahjE4N26aZpbmOred
V4OaVO9oe7GUd28U1Prpt4B2XTK1Ivy7wQvpgUSxkRJxmOlwjyWkxf3vqnpcYg81H85ed7WGvF3+
VddBaVtFjYseDjRPqF7RNGNWpbn63vaIlAwRuKYkXyZEr9+2g60EfPjmB39LgWx/gf8LfRycpZm/
voKTOAr25/vyVvJC1sNHmnIZ4ua6TQDVgzBzK6+2QARVjl1bh7Q7JKxzHYbgIx0asr05bgCKrDrX
cjimTSD6+HKZjBHSp1DoIG6RArgv9tLxLGUZ/KvSsMeXhwfvCbggOx5m+furh1wYKIIosmaORV55
wqcv7t0i7t+MU3zeGkXgCFviBU0wbSV9Kz3gI9H5oKEQLxormpWYxZ8wpKQ3LI/Hferi7ocMoAby
TPMOQYKPEjIIJ70I/M3TGW8TwOChCI2MFGpYOLs63VwZcGKiub8A0B8SjCdTIgsKOrrN3bFA+X4q
DNApvB+E8AQtjMMOkOFmSL8hMlVo6PH6sBiO0QANQQCbj9znx62ggKWxqRhrRxpJG1WeSsJHJWgi
eoLVhhC4S5e3PBr4jxcn2zHfVuuOrJ5UzydbGAmkGMYAFu9FCa4mACczVq7GjyDi0zNdwOYqiqEm
qunSx+HvDvT7nJid2vJz18LMObDG3/X3jCjQRG++1KVLxOnRvBUEU0d5R3DRkCdJrLnDSGZXaJnj
mbczPWG1GdQKQAD2tsIEXHGL44mUnPn07mSP7ww0y4ZGCu4s7lQd/1fWPGWMNsZVuPiCI8y8fIsh
lDenwVdrFX+l/3rZkVp2AJoKY04UyO6UE7QmKqFwiatkHE0RYyJJS6pQh85QJRppGkNWjOmI22vP
ft11FUtQk+vy4d/kQpPCqDKe1xD7Hwu/zSflSAwbXsUmrkrODuIupYLm63Ylfe6hLvcDMZibKdG6
2Kxf38jYd+TJcS1SVxhPAe3ekUOECT2pqCei6zdmsHIMwSXSunKA+9C+pfcfd5ZTEtki12mZTzu1
Umfyja8ECC3rKxSMWO/qa9BwABEDgErWXXXuPjrK91Trz3WWttj3+FgRLIXqIThAs7SMEdtkQFKy
GFSya4bm/1ewqwpJdOJEYd5i8ENvFdATETxMidkgz6C0EocY0iE+W3BPxu3UvuP5LU+pD74drCtj
L3ytgZwBbVyLTXn7Z0pNJeDdbU59fNRFcX5YVJCQoB2ZPtUxa3omnBPdXdj+Pz+KZRBYYKBu0K4i
m3zcZbzsHNtBUay9fFIV40uhQOd8wL/4bLib43uSJzeLLt3E3ax5Z4I8H9fssDUsCWTWs00x//fX
VwcqavNScEpLTi4HfX+wWbfqvG3pAWROY/V5mT0k4hoQjGj4auwV8dytpP5/ZnRi+TCqATb/y7ct
DrKUcZ7antATxsXQkVE90GJcDoQS2g6J1dUVb4a4gvVSS65UZQwEJB6eDBV7EyyqCbiORBNZvQ+A
TSLOGUJPAmBrzhkrOIHhSsiR6sc6oESOZhOrRVFeM47ZZ0TsE9nGpJTdiXSVs1JQakYG9EUV53Fq
aVksyFKxcHx9qbpcG+ZGrWmULofYi4TxdN/gLBn0VeDBerxksW4Seal0g+BziuiCnCCQjwhyCzVP
hYpvRqwN6fj8uEo2vIa6EKqtloXIbTaWQFENm7IJC0gPQsRVimPcyJWyYPVs0W3pjMYoQP6XZvmc
90V0UQ6tLDIi6M48fe9NW9BipPRiISfjxzRARSh7d9OcV20roCzM+/eVu7CXJM80Z6MGquKlp+ID
f4lGbs+wQG/3ouHxJJgLyO4QeTirImlwFxl/ep72vhCBkcrzjnhbQo6xZGZdj7WjsQOMQD2DBasS
k3Mnzoy/sS9K/hpVr50rqQiOhelIET4o/7I1jmdPhOVeA7JmQdctMBVltYV72uE1NJVgzrDUIsXL
18I0bLijoh6XBq7eUTGNckhFBg9C8xL79XPfJv1irxKLyB93NqZ81BKUuxkup3b9afsmlXEntAmL
p3855kj4Oj7Ks6AZhK/489oK5ACJGkMoF3FeTMTJr9/phiNBXaM0ZsqZqihC4X8GVWLgNQqnN/Le
FugFaC+vaRRij3YedG/M0+nt1B1SNO6O33EfSDN5sdMb0bmepiEZqYUqpLCm9tYehI33ITbEsIRT
b7UaJGc7q0uQyvwDNa02rDrZhQGoym7WJP9cqH734Eerwx3XIh5fYsHqT3i9ED2QXDmS5peP6IJt
Caj9TpiidPMYX8WW1uy8L46zJfvWP6Xc+dc0drK4NJCAqNBKcOKEVNg6WXz96U6rDQEkJ5M6/CZU
9lj+qZQv+gZOn9pSPOAtuj+xPKaU4UjA2QGKJ0bbCVMEdrXgcrzcQ7BiRjVvxaR9VGCjjVuS/qFC
CjrJ9FhDsc1YzUg3z3jmLfI7/BlQqsBad3r6fmmTcdkmv2NSXreVXDJqs8PYnAKglu0UqRMnWnN4
5W5uNGBJcSgdb9GJly+7qwC1SYx4AJxCl8Bl8zNNT27SrIC3lx8q/yunAQ0y5LXec1QK0ohDn4+P
I90vplo5m3n6L/1nqGYHOkZYOHspYGxMtFXMuxDO0msQj7H1jNn6xQo7oW/XBQM3QkLx7zWeGzkV
H+fZrk4smYLeaUX3BeZPGQDWMw+wLxIDKpB56fRdwD+S4x5g+LJXUndzDNngJDP94c60t6P2BN92
DEL8/nXjgiLSkTK46yerL+y1stH/o1UcHHhg4pV3e48R/ZfvYrq/C3tYCrUrFzkuS63fgNSEac56
3ty9xKxXRVc12nKtXwTD9DyZNh+VCxrL0UQfplTNk4RzQSdkhyq8331wwbpUUSKTSzxecCO1oFjn
LHdaIgKZq0KqIgB0SRqOe/NpaZWBI1IxDUd6p8reZgvUkmIEOl6EJLvjjfpUxHxQO18FiNM06eKE
TBDMXOBJERUEyYCmpqGIfrcGUusph6UsFMSbsyZ+Orao7Z/vJ/Oa3y+Wys+6WYpDq4vH7GPsc7v5
Y7/YdnDwQonKTmxsYTcCesckC4zNm7niH00MEOYrKkBtLwJpcgJZcl+QbAX3ztpBi49WFYDTN5VC
/X4LiGPKqJ4UUu5H2ciM/66g6lWLvEIWbg48t+flQSSKCXwSKbM8b9619H7ByQPahJ+RajK3woXx
7HXicJeGWV3MeddrGQEIo0CLD7m44V767JrmAzOotranPlCMjxwCysqRuVFwN7eAdTWxc6moKtjH
YcSOa+RNwW3RrWtka9NBNfHn7XRJNj6x6fyxEFIrcOcq1Cq/yloCSnMNZGB8QP5spHdMDhISYsBF
UMfgkkV64PdM5m9zckJNAgrZ/nCQ2MRtD+DEXyXON+Y8BjK9LOe3cqWvy8mS+r21XPYrJFiTdM61
O0A7vLaDSdXiWI4brVBF+94eH4T6Vb+LsEaZytQNP3a5VRj6TVGmFkLLLz0nS3ANjCqxHawxFHRN
PP6aNaPanIIYsdz4h7HeusPPpx5eYKRa6XtjzCIiG8ZiMA3l2YWefa31sXLmObcPSyDi57kF9co/
kFw10ZhLr0N6ybMOCpFEt36PJI7rCAKlatXixILq7ztctP3cmvLj2unBm9WkKfoQl2lxYoJkAk8E
Cn6FCI3oB5hiDtBZGnoF5/wwLvpj1URwhN63GxWdybVLJwIE2RsjRmod129itfttWGGQP46p3cw+
zj1vhZhtpSVukjgmkOLhfnzDHYE/VjNaMGakVSwC2UjEGoH2j/qANndNIds21kfPNnH6cRRDPg++
1LYohC6hv0qTjMQ0tljLzrSPT34h/1He9TPehmFnQM6XWIi4J3qPByUSBTXkZTIB4iXY8coYFbag
Ghk2kmq1y0oJdJ+lsJoadaTu/Q9mjJl+dokHms7L6zIsGh0tzZepUziG4lrwM6hQeFvKErKMoxip
pkzxkxCRR8qX0/FJC/TgxnEF2p/ruFRr9wWCQNWKy1/MQHX/NjvQ6LtQdmtRjxHSyq/9aaZJD7XZ
f2IAyE4tX3KQVYsKE2Dkq7jc0eJlEMlEIzFBPNDQOEBSz8sXazLcBDK5JAI8XvQ1Fc6ztPuJy2NK
bo2h2OdUnfW8cyGTy0hMepRGsvID65HPHXZ3sCZSWkKyfi+dl7rMovlge4kABQsmeiy4BMGs6U7V
Jdsggqp8PQud4REsaSW8Ua8FiAWBL/7uW+ZKElSdpCMB4ujHF5lv0kLE3LmqgZVYh66/ylWphhUr
amEjXacpvcJ7kI1b+ocT/MaFkIaj5JAl5gWR9M/heCyOqGVPJkNUIZmxKGE7K8DlVLu9IlZfAslN
tP2MYq9moqWHCxoPL6apz0FsYlg/ULmAd3yEZuZx9MG2Y4+ytGYkeApMXR+gQKduZRGo5fPM4ww9
orp0lkWcMuEz7ReT5MpXItjSf6RSbaTjqCpb4HhrIeU97nA24McBihnJ0jFsCdFq/CQ5YWXeuZg7
7BfKz91eufbCsz/7peHvSm6W7KJ73+m/7nQS2MqdEbgUmD/rMBGnIycLYRQwvrJC++GaUlF6XDyk
9HU0rnzEC/0v8VyXehsKBkmd05IGlP4fG4UYQQNEtgLksYNHiZI0QYwezFTMSzJ87fi+65eoj68C
SBoBqD8RqFG61Tezg4OrrTCuoQDDrkaWl/zLj/M7MmuWXLQOoiw9/rC5eMZShGvhAqLIazHSMP+G
6r8ZmrzWm0EJJTSCeL2CUI9ZhQ4gX7MEqp7QnhPqPQ0FBWbwAq3mrLyZJGAJBYKfXYWsFqnlsS8+
Iit5balMgBtm8HxwewM2BuHwt/VAKAvXGuk2+FMmqh134pGCdZ1Om4B+jBT0c3UWEKpWlN+sIAdq
xLaIWJ2aVNnaEtMPskE9EcnAIumSxCqlV8vwSdr32zE8MzeqKThI0tQLG2cs/0vu6uCg/XYx+w5V
yX6BII3PWu9xzMnuGJJX0t1zLZq61I7MvSxZ2eydrkUA4ULiwFN86n+4nVW1o28xeLaqdsgpeMmd
GUry3ZkGqx4uUDtCIVXgNmCUdV+eB8zA1xVMxuWvmGvVyk8Q7zhHfIVn9g9SWAU9INydOlLDBnl7
KZ+gEb0irUBLNDFm2hS+chDO+B+sAdkMFBsloPs7IBr11GjqLcIyhlvYtPa9J756zwSmGEmQF3Ud
jFEHLX/SpvCxoSO5tTb/drlZ0FNV50jO1hVm08SIkrQFAgHUQX8aVBCnil/LlxvvUOKJyHRok8IB
yBtYjMQGZCZcXyZVfRo90Qx6LgP8Q9w/tkmSz0t9AD7FcnuNrD6tKkR5QgZS+C7QZ8aFXAb2+Rg3
OHXZkMgy/nAmq7YOM6NBinE5r1/oIHjl94a+AQiJlKAdCrw4kKL2ZVoUebO6YiZMVVyURa30cssn
N+All8bfNRK3Vrq7LTpYDirdneG9S3CfTCUZmJSoiiUp03JsAOFaRY0qkCjxBL8P2Uuvf4n23QoS
oJajkFvDhdrzaDkm54L68ZEINoOOTFZXFW+xXwrTYmtnP4/RwaS8YCm1l2GcFnPc4fLeltdFgNOc
Ev14JbD+qLUILIJMxhTn2ibzzweKSogQ/i+y8xvOtrm/0Cr1HfSl+UgmXeDz92CMsvRplCG+UXp5
khBWznL2xewL+mQitlwn0SL+PG4xr6I+5F2wXE+pAjCIxDg+XzS58HjEIGa9gtOkcThamHPh2gxy
eD8ADKjolIdf6qrzQPBj/zneuXznwdWiV2F3zE+/mH16dK1NzPyw8NTPgP5MxywojRtkS8Jyz15J
2mhgN4yd4EQfnJ5fBCECnoPTW8dJgqgVYKqZx0wFm1gFyMf0kjVO5drLxGVC1XW4aDSuDitbLxI4
QYHI1jddfggOYO585jXNyIk2KcudIYzPl9JY8P6pFm4B2R4yMf0zx0ESzLPajzQN0mPjmzI5aniP
2vdZQwgkDr/S1zE8Tfp9HzEoEg6iVZgVSM89T0PFWA4r3Qq5zMHO9Xb5uuPb11UaKkLucrC+No4E
paQ29YjaPS3nrKHA/tDtR4g49U77QOpBXbIAI7hi4Ud9FNHecwD6LDMbJpjSK1xvXPuhOa6u4XAi
UczJm3KapucFaBZPtw2kyOwP4iLSTNHDB122bdPb9EfLVTz2mp+uFhv8HnpjBxtxqfIcrs1rINRv
RPBJ0eoqWms/ALjg03MrhQLFJSDzJE94AhibNWxRHyOmZoMBXq++s+XwdLb9QJ7eZfbrwgyjS0mb
14Fz/q1ZkGTICaa2wLojJ91SilXSf4AF41YQZMTpVAr39dwAqvnzNkMf0o1CCSkMrP8FGPsW3HJV
6fQpIKrbkLfW/kYxghRxMOFmZkOaiyU6fc4+nZXL7SLvKXJdpTrRicvMHrB74Dk6mgKwvcl1+WQL
wmz2ra4Uy11HVGCdHUoFDdMe0J0NEZ6GHl0DgFoFRbiukPKx/Jc2PTpltS0rQxJnMHU0HrffCnQQ
XpoBG+Mwqsg/ZH2B+2hqOgeR+MyCNKiz7P9sNqgm3o3s8aoHFPZ+JrkCcHIKa7D+p7u9vMNQvyNQ
pJ1Dj1+0jNBTap9kYYkFD+NmDvkEVqEDdU4Nhz9JRlnCNnzMBCVukZj7QJlbPRgemxgw2H/4BDAn
tXgTcSLSh0WRtTQAiHayePRpoLlEE0Mm178zBBE1Q/uQWYOq+gMs4+ERDQ7LIy6kA1P7tTa8Vlnj
T9ofb3WkUsdQIud7kgRAhxxNDuRMGk7UjAjWkMvaI23d56DKQmgdOXh/hJPPp7i3nDzVeG1F2lVl
DR+QXxGhKcINOHB0Zl67ku2e2uhUycQScpYs8PlZDe/L44svU1cJ867/dGCZ4uR8tVjC5D5Sbq1u
Jn3+key0ZKh7xyQwh/TDBHDpzEmZbpiuvhNb2p5v4B2+useoKKd5XaHjXcnThfgqt0vX79orSYfM
T6TWVJuGbhU8fIU2FtT+oyNuHQ0pvR6y19Xi/3EIjFlbW6CzUji5cyTjyp5y3zPQA5a6SOkCW8KD
uNJsPqi2ZUrUowQEKYhlLDXjw5vad9VBcSEV+TBC2Qk0NFU17j6g1ifHnFU1fBcqqsAPjOG6EURr
j3jg5titEvrd3yE/lT8nyGtQg9wtJBaK5ElpoWd6MJAm+hBaHKLjzXdF1qg3ywnCKQG70IQCNksJ
hRxGLhOE0btzDw/UuqXZ9R9iFC5QJeuATXSqi6PMI0XRF12G7RVSpcbuO2COkIZOpKVuJ6/CoJtw
Q6SF7AmCT0swQLhRz2iGy4ZWALILKQafholOeQCreykY5t1ovJ4vCpO9K1zLuXJl+vU7A4gXkBQa
2wFuy8JW1M9oE+8q3Z/1SWEyQsyDIWBR08AtqMLnCf5TcqkgNlAL3Mke/W2zuSATQRKQCkj2Trq5
A6RoC7emtPmchjuRcZTfG6iCmeeolApp8kbbS73IvrOyW1NhDO3PiY4InPdxBGrw1R09TpgQcpwQ
Xj4IzcwMcIZt2eK0ioHkJ9+8CYbwtK658B4HKRbrbQmmE1Pzp6qoAI1XjgNXcIKA4oXCz20cvxJJ
7R5j8DGmPxNoaNrc9LGvWZqJMEKX/eAHx8S1llfPlCAFTJlbq5PJDrE5Z/NsqWC7nKB+JjaGc+UG
KgnEgy95iYhcjQGD8yWKEEUeAu41Uwfhj+mQERoBkMypb8wn5MyAoHbgvdITW8GhVnsJcrAHivfW
1y+Idtb9sKONyeZNKbl9RikKONm+7w1C1dwziIULtridlPoucsuP35UNIoDYP8JsbUpGOR6vDA3a
3WstflKNjBYnTPW0b6AxQhcRe6PzoKc222/+QXKEvSAu6jsD7YKHw42jOVaqgoWIXBESA8xphM7U
ZmkWm141MlJYvAvlMToIe/wD7AbiZdN+swu+qIW5y1OkorY8nWTS3hzFvXZ6sEsn+MBKKbtsB+Vy
xhJCu9EQbpDhk9ap6YSUlG17QctSldYMHzOx5Gk9k2IwGg3khFoQeLfjHOaIfGr2544dvyet/jNv
/h5o82wBx36162vXPZZcEA+q7R088T76s6+i6fU0uGreTJypxWfTqWJb1irsrJdVK8eb5DQMaNUe
wr4RNSnRDmsJ6+zguNWfE6cbM9rojcpz32HQZ+rT+R4TJPwgmzpBrl2UFKkmmrvWVqd0N/jrfsBX
qxnyD1hKFiwcAijFqQNaP0OEtVRLy4mHcJ8fgcgqA9zWDJvR/4H/pWiHWYvvCJHCD1dB4lLtoTyN
X1ZnH1qGsR8nFLBu2nWNU9ps/OffO+LFOW0RjY5EgMqyn/45drSLAdwMPTHKSid2sLJQonHMBhK+
EMQQNBG/Z3wWxA3COd+YVxG4XpVh3W37IAEU7ghPWvHHxKIqe7tMo6vRqoc829tDEbgtfqFx2bec
Bi0M0XVZYGmTDcrIzzHBoQ1pg4Bf5Iuu8wL96prGjhZkycY028//yoarFTjKYh/b7mNTmzi28R+0
u3+cGhN3kp4E7JUkRP902dWmymHCDXRegl5l/a8vqgZZRZI/U0qLHf7wsMIYbhVIIvRWA7JzQ2BF
8/yLDc9GXzLniP/Y/9eT4QoT4ribXx4xb9CLgcAg4Bl9wnUQyB4lbjtN+iKzgt6DlI6Ab9KeJt0c
SAklXjxjWoKs8WwzDtzxsnhejZ+zqxmmx78+EN3jK8W/pa6MppZdiKImfUAyb6bkxryupK5Qj0Vb
T9BlPYrwTEcAnSjB1ogUuYatq8DqVPLe8HVCA2O8mFHxy9jipeZJdr5ZEABDZ02LzYG2qzbbmLy7
9noVj2AoJ0m2+1w/KzBZjuQcl40r+pue06zbLGu3xnGK42rWZWi3GtInH3ryVLo9msq7J3w86B0m
Nge/cwhUO+8ambKqYMkUSMng6zrxsU4mG4+OcuBFJ/zqdBkaxhWd2GfBnmu2+rQO1/qhQYUweDjC
QP4mub7HzpdrIqXyCfk0ZWj0GXVRHOeTnak/oenUeLcE8ZZMF03iWBDOw3omR0iTEXaCK/lgOGdB
bVb7v25AC8mzKyttQds3Jga1eCgKe+NX1SN0X5tI4QcWgN0zHlud01vl3HQCDEk2mdQOZh47My+I
4IsDEW2xpCl9KZJppqu0TX1oxLVkpy3MiNUlKrVLA+DVevC4iajZKmUMyZCF0M84Nu09iYyQ/cjd
iaIbStGiLZdgh9+4h1P+9S6WumdMDqFTr+N4lxq65j7JhcP61eB67S+Zq7yWwyHCNoU5TROb4Eop
fGoPNLOSKizg6YJlGfbhp0QelaTZX1MrVWgMpGfobEux059LPBy7R97mD3AvK30M1E4WDGnHViau
d8Z3Csl/CB+CYi6Z5cWFC5brfaWyYmOOlkrpSeosZ5OKpb5+HkZ2d/97T8TAeZHDJrvIm6cTEjlV
E8BPNmwx7xwW7Ghti2G6jTr1yFCxgmVo8simUjCwmCOX5m0YxMpiB6I8+Y+ace7Jy2zlpDKoUyeN
Jvg9JMW0l9dN4hDkwfI3phhDS3DzKq0bNnU/6j8shhLix89Kieojhop3bTcwZDxADE2pG2ZrE3JN
agdp884lT5VkG4Tb0ra0xuGGhJvfwSH3m/fp+Av2wleZuXUXuuQyanFyDg6r1k3T3lThiaUy91jo
cPWlemMOfws/mXoNSeyFYunRp1LW5dtSh76n4iCvaBkN6z+TZBAoXkqSS5kvu8O6o/yt/d5E8uXZ
7W4o2UyKogQ900X2u0EHwN0NSKZwLccbBkZweCX0kp6RleuFU23mUdJBm9mg8p6ffVL42CpCv70U
ybFlxvS5Chc9raJaCgOfGzDZTUo45qFXzfEpnQMNHgloK2KS46ivJl0myKUXmhfaSor+5KbjKQat
w0eOitYodRZKmqtzCVE5SqMULr+VcFrTDCVWw4aUSOUGKsdH89LhIyxtbn56CrEpZRF9KzvBlYwl
b49KHBFkU+TUJNA/aHRpHEdGn08tuVuMqG2nS+BMNaFT7OiqgtBaf+SQ8Kg95RQB8vMA9Edajygc
7pGaPHgqexMicIOdcCDKJSpw6GlUJQj+rFEuLTWr3wjyxy1gRDSFCANjfHK4QbgGnp/GBQSWGA9e
PZhkrBK+qCtL1Pu6DM4/Z0TsGxTuSXLycnOJzV2wTuM+ZO2CkzzocEAxzp98isEqG7xbTjntlXSB
p0LZzksLtYFb+UOjtW7a7KGERO7jmcm2Je9JEnMGf1hCEKZVjoxJoQeDTjCGFi6bNhvA9+zoN3oO
SS0aWOJpUL62GRRYJPCXX46nTxHCU1p2TMCv82HSHyXteSkftriTdL3HHDekDBxQMxaQWVzpDDdO
78Swle+31in0/fddCVqdyln4DKPVIb7ArAzJdCZL9zdLbg8xX7Exn7ITs96Ixkwtfj6jdJxdgFw2
PKO54DxEhUL1O+Dgt0aMCqTdeDI5zovasT1M5fldXiLSyMofgOD3jeN8fig3Y3eKV5VjDtdhU9Cw
tTlU+cnlGM+hP25+yLgvaTJq4zWuI8MGdcLiXfhTAzGB9kI4DhteX/EguW/lC5bBOLWl0aV0qNSo
XQS78XWZL/XZBZnFs5T4CBotyWymswXdL6xlpI3o3a3y0oWYFfpLhjuOSI3SRQ5Qaa0jKkUsMUXD
DNiL830JihzM1jzra+5jX5yOuThJ8Yy/Jdlm7VgzpJE6HecxPx4Opsl8zunKWeZWYA7nqS4gcjLB
jxWbUCsZOCn+7t6aVzXuXIGo0R3Lms6oAC+hDbTkX3HvCXGkcNBWaUmqjIIsUBMWEqLWs2JsBiKG
XVyVpDzfgGapSsdyVuzOFHqnt4LT4cNQ7a/LEiauvDvnsMHjvc4OxxNAQxTxX57tLNezjhik9TWe
lJKr5ztiL4BIM2f3YdRM2UBYFC6sl6ihWBKmvrFbk/Bp5xVFRJ3eRhqRp8FGqxpHukjgChbSkdJl
OPsQ3xfr96cUWWH0VO7jhCrld4Llpb/fgQInRle75ls3vnm2ZCPFmcDSg//b0d57VK3ObaFwuLTG
TGrHUwgkBc5wv3OeXR1KlT/c+D74OJTkrAjVnCc7lGz0YZfBoWaGiWoO6M8P7eTdQLqD4R6ennUR
VaHNOa400L6lwpVV9qNHtgOmi3TB8oD3WziQgOa6IZDS5YvawdJm8v6x9eWvWbogLzo5oyIXXJqn
EfYf+nqoxpDshC+Sr428AeT9hX+XEaRoJF/fMrJ9LPlULKUeiKvxCZ2bJtGa+xpNJXrZ0HsWY3Q1
Trc9i0hqj6QncTV7iilIAHbnvPCh2eNNcHZmqTZCWnaXD6NTXWbV0cXva++rDayZoAPQKojoagKJ
KlqNyk+u/gtj/RvG9WkgrIyV4y/rFZBzewArwUHzM7PCQl9GE8+VnxKzAy20/Kl+9lqsxiac6lTu
8ZWxhYv9tAol+cAlEGCGyRn5phjRNpj2AHuUYDWGJuqId3nCaNjnxRCIKoXWWFAUjZw4Hu0hDYUL
3uxxlfL5GJ5b9xGUQM00gOWbXWLE6lvBUtNt+zV7R06TPyKi6lnMAmTca3q9d9kag4ONyBVcvVHY
ONMFKrbTKJ0qTwAE6oMBGalRIiQdvm8FsXqyRvZ9/jStqcjJ11fOTFIsGnMHQ7Bc0AHenK7ug0Sv
Gt1qEHsQbeS3iHOhyYDwsvM92jxSRzAkBUsBcoNp31/4lbc50Rj+UvUvl9h2zYUYmbBJiTMpvFRh
iOpn4MSm43KdAcSy+wcaluR5GBJUc/wWulKU0U+jeBTWhO6sSxtE/CeeaWnsAWYMlC6vGgqbh46x
+i+WZKKAGOcgx1W2KxS03CrhWSPCS78l4AAMZfU4wU0jjAVyrqobMwRnNCsKBqiuOG5aAt0Ud+SL
RNOCjy9FTXWdJttoQFaFX5suKbkKtfmndGyBWkBJvwYPqQSN2dRixLLG8RCu6GKx9WkWNhhtTmR0
DJXZeKX0l8ueHXYH7ENskIS2C1plHGsgXGsOkuFLg7Jn8ByGgqjJo9NNHPz6reCj5DAU+FaXDOHv
Rmwe+cUa04QUJOyUdi5tAsHEv8w0zzs1jObyVvon/viRWCWA765FC6qRN8+yA3rh2FBlACJQ3nPf
hAGxeBFl1GiBfou8j2+5VHQWrJ48PUi4jP482Xkiieie4pFnjZvZNmj89eVPPjxlnHPyOimGfRYJ
F4r9ESHiPksEsSIc8WuTMpWxxAzcdWdhfvu/TqSSG9BH9BPheNu3eCKX203W5sv/4ZhnYtjzImHz
jRteTJBLHJ4TiX9Tshent5rKZekfU5/YlMTonNkBkqBYGaDuj/hYhl3Svh1tYM5RUEROm1GQ8DYF
rgQHVZZYyeid2OKzdacQYDfbViIl6SQDZ9TW+oEHvOQfLnklSukkq06le4FP2scsRpDY6SrUj1/D
3npMcNcr7mhytvjtM7FpKIPrZmCX7qiYPk5vWgUtwxWs8lU8x2ttHxEpcl+R+A5IS0hUA4yC7z7X
gRkFql3XgK3WpCe8n0i40KxvFbdmguHDbRrL07sOWI8JKftdDp5bGj6nmT1LHrI7IAecZQmc/WSL
b/wmlkHIXH7ZxqtVpq+73iuYNgO0YmNdA4zDQ6GfchV3tnQGDx9LBhReziv9bHgKp3Hqk/GKYrO/
wL4vmdj4yHsxqjT+SlVl0BCkDlL7lhRMvzEznU+0VNI4rEgjFUwaApMMGmoiWkzlfNCYGprSWDki
LAb0/uNvoSL9iZdrH/GuwEwdWLebnPxX8IVvdj750+KEHN6+ih0exhX+2ESd3aerhpt/ENisO5o3
GGg2EJ89K61sVT7mwe+NqaMAWlBUEzr+Txo3EdBRdAhzSkW1iJnvilyz7BuwidpTmBkJ9LrugzXw
KXaA15Wct0fo0fSM6LKcAvKGeLzozPhEQC6zNl/7crbTPSbZ9vm9GNm0SSB8M1jHv/3ajmvGWw1B
KYFLldM26taphQ7JiRkaqswZRskHoqGAMHs1+nqKew6yu2gc+yo+Y9VGxfKG6j4nrCxnK3k+G1JG
g4JikI2bvGQkltVKvVS/TeNFhCu8e4uSSpydyUqwrysxEG/nHdvHGSupeCXcVB5fie/8czk0OjE3
KsvIrrj24E54Pzn1bNfbN2JytkosT8o1k0H83UmKRxhjKluc/zH0abpFCJzY5/YnXPgkF7YvZVhR
IaK+1BtZbJh2/oZsJsFkxrIiti55SdPJ/SbeaDSRwC62fyu6gc+dFsaEysQYuvgPZvoEgGH/Ye9c
bHiPa1z8EOySVgR9SX11ydYxbRHbsGE7qHRyjQcvyolpeqnc96banixcASrQIUFiA+3ta0BR1EPE
6WWuErP61gvQvx+XLz8/0YwrcQdop6oVqu9gq4r60/NOXhINNZaYuVbAfxkiuywpIKH/XXKtuPH9
VdG0sC6bXfHTK4WhD2h88ibtxA7aTfcUd20FTXTlcXqnxEZz2Ose4PweLx6o2fCH5/ETLqJZpK/V
uVy5TaNeGUrSeHHCm0n2kDr9n+3LUABW9Gi1iD0XSjJmW3BN/UnwM2Hga/L5G1+WWGyZzjkUG3wv
T+VVg3fRzDoZumFP0ZG6ho54JqUaZN+8t33v9wyTPs4C4AjybIXe9MMCQ2uuvVv/fRsZdcT09AW4
MtdwJjMUs85+C2XWUqJGHh8cc6nuvFjV4WatfzYN4PDUxNZFDxVEVr09ex/Y/8nQF+DOuhIY2zwD
H2Ylwn1iJq3rqSSZHcDD0sTnCIdMiG6Oww1IZIpKK/hGwpoBs2+mfZyvi8+1JBVGlMd5inlAhHDP
dvAX/7hN3ClQnqYZDkVSn83Z9vH7I/Nxp/xbu2/zKy5EtYKRSxJGOmR93vXygs0WT/XwU/8nUxii
mpQy8xQs+pOU5abhvgEbXIPpeQ+5MhSQw3lXKRulde8fwDQ+c8D7WcdBCqfYCi9LJ1Yest7mL/BN
y0B6+lWjfyyTZ+C6HmSzIds7TguPaKq3IjuPFXOLQxRFdXu5l6cepMGITouyK93QxzQ+yZ7oaW7b
R0Uabs/tZL3pwuvnzVrL+pCW4MrSD71jaSKIQh8i2rtW93PU7GPvGl/KS7HGUGjv4aoMG9HfEMOA
jBB8cWdpBAtcbEnSEP+k0dkRDdzeQQExPttCLkrnWG/LIjDAGO3VccQHDZ7g7hHmzhn429KOiYHB
OcoFEFbNQ5CHeepoM+9zbdpMARHoQcPCbch12tz1Cvv5hTwyno38iHXlZBfBc6kXL6rsF8294D99
lYRrpdvMgK39zDKausHNxKUPUCFoRtQHLTvzaspmwDiJ6lqbERQf2oDAMzURBf5w3cMoVIks4puU
bs22c/mI8Bg7/ABKOcvJdgxAB4csmH0ZIOdhir7lZ/CxYF4Llwme3FAHqYoW0Iuw6PeGL2CXCR6w
hE+mhxOjj2X/pgIVrp39N8Vk+OkWjQQvWYjlpIPNvAhi6upncb9JN7O1yEnzDTn9gjPwuAFGYuKv
GTIWKVtbvyepd4HIayP6YFNizR+U26VyhGvtO0R+DsCXr11UdTjK8HXy8TWWbb0sssr6Wgmk+QoQ
Y/wKBpJsqj5y0nQNIaeFlvaAuNsp15idx9X2z+rzwQ1IV6n5JMV+TgjoTT4mc47Pw7V+ciCIWbWo
2z+k2tdYYm1pmqPfgw7md7HZwX8PgU1PaK/+530iP7XWNt1/Sk2wxYApaApkdpDUh9GSDwxT8k5e
bsNZLnCltswXvYHu4Ef8GLVwdJZ4cB63qFszTa1TKNbGWmqSSxNUmF4zKRXtDdkWRl1g7LvELmN9
kiutIBAlKrWg+bAOX1pYNeJRlKaI5UgAAKkQtVpjujWYz7MqXwjI5eA31YP8HIvFyyHAcd6/9mvG
VtsxWR8iLCZD9yk6ixX8oddXGT/HSDME+1Pex2Y8RYQtJIpT4HIIvBpJ1lB8K6otCKetbLcnAyWy
HXPJo0OVVVz83j1/uOy5XJMn0OyvBdRvvWhqxu6K1ZxoJuiaNWTyWARfQz+hPHexKNx3t2eUXTPo
iSzA9Ds+jWR6xQFnSFWjrgqX5kFUYEeoBNPtu0lpJ+B33FYp1bUpcFg65+7fI9k1x6NPWyxNRk1J
twBgJDCiEtseAPIwCTA1nsAQ+9SB+IUOGqyvH/fPUUcIdvsdRnseVzth6ePE1VSSszxTegS8GO8A
ribJK05cXOsC2RGy3MJKUwll/0Dd55VMsVPRlIZ13fiAsgxwJH7e3EU2a2ACMWjWgJ78Euwa1oFP
kXsX7kykZFXXDP5oAeN1Z67N5dSo/BYoCjdQg1pK7a0hwTRzsgYaUw/VjbTX6MsfiUREQmuCqlw4
/a33ZL8SCbz98LicjcW76uYtASOOedfkNDqMZW8Ast+nt6G3uPwSthQ/Hj9E5WrrQo9ly7EqQ+N8
AKph0UWbbETyRq0cd9Oqv8yeuqX/5mXdDwXbqm8NQLi7a4L/GmwkP44O0gXkL3EJr+XCw/vAOoG8
c2+SLiobec2mAst8ekl4VLvdtz/I+UC9ZvFftRuac2QdnQF0Fpd3VREc/tWagv53Gjkiu/shwo0x
FU2XX/zozQmQWEAD7O+lzBN8i/BpeyBiUHA2zkAz1WPPOzbGBRUd3cju1gEK/uiRf6/f48Tw8w97
7wtqYEC67XLbJ4x6zX3C1Jnz9P+ALYJpzWwxNm7AEWO9mUNPbSwvc8C0WBLA+t4AlfwSOeWe20Ke
p/Ck2Bmpz9N5OXP5ddO1LAPkAh1ZFCIKy+NLzOtnYo01NybSawVQiMse8qFj9EhNkqEh0Fl3XdmQ
E2C67GC0Y31PIxcbhriAmyMFsAdc2+JEJlUxtRv2n780/ziEY8dArGZn1XGIMlnzllPDVAsXEIYY
3CfLA2J0QAdN/5XYRgKfSIO6QqgfyBaTlqcYonSvvB9sp99jNS38hq/BzOHJyeBJOdw2nEATd5WN
zGl5nf6La5KHRWVanvXN7Nmb2D7OteYGIo5Z2MA04URZVR+pdZjlIvkgcbPKhy5Vs+m6Q0r+hTd8
9+rGD9OpEdiIAOkiritLr3bSLuZlP4eJW9Y5nueSkZ8PPmKnWs9AT/gJx/5H2BaMzaXbLa7VtuKm
niAmndMnd5za/Cg/FVM02uLCGnYdJEycDFlkBuG7LKFu5k52BfFCFal+MTBLM3IEnRYqOsuekTCN
/Y7Vhdmu8oXLuKwOYDlGb3857xswUW/JiN4u9Fc5yOA4wDJAViKKFPQwE/suyKxk8AxughNUhT8B
qYQC7g48OT4ZEr/HfFInZWNShwtTE7DImQYsNI9CCh7lHiitbk66YzgYk8z1mV17uPhLq53yKJnH
XLTbU+ZLXLG2ivyUkJj+XJH5/vXd51cWikI7QQ2A/G+TtMCP6f+mUXqWPnEH+Pi4YNpUx2VDINQN
nXyPTDY/in6ypxUkRJ6lRQ9Q0mMBAKq4TAgZjsBp3xgtWjr15Nnd9+YFH4gssGQYsBWRJYyTn1zF
84/UpdHX9pwaOp0sXrMCai8nSONEnFZz20zkl/D4jdxzz9MrbxWjyeIOXSZpU6kOqfKB54tses7k
Lh48LySrCvbtOkGaOA8Ai51TG5u6iCi1VPkREzA9NJpU2fnX6enbTPuO201s7H7/76g9m5ITVilN
W4J936P9LTfEj06xu0zBuI1UCga8LxhtbvpwR8JxxKpvZcAIhUqzZmK13jAAPM12Buv39ACWBY7T
TF6a9Lzx4hYmBpjxiDvhW3J+3bhNVRJ3GU/gGFSqRrUXjMUCa8f4Qo4rQjQuAGBvb5J1CBmx1Gb3
LQ++90g1+DS8VtIrUMLypg/py3c+EsCcfwXwK0hKEW0yoXCw7+ghA7taqB8pdBP1AAjd72wXNpYO
9AxIA8gz8dpQq1fXpuRUv/JItQwenDckE7YjVVOWY8Iq54fGB74YbdQkA0h//733ZxBNICJwvnqA
l+AQNX7O/Xl//c6swnqOXe32iWfY2iVnNs/1dTUKAaIdYurEykV9fFX/Oe5P3O5VjJP1isM7CsWF
JCiDkYLyAZWs3A9YN29d1SpcNklarMZ/EwWjnpBZ1GiaUSMLJc1qjFn7y6V6TmCcJZnk2leXeGx2
iwUesawTESJNrx8KBhIq/IqiqNilcBgG09ilbL73gJhppFn5wqzrUxRV07EORl2sEPkHt/tI9FaJ
EPmizmnV8eMbCES5G2OskyOC9nLF+fKcFYl9TvQq1NZVTkQ0hYVv3Zz6nIPfQWV+VGneQeI/lFJG
TporKmQikSnPDWs4LNihG/j43HaxmekYWSYCTP+MrYXbGLzQkQZNgboWEnWgk53m4GOULXVfW2bH
mDhipwZciPpEg4vQwPNZblAYeAPlf3+g4Ips3ij3JMJzH7x69nEl26y/B+98/NV+OdfbTZ48XrU6
KtM8UyboGEg2vb0fVkPiM9ZnezOGdxaqHkmM6sovafVbKEMszUsY0OhdYps6rSZqpnTab+8L0Owb
ukjX6+lT37XJE/U3s9Q1//rIKWyjnjnYmzYZCn73Ys/YcTkpAqM5U94uT4SZWN9HmhOpz2p9nRpa
c7zPPyBhiMO/x/00x8Hwf9AMm6XwWmpXovnw4xoxD6ZIwZzZ0cFqKJNJ8XIeJNVK2kZaGPkImy7x
fvNbmSTzHeKAS1Hwr1Yr5l+qVaX1caELDlEsmwccmd+7wTwq9SiXoj99EHSQ70KKii9XSvHPR754
BSM4fq2zXuQO3pkK+Jc4vpsmn0RbfhYpTOWOHjc5gxdwR8+BLnJ5Plo+2WEDsiAzMqYE5y8E+Iin
ArPWprvnQE9EaUIW3e6MshASQ+ELUra+FgE7yar2/2GUE2zV61BUIr16jEFlTIdYXa635YT+fSs1
XKj4MUMXpSKsahDS95YbnRpQ+nK8/0d1hQjW1nvPgrVZ1mGSZ6bA54q/CwFzwW0L/UlZ3fHa9f4D
1x8u67RIKKx23I/yeQICCvWkq2H63zEO+GImixXq5fbejkfmyscg+qDHNrlBKcFscXsTFM2OOtpW
d4+fSg0ImU6oSNxBLLn8C2UCpIxTJ92OxKcPfk0GO9b/tDygWXAbw0PQHnN4aQvYQJxoYmgf0SM2
e3PtfAYM+8ZQ6CrT7Wg5ssBA585upfz4Mw4xyFIjUIferoTvaB1RaY2jHzfRR/Do9sgOq7hPPbaQ
1n6Ajk2BQlU9WIzTnxz0kVHSOevJ8wzPxTc86DQdXagl2RZhN0HLWs4GjAGHRVVfmWBxslP82vg9
PzNn0XKiqNcoqQf4uvP/D7ceGr3XtqntKq6f3PzP4Vpn/9fj6kcrYaqKvDLWhJUfVcixYLtOHQUU
QR+TyC5pW4pOhbQzwpHrkukKdpgHlgvcR/ee4M/gE8Z9NHqKJ6Hx89d3NPw/Ec8XzlVvhtru40kO
9MiLy8Y9nEZ7O17AyfilmelZq6fBAVL5X0xHZuL0ki/kHCKjEWi5l8VwGLSBGzhiGRyRVX4ddyoG
sw6w6aQHf6GWRzeCDiBXRIEfmKysjgB8qsqEiWoD2GVOivOVVbPBqp7wqW5XolSCIxw9jr2KbYJj
m4/D/I5n3rf4KgsP+hzAmXkEDjzs2aniUVxZIStyDNoeOqmgldZEgv/Wl1NakwpUGtNj9rjSRI8G
GHsBwG9+ncyDhug3cJg7V3SAlUg1Su4mT59CmgUBtJI1trlUUvP3uNhJUXxZVkq+AnQfXhu7SKGo
i4xFo4CjE9ImxoCyUodKowcdj4u7URZrlf7b1pZDbteO8LrjWfu4jITlS5y1Mqgud1uIFhrYzJxu
T6Tsmqj4VVv6A1KZOpQjqv0Ovi9wBif36SN/2zlUw6aOCrvGmMsa4e0k+ISsRwQnV0NWpoWKy1uC
OXNYidx15PCuBOp62qa6KG/lAVEgl3tE17bPvCe+iuPc/BqT+qh//XbNcOGFTe41ufQ0OOcF6jzR
S9YJRqVAW+iiUN6A+UE19iERF4HchNiNaNTAsg/JLBVmaaxlknxkH7AF5oL857aHGHl2SfF1H78d
HM8lGg6U9wKTcP3E13WV6Hql4f5FpWybzzwWi7zOdL2awlEcKrsAsHiLHIWq1QmO//nAHnQMZ5j8
NpRejzPXfaM1pVmrlGICNhRcPjqZx0sc8LHYnvakJUalwKv9UZG4O0SK1+TXy1u7M0kAxpItUY55
UpwFrV6VEEQeizSGME79ki+T9WVlHh+y/KgShi9Tzy6sRtaR4+XElFniirO0tSecaeEsIsqfhXt0
o4i3a6zKW7kQ65xt62o5dOjmdrfMzCqgPeFBo+j93WCxOisxGUC4aivlBKoq/bp1iBtVN6m+NbiA
ZAksSl6T3fgcYliaaZVP6S9yxbJeFga9TEwH/8irhfo65hg4lW31WI80UCFr2BQsfxHiniAiR+/k
Xb+LEc98uBJqB3ohWV2QyGCOxmr2TUQWewkXDltLxDrEPIJOWgRRA9hBlik7Qt+Li2ua5PoQM+1K
tT/Sqymj8fmEgRMYDOtAflQU6y85XvnznuMQkSXHdtkxob8Wym6MOcHaJuoQfb1Z6FrKmDZeCS84
uPTJpoIbn0s+1yka4OrpCIb15bctlm8/3t3CLIEosdp5O9sQTxjwFp853NUi/dUF644un8utnrht
Ys8S7WxxKJgnEPYa6dCvNiiv6VvZJNRnB8cPdxBueFvP3DaTaO4FLcjBkYwdI3v3+11zmM/4WkMa
nPn5EzwwFgqV2IJEkCUZgH71EV8Nz+QQ1TTuoROrWy6QGFL26uFV3DulBelLj9Q56WVqh5Kp+MD+
0y3g0FZlx7v/VI5jS119RKg5XZUPtfV73vPj9lr9BbDlArrDrzJa7T9FpphRcFWIeZlknRzr+fjF
nEYrFra65Bb91OFDZv3hmsu50BXbPGZFGhT/lLGl5ztvbfrU/0j8krqaxTJil0kiJffkwiOR1PVV
4EEF++u6X/jCnHZlLeZ8O9jdeYBjWKJ5BY1PToWZJ/FbvnwPp67roEHKfz3AumBmNZPfIy83kgs4
Th8eM1dLQ75quhlPy/o/1/iEtxgdpFWRWhqIy6kqGeF01HeX4oxzQg14TV/m6bnzg21W7pHOkyZt
u8GIASkHOb8aaahBlibyKf+BDGcYX416RK3ReM77ZxRtkfPJEnT9npVkhQNcWRR+GwVfWwIEBWu6
B4nvKc2HdqLkBFBpVSS6gXLnV4NEvh0uO2eLb7hgUslGJYgI7z6nPEY9P3bRes7dUqiGkNsauvIl
jNOL5pnTpcghdnEEseRUg69X4roZsaVAvRKPxIlaB4Ojhz2PBqVEk/H60T073hEh6+HROo0xu3fQ
GDnVjnPESUMK3tUO9WGUfCJCrCUFPRX2BbSKYLHFLkFjHWNmQm6L//2CEFn9g2Wm2TbOwmwRxVeo
w6CCkNjkHalhtJ+eqWOdhMLJNOwxhBVrJpMZE72Ny9uDBH+/fcPspkzkZIB4LpA8QX9u2XStT6HW
BURLdnm2kSrz1EGMJlXpvczrb150Mcg+ikJXrYzKoJ+qcgWgXvBx8he4uAejIeEF11j9NBwyTWCe
S/SrTwRmvtjZ7WZ8HeO6dcvv1Dpe38g1/8kED/zwmhhc3Vq/T2LAouKtpc77nUfv3i4bGoCWkzKz
2fcnIeUnAXBcSbcclhWymPUdcSTiJ/rzAzIuJCZO3kdJYvyCvGzyzbMJJT6RuHca9l+fOOR2Uusg
mBtzmKlhT5CagbfeRmjb9rnM1hEHyrhlvvxmgetFBr9LElfeD/Je8glAwstF7YxwXr0pspLPalCu
ThsaM2zP1MBOtBeWtM7NhKIY/ZxBFKQ4grO20wOq5C/ClhZzVwXM9wqubgEKpHmOszR1Ht8TITrJ
zJYaVOxrKnbllN924cZhrz7b/jjvPRZTNpW4xffcS0WtxRkah2tO32h5AyGyfN2Cft/fAzuwIeW5
cQWEWZii08b43TMowpmqXzsbJO0S/TjTPVST1RD2xu2PLpPhRw9zgehGJcpfxwBSRoW33oKksq10
j40S8tg7WX6HHd6n5KynzxBs0Q3DJUgGDRl7QvAWEqHEXCrBaIGk+D1RS4bHfmLNzuXscdsf6Krl
zDJg4H/DF6Zg8+dEUgU1GUfK9QVHPWQO/b+vi0fnE6zayt+mgAN3eg5300kK0d7N4bV6c52YR0tX
+5tu3859L6oBKun5n4XXrU0h78UjkO/q3OBMRmDSKH2+UXAqlP5wb0t64S6l9I6LGUVj7EZiYk64
3rXxidrNeQIoZY2cLJbRRNW4yTPQCyMNd2Zej/GcatC2+kc0sRaYDw3ISoYFUfQCZbD09Ezp7kG2
2gWRXyiI0wtRqyjb+0UKL0r1KKu0k8EN7rYCySISmC+zGCyWr8fWY7+/PG/MUQK+21/9pFczKL1/
Kd22LneTSsu22NL6f2z5GHO4UeP0cKFur+a4+fB+PQHv4TjKlfBaNylJrSjSaY4yFEe9ip8kqluT
lc7jgSI0+/lJDvBOHnE8WBR1Fa6NQ83LWh5fNVay9iNrUXY/GqSKhN0yKkDLzF0kE0az+k8deUnh
W3X74NTJDw6RVhKdBZF42G2yZRLXdXJCgo4dg7GeI28yWw9E2Hu32O8u9u8D93IIID24qmaJ+yZG
a+UYGjGLa35EZkzzqM/wv7bhBQ1u7mPs7DwAEG3D6Q7YBObEunRcQ0NyUS+3bUO4uU0u8pZanyM1
bi0xbIzbB9PPd5IB+WFrDXS1rvCyHpFizbhfFjF8vvMaTXdt2fw05ti+b5eGEWNLVbi+QKbMKYDv
egb45vyCl1dM0PJtxkVhtIbg328hg/2QirpO8Z2ClicNyCtiBfNAHuCoad52qUWCLeFz5ivsS4bZ
MMGm7qiGRWQJMUVWu7H5W24LzM4bmy1AHytgXJ+x/Y2towOXtp9Gw8cg0LlpoxJqBidc/ASlYmn6
0UfOj5v84c2JJ+AL/fuAh2+iCmcZM/c44ai/CbylGw7auxWwV1GLmiL9Ng2zGyIVE7XTghJMpDEm
0zfZVIsmX4+6JGB3qk/zC0FQ3QRwEtwuWxwePPypNFwIrZVDEPaJd1hFIroOlV90bsppXOFqqGN3
1cbxdF760NB52IHM/BvX1iHLDD+XmxbOGBrL1RhGc4J9YAKmQlwc+mZBilXx98byH69RBkfWXSL3
SglDr2Y9zzQ4B0OEez+4+jNFw8BdLw7VU0pep5GdvgpTdpb92qO/gsxncHs01FajCxQVRBsBFHzD
ndekYJA5zfUEV+Ob0YP+STw7UIWUr7gDRzeT/u3lT1lJYp2eEpRFSCdGceKFi96K6vOBr6Twqcvd
DajCiReMpjyRbiOS9BAOTrAP3ypVa0Eon2wXvy9Ju8NarKHD218WNQNWh2OvhPv27NmVpC/j/qLO
KoUFzsqmLVLdggv5pj/5gAUSiQ8Kc/RxvHL9Rq+XEsq9hGjJTHAnwxYdQhsXVQCcg2Pdvv6t2/rj
dwwenlJL8cMPqZyLJ/JIs54Yatb23pqJUbTkWBMwZJG8cZUTUyuO4rmazo+vNRc2OG9/kWToh1H0
95eG/U/msJ5PX882lyPStyD0JHCT2DcAw+r6OQO2VT0BplUmPu58j/zlX6SVlUlwTQ/LU3MUvYXF
VXoP5s5GmWZ43PWDl2IdLXefEpfG7nkZaTkr6QHaFnpCGUrppXzj1wzKKo+rH6R0klN9zK8mBZe2
ttgXJcFY02esqBvt+hWI0NrB+9gA4Z2mFtDg/yANeW7RTGn4hulm1nsDvucWN8Vh+AATXX1/3T+2
D2yJRYh/GXFBCT1yA7+OUeOG0hAJoN6XhwP68922JdL3R2ZS6V78ia9SWOsCcnjmPp2SUbGQWBPD
V+IlKqvizwJfpbHhRY0fPrdPokpqL2pGv6LK8gQnQraH8M1iYUCmykWK1/WShlwPoWEamjwRibbY
NI5KvIZ1ZHX2rDpsa1rsiN51o3qmGI1kf7Pq51Pp0LvGRVx8dHlHfJ/j25LItEKiHTsUq3pMuzfF
flVXyYEmbA3UQIOOjDgtxb3g7s8QrQdeIEhVvAjGf9PWyEanQ8WDZXpa7osxJYRzbfiigSII/Yry
pGrHebR3hV354s+Q0Ua0jYB0P9ahbOaxZ6NT4X41R1QxohPOGkNvjezUjCCtCj6eWu0NG71ek+mR
AEH1m5zhw1vpC/NOm9FJ6e2Jyr2a+XFZAHnENauJTfzHMq+41NLDPXnHMei0/uol6Hj4rZsIdPfs
sSFm2In4SR4uUSVq3TKSdNs+3MBxtj+0vgEr9WQZ/sBn6OfPVLd1g3xbD04Y/BCkkx8uw3gApsG+
9Ti4w3xGSkWTP2gelVq3wzohGWmjPrSwtHcj+lqr/ohn/M4KmIEQeDHejHFo0GVYcmsw8jf4XE40
FjaaRTm6Mr1xMpUSRSHoNMkIyY3rTYFqzKWrC3/HGpEDfrQfv9kk5Z0icoGkEcmI+ohqPXsByFVh
uesAjklIRWaTc/W0EePK8MBp7lEPLNicgvaPndtv53yObjDEs8giAibc/NCRECmLGfN9pl43+niI
vSjIUZZIDR2zhbXbl+4Xi60wltKT5leMcgylLafm5xW3JPBAEsJrxjfEhjzUaSZgH0SrL57/f8T/
hsVBiOJSSqns1GtG/4OS3XCXtu1Nx3EuPpvOoLQSBtPQCzUARfR9Eet+lVOIoED6wCXvUNHM/oQo
5Ol71Y+3P60YMhC9kO2BdHSRnIkmEPi+/jbWSGtN+IkR1giaehYVzeXmPEUq3ekwMbrIpv2P61VB
Ym3TJ3XFBBJZr74qiDy8O+RRNFvaR2DhunGUcMNHTj3aBsrfqOkAoUCicJUGpxOddlTU9Ay8LgJU
nT6AnlGxe5qqh+7OZcsLabBhL41Qa6VWi9K3j5ceNt7qV/jkg5SZ+RP3vf0buztuOrOYi/Yvl7CC
MkqCg+yXmQX54EhJu0rhGheitRoZuvACRwdXAUPdMbZ/xc7BxP5fa/ecDBRcpusR+9ZTfU5OYCKo
iatE9jIovdH8SAvWiz8o2kBpQxkBzxKAUWrcurspvexwNCi1ATYRS+wmVYCIHySkP7W04+zT1Frg
xgFW8A06txU0abBOE8sveKnQ5VD/zLjpY4uIMVIr991HIJFiMV1rZEQ4zZUcx25Opw/8ICDC8aur
SvLJjDtbvPxg+BNxOlTMBHX1wn6a6OBG2bcX5hCdGSl2ni1c0Szq7Do7Suvp2v82lK0VIHtC67Oe
PeNdPMsyPx0bwlnhm3Pzn5uRHEQJSxfsjIcuBQJUrXtXWNzEfqWQIegF54lGcpYsFC0S5mYnVlwm
D+WcZP1dMQ6LiXelQs6MBshXzM0KwcnITyAprzk4i4MwuzPsNcpYzubhH9/SWIZQvt3bc5/g32Ls
oeR6SoOAA9mOsPX8dX0Q0t/JQMI9tSjbtR4dZjzPtaWH3nrGDeXbyE+WWkEA60ogbhz951ApPiCQ
vF5CKFqbkLVlH3OTAAiKOCnawukbitwmI3aEKc9oiWJtL2Wp1lcgkU4zOA0hYsyirbzZRyLOVQ8Z
hZTWXdGxvCILK2g20TAB/Z9p0pg2J2pOyGOzP94jAAVeFChuBLZAajsdS/zk0tESIduz0ZuIwwu2
CdRJJFSy7bdTsHYIFqgIZVBNVJqpGIox2YAuHgPC+iO35iutHClrCo5ty26kCDgBYjgEuKjHZwpA
tKeMdbqJOif/Tsvdwc5vfjGzpXoRYyVcSLNR/1M+fcrlEKXoIkpO4j5szpffpAF1p0NxuoLOxI3T
HXi5yH7Ch03UV4D1BTCWLI8msv39yFbemoorFQTmhVvQ50OE1mYIJqfw+m9ibA16gaC71vY5/Z0O
sILG9LEWrTKqolRc+s3Otl2crgZmKksUtlnT7KsyVUTNc+gGAUFV7xKzcieDByM2zEYFAvhtDf5s
R/cqhAz1zJvxALxMEEdFd1x11FCK1vfmsEIsNl45mrdao7aBPZq4+3BVcS9iNRBZ4TCC3BfDYJYq
gsGlARk0t7p4PC2axF3iQE6QcW1JLpZlAy6/nEFCbaYoY5l/ENp8FbnIWIArstHj1394645RbrNS
ZfgHEqkVMed0hTt6iNmPyPxvl81GNyEpikxG/FYGGTidkqBkFsHjdDfKvPdKcqLnOr/2y6NOGpwq
40U0zZFWhjg7qO5gETk+15rrVTWCtsqYcxR3lam9g0P4BvMWnCdDWZoKjyo8sEVH5+46UXdgSToX
pYSKtVd02RS/cmHZH8OOpMbsy7D0o1c4bl6tsb58XQfowku6gJJCcmAUSz+gzKA/sb5oiiuYBruh
YUnIRqcWnSyyY0uUHt9FmWAJGw0HHwCFg2uM+hPhkULFqc4Q61JxOis2o3YrDh0ksNXwtIFz0p4s
ep2eXcgyqZABqN7nrzb/MYAP3nzKIk0CRRXAfpQGBKc4HcLGLm21DFNgK3HpYuOiYRJS2Y8RnAkF
KjpQ1ucnZHDn/Cn572EWooLpS0l4k8iuKGGMX7KOoTZUoAfpL9lRumVHAMpvf9bCf0U7EZFSSnBu
X9HzzszqKMcY7Mw1DrOTyykMqWmGUTk/FxmWkO87bgGSLyX+1pdzcYACDy6mtP6B1w5PQcdHDZK/
eskctbjmPtKjNPECAD3gAU3t4ov/vx6UoYZ3+Ny08Jn0ClLK7u42hmSMdgbUsbLOrByS/zrBiGJy
DiAMvFmcCG4DwGmJ7O8pU09ncikSZdmSPjuV2UJJbtYZQOLCd4zduBLihkLHyAgA72pqhFSFeBla
wFJ2vqzLHMScffjgwhTIpjoz4FskqQ6zsDgHmdO2vbJkL9S5qoxjckhD9030katnViNocvv8ndHY
0ngaYi22xRW6fxSAkVpjLAlTajXG8Wz/zg+RsKV4yoLgXLw1E1+/ky5Tgaczxak2dxFNj6EAhUKb
z4xcxCnDsh/pDzJcHrFe1ql4myRNQkRo20xzmYh/GEdEasFqpiXbwooYhT8OXz37zB2jpbhWZdt3
71xuEEjgDIfAVPATf+5ZZNRcSIQZGpRV3jmnkyqCaN0sHPh3vxAS/chrtSY+25Sq5milzZ6sND3a
h25MCoVvMYmhBGGMD8/ogscn+gAQ0sw7JAGi0lr3F+ie0gSHAC5FfOJANuK+QLok6GYeo+Xs2f6A
arg/zeU4JsDyRCvTfqev9t4MtXVlpd9I4IbUcohsS+STJEKJMtx2/2wdFIsspSa+4ayMUWpMkbFT
RcakfQwGZhWeXALLiOJz+PagvFLKw6SgB56fAhFMAaldknQUE6DjXlVs++p1EL2tllyCcWY2Y5gL
Mrgd8Lr+J5yS1isqc3l11gs9iNqPaBpRLtuUkBlw7G6IIxojWRN9pCLPiYJmsLiMqNUCLKiBfiGJ
4lbPHXp4JbPJNfawhDAhBPkPGcCjumVV4jDiz1ERw5uyO8Y/I1ZCRIL0ECrqDAYbVkp87t6CutEM
PrcxpOLMqzxO5bgz4tU+gXmk9E/szI3GKpA+pe+0uRTFZTgHQXc0+PDPrB0eBxNcCviorpI0N0Z6
NbZR8XhbivhDUGlpnGXyxiWAPr69H9XICteMRf1DfogeAIxVJEdXKTm41fYX47ylfuNT+c//MGae
m/NYMI2uVn+wf6gE++9e/9sEcYYEL1u4vnZJZPzJo6bH3519O9qebOTWT54xbtAyCrDVA5hFfjWr
BSKN0xaSlws0SnbvJgN9Q8sw3P5nWVqegGmBd5QjASVCMpKzvzwgaWy322lPQ2yVokInmvv5DFrK
pmWufX49odEkIDcUYg64PFQRBFZHIgxn3FOGBFTO03RD2Ho1xt2uZ3iEhNF9gvw2IrVcUSuoObCC
0njuF8R3UENXmZUIhGZPK4MVH2UEpGGHodJEJAI8s0ZaoQHqs6sN2yxIM2h/FqwhPspkgrA/qK5u
6+4vKnR8uBWBlzPVI9t/y4R1/cv7EfNclRPoecjFuBpJt728RGf3ndQWqYUCRP+RuZkczCcJ6CyI
NCyYCxz35Q7iMeuXzk4kT0adQ4AF1a+RKjs2UHJs7ZYw2wvaaorgDjM9MIRCfQyNeFnvI0yN332V
azyMfthbhMIyukZOsNtWawdkTBbBY48yt0nqjrLejCr+kwo17W0Cpjyzuq1fA0++vjwWcBAS1Mje
du6wh6OLVboX+ttGp4Df4fJLw7WALLU0GvX2myII+JRT4ZNqoF9ASUptVLHtNLn3Tnyi2Zly8nup
dePLHNP8nq428D+PmwPBgTMdy+fPC+Gr7Wu45z2aU/M2GPCOklGR1PVb+gboDIbjvLokJAdwjgWf
16qalLlqnX5x4wQLQ8U44BNCuZ6d/OA8Lcr8WKR2qORS6Qv9R6QwyjV3DtC2rdHxeo2s78ns9l3T
NwTUgfLU+bfg+mlvKqtW0pEH+mqiNLIw9ZZQshAVnCSKzYJ2i1lK96pfjL99JbAkYwofr8rQjFdK
PA8/75lTjM6hZbZgtB5Urb2Mb/0+5FKcBoAF147SAEEYJHGAhVHtm4sdwmyz6d2q0CoaKPztB8nH
o7XGY2+0nFMEUN3IFg1YvRaZE0TS0tem/AKwwWkJvgzOxQlqJhlEpA+FNjz3+jgdASXgz8AJ4z7g
ZKeuByzCZztHCx2gnTAcb/iCezLoforq/5r38Fx7DaySy5+Oxzp+uiFhjLSQFquNAoXCxCpn5+Qz
4l8oCDcCVsuVydzUOqqbPpZWkOclVb95KuevBTtbqUJQf3KZyg+j/0hQ9YzeTHQOOKDFAdtmVwE+
p9QWQh0u6WBgibDmXpaLmXZO6yNME8ST+JD3OVURxVGAIaF4ZL84J6PnsMpsDiEu8gbrWAhmc0/w
PRWkgML/6rWyk/FpWEROIst0H8x4VaqAVaT0N9CnKuBepqjvi/WVp7o71KFCZZW/N8Ta3UOSGdjc
Tdiacouc5DZM4IobirxXKBW2HtIOTiOzvNANSXvy3RS3EdHriC9mZSZVz1da6rhx77pdLqBf83cF
gxJyxC+HiN3SlFLz2SBJJnLMKDd0ftmLJrN6/C3dZPN/ZbDT8BHDcG53AjJXIpMKx2VFxmw0aagi
tVYiEh8lDScXB+GQuaW0OALbJ4e6fFxd2d1tpf9St2UQrDJKtMtuo2p8WdKNTajdaUYTtUW8Ec0c
ZEEHXtKXWKdgDpFdhYp1n04JIsoRREWH3/8wCNrLkwWL2KPbBONwiyvUil5c3byJq5ZxPQUf4ymR
/yzKM/v7XZAqPrX1zrkw4y1n2CoWYw4GYntJf8QH5c6vQsbRJrW4HjY0bdpfveTgr9lS4S0jUVsg
I0kbxUWywpxVufkiK6vGq3NdGZfWKsP40IuVjVbtJ6hy498nt06t2pTKjhNDxqzM68i6Ak3XrVDr
uHL8QU4Zv6ADzs60D4DU0uRmDWst8vQ8/81/2J0t2HPbN04hYmvvHfkTex1rRVhT0ZvlDqUob7iW
udpoq0+St5pLvsvcVWXbTydNE67uOHI3t8Y0lp3GiFm+XEOnQP3w69yM2+YkQ6z2Mvgc2KlVXpsT
1fNf3s0LbvKeTPfpOknW2H8ydDky3XbUsEgGfsxBrgQ3tI3tsgDzlULoNU3sJ/Z+fPvo/DFs1KAE
DRVNKxTTXd8R/xtfc2+AOzBiQ1xnQKMfkE1qsL/yIeI8dWfDk6asLfQ/XY1YOl4Vt35F3U96o3c6
U63IOqnjc8NqzEc55gaV8OokDSO8OTsUU5y3EbkxYIGJVpA8NgVKqHWsZcSOEk2ehK4cP165PKyb
vPnBlqlLCaxUk/zVEiwJTzoaW+mFATbT3JNiZb6K+dWAnT8NJlwa3yVRu8XkSEcY4tgD0ydHGE3A
jxCdFGKnunFy891AJdrBotQFk1KaGH2fDc2t+2LBBxN2UcIAJaBkI7OrF6nAdmO0HXIzsPElMWmC
iOS/CFEquxAx91FjEfEWcfDz7JlCXbRXobhn4uYevZ6tvGEbHzS1Ij0Zb/rT/pDMDDt/HFnwKAzw
jel+xoKUCGKxHZB6ZNqRuoRcDWK7aVT5ARZOYFd+6A0ZRnCjQdm5HuKvVljBr1jAn9LwmuT42PSf
4RRiu9KJl0+yNKTd8EjEFA0kLE8nmTHxTYgmZfMhgyQZD4I+HsZnqStauqrPY3hFI8xFrxT25ymR
ux7lSjqPaWCcCPywQW/zojXeAzaZyJrPk5NTdAWd7ajXIeauTB4mQBvY9CC71eeEiJxe/TprGEDi
fk9BPpJlBon6/ZPLBMHU79xpILG1tGANtHNcZqi14e5903+5zgu5QDtKn+yz2/ocD9yBAbqoawnE
pAXMyJLvwIQ7h1Sz86YcQxUQV2eNpgVtGmL1yh6wpO54ocsXiCs1LxO5uvWcobHpSmroivlvkvHm
9tyG3Va6/iSk+rP6RtklqR1vgKrJiq+gXnikSWmc6Dr8Ph0nUgO6W7Ivm9aje/+ZS5LykTTAa1yh
P2W+mgcs2iIoRpt00zpdozaqboInovvwoZ74nKlVdgLbnYbmcyrqMc2ESV9Vmh06QuQWkWnOqPW8
mYhcGp4S/k9ydvT3HXDknLqQO+9fjVD5x/C+ulgkz3xSgKe31JOv8F2l6lwXjOhnHbaH7/4DY/nJ
hDz0w81LzKj9FF6Ik+qOeC6cE2RSPyRjQKn1NWXFsylWxmWKTXnuVMjdI+x3vdbpJZ+IIYw80+Bz
9psPWZ6fIa6FV+uyo7ogY9j6zZIG+J24GfTdq3wW0e1GUOlEBOxxmjp/dwysKrtplD/zAvwp8ul7
++Pk2WnryJ3xEKtBDk++g6u0ipAv/Wq4TR4INaJSBemForKcP3Hdr5+FGPOTB5wtsI2OA4iczjcE
ZfzO71zCtYOC+e/FTeXQECA25Ds0OgX7++NtxSvyQJO0LqNfzp6mIYpYMVUeG5T4gAFE2dU8YggN
9+MvdW4H1Z/rUIGP/GmRLngVnuHsv7fLKoIPnx8Vn+0AonzEoe7U8BxiALbHZbF8ybuOosBZRmG5
euKbOeREPNrmCr+zSCebDvhS18IVhM7GLUV09EB+MeYdxdymP5fBir91vrh+0/PV/1RAVdvxFsua
1wsOpANUJYeaiLiwIaiKdDsF9T9EoilygvpGvVPnV4Be4ZaaCbgp6Ob4aHwJRZItG1kBu3hZvQdz
FobTCONw7It/xUgB5Q1KV3uhv2RJba+36C97dCO0KTz/7B2q0MIgYcNqVmGD5WUWag168lIqtigM
e5w8Rt6auiKrKb3DrS2J1NDLE34s0PjQtOEkuE4KcX4AUJrs1/u/JWL4JaqeCOCGn84bQ0hLldAd
RuJyFprJsDURdDYVdc7JFI+noTOXpKmu6/wxfZCQpmqriPY67VcmzeeT5VEHbzOOf/IjndQmK2ZV
xuihZoajKhKMM8OEZiKlVHjyQHYP3t2l8VAAlr5eORC7aC7+gsnygCIvXYBWrhVr0gwM9MB+agel
HLIp6NGLJtQwOGgyXYFVKvexsdh142+DJlxOReTf2j81U0iBZ40W5cD3dBlZDpBd3mKdSd0zOJQA
2fM95lnJ7a5i5xKMcQqDvLwhEteD2t3838LBE+bBIDsnBAbfvEDyE9L0guzQPb5Xx99TIQwpOq41
MjpaAwPnbrj8OGv8ED574vNLfVR5UImpc0kFsHbOJGRj8qJzc6EbeJX85o0sxxbbR6wArtvCjH5c
RMOD9iw0DnaeSxOEURkshzer1BdyLkb79OE9YYi7E51wTWZowGMXhwWX5vCS4nJ2HSRoyyE6LKmh
N62AZbqzFfRRNuBmYKMD3/xkI2mK6URSymmNJxeDCKCq6wiSCOtyE7OjnoBBqovpRQinb8MeKZfT
Sst9uXmQbcuYjIbfGvZedrlb6oQTrFxWo9d9+O411lsw3NAhw2ArPFwNF/FWd4tcNmWt7jXhxHp/
omRVI87x64UfB7dNZ4MQPVTtmF8dbC/7a3xdoDX1yXknQb1ByZuRSxshxOXCdZO0jH0jePLel/3V
VOAcsiNu2Ynj2pIRpe/NeSdbK6UQIuWyjn4FucnpLEEC3go5ou6XJVWOhdPim1h65o62nS66ap4C
Tqi84BJcy2GZ+evkxOxM2xX/8z+4pMa2MDrurdzQXRN7P0ekUwqIzurnqY1iVLz6/+U7xao9qe0U
eIRmgYmBwFqMMNGawo5rcvUZkbCp7Qwf91BZM0aitogyN7UBSHp319rj82sgVXZWCs0VgIpZwq+3
7AYhHRZdyw53GMVBP0i1/hxpW59y04+b4+7LNCBkWosqZGQ5KTjL3+hfXzDCLnFWWCGR3d1Nz1WZ
RdjTG3fNSsKMTjhfk70P6ljcco0wqubPqVNAsUXq0vpZg0lB3DDRpq+Kpw7b2QRX8m6E4mFXAb+A
K58B9hxOS28hsDmK3njApQrQ4kgXLHgyhuCXCnRh3jZR0m7JH3/wS24ep+EOlt/BW2qCMHthlqkt
P6LqY5IrQYWROXRTvsz7mfyv6rR/KpBRpuqNSa9+8htpFKhtGVls0uPhRawslACaTpKJyCOPwKz1
88fDaOmcZJiZuDgVd0JG6tGyXdnzA7QWL7C1qmb7Rwod0YuV3mMaX7AOcqPXkJLkpejGh9aPxcoV
t7nGlJwedoXB3Vxz9j7ecGgQJ8nyTfIPfUK6lOFAXBm+KPJ1soPVBAnResUU8KNvuIewWtkNZ/Fm
8fT1LobBEldTNFmoedGExMfRF2TEuEMGoupfcQVyBud073q5FNtg3yYpuLldRBLGHId2L6/zRtJ7
6DyhulgoUaca/QZ4lSr6vx2XKeQCSJn2XHgQ/lz57Xyk8RaUkVg09Ow70nwa8rJYqdR2JKXAyV6V
7bf+x/Oj8Q6SajQeZG+xfZX9ek6twPCAl+gZfxV7K8iTqgAvjw5e9khhwyl2rN0ztpcjQEzsd2l5
z08NQElTNS6ZJGxU48NYz56SyDCS7098aWM/BxLo6kZzi/rdDozbx7+svw4kWV37NJgLqy2H4GjM
Wg4UPypqShI6ShzhJHrxQC2LdXw/rHdMAYH9tPucI0gxF/OrfLbU0ld27LNc5iEtyrEjrKJZs4T6
AJziO/bpOFcqMQKX5y21+zBia12TZ3OW9oVSq5Qxu0ydQ/oskKf/4WhAhWwgwjdCdjCP5ObdMgKv
8xCFyWyG5SlFgZjEBgxb44LcZ9J0M4sON38Stv1MrI297H3CQWsaHwwe1kXf4Gd/UNDBPx9ll+vc
jg4VXIJHmtkA92Pi/EinMz140LWt+2iqq4g37f9dYRYVnL47vRvfhgvC8Cy03zKB1+okPwLFDhru
Gx8AJMJCedEDAzxYVnjj9nJnjJ9cA6iipZ65pSTTt3fqTF8HPEpJzQZ4GXwpaF9PFeDhPQ4t3vv7
2c6X7cLTIVg4jccojxNXe6mWaXnJqxV6DoeVS8Sma7FU5JvsZfKK7fwO+KRxN756WePIqLxXYFlq
mkIsyE1ZL/Reh33Quw5C6ViZXiILs0p58qT5IHYUobHzVOCas+nVI2AktfbLKyPmVJRTzKnIHCp+
sn+vsMZhRyTR54ryk7Hctp/Ccn/hxTLs8gGL+95cJg9zLUJP+pdW/PzG5dGN6vYrVvRYph09hj2L
Ll/EVMa5ZdWNdZG18UIYLmaaghxXNtSLpd4P17FXj415NFXSRjIeer2eUDB62t2G4W3vWoKmwlVy
3mxenlmCWiCEoAUHPjt1QuXHCeILxH2KMzy9FmODtMiUITjg/zzvDqT8Wmqtiwdy1fpTByM+Rqzd
PcZaFv1Uf+yzdKPVISPvBG0hVdackTydsbalAR93YB0QlPWZQa3uTtARSFGy2hwOhKmMN7UO/Lc5
YKivHlwRmT84o+P1Ssr6Mcl/apDfkERU3YAkMYJuVSQC/lO18KLr3zInVKM39ddoWdlamP2fLp+i
U8ZYFNDAYwo1w7IKEG4+mw/2n1eb1+YeRAsisoa20Lg1RcgLMrzEFmjXwVHCwZOJSNkVTBGT6Dne
ZTtS0FyBIB+aaGAVuWVRlU3lnWV2H0IPFUUtlB1W2nNMZBQvfuoeRxYV2Ycm0xjqmapSW45AdYwl
1w3IAAbUznMp3BnIC7yEVKQ7ophm6REJftimPvuVSBBqsCH9jtARoVFNrWGk9nNJxMSG6l6F/VNR
lg7vD1zWrMuSw37XnaGwoH9U1L1WN/Hvh2VEkm4rDfF/0jviolI6IY/AsPQZ4lrWmwsKHp6SLhhL
PK00vWgIuQPC0KrmnO6qm9w1ZeXl2PNiNb6ZWUWGwolaDpq15WOwxjKu3B23ris42Gv7OP/4tTFs
zcoTYQCLjsbimp5bSbGZ3ZAvmqfhHzgvs1qT+/u6V7elSwQBtxdoRqNJCxr6+mERYtMji27FskbJ
9HjfAVjqthtwhlgHRfR1L8d+R+cMntmzhCmg14fzuQ/WKTkcBZQxsYNx0xHgFkqIUVCE3d1AL/Wf
rgPXBbIXQcedxob3VgUshbqy3wFxfxG2Sx/GtnY/drPnOAZO3dc3SVMheVDPzRXEEQvzxziZExpE
AOzhBJTNYhvEqWXDS285i0ozQHA9CuYLP0dYIh1vZbm8OHHCV14qB8eTgwWRlU6JgRtUU7qeS7+d
T7qhrVK89k4Y8ZQDXOUUd+kVBrXuA0uomt6GqS/NrIIhKwZHkj/WodFi6lIUfw8oQ4lwU+jjoZt0
7JPZOK7PDDvglD+eHkcNMZC3eCK8xKy73giJOEpJXCTmnpx/J9q2ZNQSYnmKDPUFNH3SaYYazstM
O1x1VF9jHxX0zvxNTKexPKN4r/DMkdpHn2kUYvVyPGBc73Izzy7AmrVoV4gEFsp1ERr5wy/cTpQO
WJhkZdRYXGwV79a6sknRNU3HXoTQ4yYQmFwumh1DybmJcwh1MAS0PEUuPAow/OrmkY1yVxSuyRwo
QedT9+/1hSX3mbQ/WxlkgyKeXLx5/9mnqg3Ns0nXWUhX377pLFpShXG0TMT/4eY+te2nmbdQq+xR
tWkgGHvB6JhKWJoSAFL1kAt2AX3W6MhBaV3c4uI8xA2d2flCev2h5nUoqJ1PrhkFCeyFxkZe8oM/
XK22kZ2RpoWllj13gNfRbjeAaVPTQkSmyJesO4ZH/+u0UsOA3bpi8X3lqwF8a5F7CJCCRP+uh9Ff
ZG8cLumpOCWRZi7bKIRPR+wm6mMoP9EiDakDKvObRBWkWBy6E9y5y3zW9YHJ+NmMnqSUuMrcLKff
HlK0MtqZ5BmANR2Z6DXA2nJ+9Gqkx8Nb2DGholwJiSD2SZyRvrm0DZjPoybofMlfSi/sWlG5p1l/
f/BHhe1r9pF6ziOfYFM05u9/MOflsmNIXT7Reo6Dj2PQ7jEo2KNAjGhf2IH4qsEWdG0CZ8ePGO97
LaXHwAxZ57FwqZ5fbScbUnmyjhYT8wpgeR4C8cprUwXA0HxojeUFh8cAy0j+CzIsZ1vbk6Qu7WnB
3h/aD67LHMbAZIEN479hH/5Zbk0VaSz+WLh+jwixFtLtM4ojpLKwxF3K2ZhiJEJvuytv8rl2bnWl
67zUshkUWsfK7FiSKHXfv3mERRv1/pWyv0aRcBLuDP7CEwpU4GqnMSWNQ/exbgVfzFN0Ifj37/B9
hqeYyXiF7cqz1jH08SjZu0u0DiSQnYZ9phGsFE/L/Y6L4VeTq71nAvItDUXZyP/0XL5o2v1Xid/x
30VojrpD7gw/W6SOwlrwYCPNsLKBBq+tjIhXa+qvtLK+mAP5a8n8PPTB+hE+LyxEs0rFRvlLooj4
3M7XB/bgT3hzIMYNLAM6XYrkoydvqU1B/Vq3FY0egicscDZliZv7VubSANXGk8di8Fc/uK/K9mWA
tVRuSPzDeTkdERRfZbOXcE6Ifcydn6R9uekcXYGlYxPW3OjEgxX9GqWh+SvHzOYf+BH4Ea1+Yc9o
s6groFo7Pq2QGCajmAnayqEzlPBsZf+wuHBanIxQtGwB9djo5YHhxCZve7tB5iM1DB/FV3EDPnw+
M7sFABmocvIFjUY/F4W6pojJrfqL2XlWwtwjjJgX6FiyvJFJpsZbgZHVcd31/MDVItVxbZeVu/iI
wr61j8u5MMOyMHwBloCXopz4E7rNn/7ccnwgtbRHhpk39KOEzrqdN4CLA2HDSeXMf+1OYHIjZj9L
a43tx6s3z3jTY6Mx+QO9heJ0E1ljgHnvnPuqiti9SMp+ZYD2jwlCVsYYv6m4qwRS3DY1Ah1ImDye
8TwkBBbxRzyosix2InqFwcb3zIoJNWROqFNX8Hw32ip0IduYkCFup+EAB4CXMMJ//ppQgnCTbmvI
MtBT6zg52kzOn9VzRRl639dF0VJMD2Bl3dru8NhdvIxSTzspeKo5VXOkBn6xHDbKKKE5hsvTDlK+
Jx0cLGrPClvEZs6tEQ6t7hyQqBGtEQugi45sHz/rz9uTsvXkYdompK3KMRBI3aIxbJ9/STir7Hcq
OwzFPkywH+pUcqkXA/POG4LuWCqaJT5NGmfL0d7BAv6JIKP8D5EvDT8561RoVsqkF8VZ014wy91P
GvvO/CjxY4DcdOPVjarYNDv3a8H8ErERnl7dtXhc3lqp+9llaB53wt6yQdxLozxjiSzHlBjb/Mhb
j9Ydj7HzjbzkIppRY1bZoHz9NW7OfVT9gOkDBeaZQdXcNpFKcvSd1RqEaOWBTMIiKkHhRcQWT0gS
3F7tQ66eMLD7YGMx4zcJyNuQPVyWNAKc0xC8FfzUpwezFnyJ2ls7rsxSLqgY61FTy8nv9jdOlK7V
jQ1La0wq+IQ2MVFXSqprU4yvAm1QfFrbqiz6v/49bsxYXZbsn/vK0ftUK6n9Z4pVyapnC/xt8KkF
4uOgpdV6bNpBDEOypUMx3jx1eal6R2A4oJx0rY6wdWguwHOGa9lw/sigywsCnMSQREho/iq4eQNN
/t3dNRQh9e/t/Ihse8JOo4NrUsQOeu4GKE7NzWZ2fxbHJimdUVJWn0Lp7E1YQyvLYaC43LhLPAHh
wWTj2y5Nc/Zz2cOK1L9193ouO3U629rucEzJXDLvX0iheuEuUvQgKLWYp6LlPAFXDYb8NLLAncTt
UVhz1lWVGCh5jARKcldNzteGUuCa64f7L5UCKbsDR3I+/soDummBVv12GqmmaUXmw8pYkfND0eJi
cO/oAQXVy5YXhb0kZy+PR7aomhj87Lf3WCO/6XHYH/oOhQKRdTdDGujRvtluuf/zU5ixdCjjs/Nw
0fJu6CDmmBVW8cosT4g9/s/CuPBoJLrbI7TFTfthAUQzKTLmv2mLofoBdKVN4NtDduIREMHQLxHP
76+91CqisXsLDfPGUWW+aInAjQVmYLQ1bQ2NV5rGJPdQTpiuAuF/BGECCZG16rBIrAnZkfUkfsld
MhHkGZ59swM6DqyQMnrYV2gGFm7p8DkRICbDUEO/+OSi3J8SSpYNH3Wfi60l/VM60pibLtKw3CJc
gECXeSUoG8l7a+lcYk0zBAFEo4LQZTZ14/MUZh4mhOzHOFCCAJOTQmHPWZZhZsrvjtZQr3sBMUih
XVyZiHxDLexPu8xSZbdT3iCjdFZAwBMhDnhSyEPKRE81klYV6DaN4yXtGevVocAALgHD0S7L8OLu
ixuYlitb2lhIIFWQ1QHl+daIU6dCAaBBrY53PkvBOdMq/Ig0GLiFwVY8bHo7fQhRlcakBOe8POYP
5i8IYtT3j6u3bB4ifkHPQFqIZV64/9vi83caby/qVy8SiUkoeZNnfpbHPkoVNRnUtNkDFm5GNNQS
AWspD+cSeK4G9nSa8q0DHE6A7dAgZA8g2WoGRp1LIRB6BSVaZT22oFjd+K0ly8TlYkb9CjEBH4nx
mVmFmYMKDudvbVWceWBTm81HsAIgpfDzsMvOcFKX6gOu5MTbfWq1IxyIVaRNdb8HgsQAmdR/LcM7
ls2RHIB11Mc5KU+9af7EMB/qgeITZ/x9Vpttm8ZjdL2iEWjjpZoL+YvTICRGAiny9ar/4ET47X/x
nYT4V/A6qrvw/oWQiHERPO0GfZzv7eBZHJqYk8TmZUAfS5pZNKMDSdAWBZ7r7PagwamXjENrA5kd
h5kDMcSmXJQIx1xi34boeaKJ/NKw00qoBIX3zuLG6wR9mvZYTYt3T+g7U3YQRpkswwSOll7ig2n9
4ZvQRg+Ldo5wqaj3PSN/UyS9mPmNu4vW5wjxl1Ph3nA7acz4OzZfX58bH3yBq/Ig1qmjOKxsXfIM
9VgWYKNd1Biuzc/ER/RMnfyexCxZssD7zlY5/B5DonTFfJ2eOH8qd+e+RwiRgYHz3POOFCqBtbB8
SGCNA+o4eBaBT3ITrSs9e0ADGlV0wNLJaQNNHapLET4eVIzYM/CpKJxRIbux7zgwR7JmgN8Sz+yl
nhQpZyBH72Vpc/YXJA5JNDUx72hcB36jNUZGfgYcfQuU84HuiRGgp6SwHgS3Kl4yX2X+6YhYbVkd
Pq1Y/lF/nDVYg8Sm0fSL0fAbUhc7Vu0cl8QiLM08KHsLxjqXi/8XVXAFQwDmcGlyuS5Xfg+kaBmX
izx9R1S5Bu+ksHf3vOG+EixdVWaqTG+M0+5ovo7bRb/+WjXOLDtk6KFsW30hrv84JtY48KhMdI+2
mmK+JpntiLAz47aiPokFbt8LWPZJ7aV6dx2oxLdkp/qRPuGGyrFlKfHsVEV5NDiD4NfHnk02t+gK
uedZwdisIBIhsL6J721V54yOi+fB1XyId3cIrBDkugmDjblpwy5RTbDUCNejwo0HdpqbmXv2OciK
sQhd/yPHOIR9GcA0Wfznio4+MFUGEUtnAqO+B4GnH3oP3OV2t6BpX+wwQbr/7LYTFcPqfG05Ykzw
y10g9dJEIt8LOB1K+l3+NDNgFfLdGwnnk45RX+8F4bZfGGGG3s3vFssh5Hg4UHnaT8Cv9lBF/2jH
/sPOrp7eDl+w6r0gKXZBlixaIMyd0WYdHFagSWZLWr++SSmh/HOKs6HX6kvOYSzFv2Ks8FeAbC3d
uO3B7SeyU36VGbVPSphVZFC0xGCxwJvJLfSAsGvZKCImgDbTz0NgzqY1OsILIzcDeLC7akodgIrg
lF2iHuJzBcfFpBAAFM2fXQStgUWqTe65j8/T20+dpUUxU8AeN5VmTtp80QYoYofw75B1XSopMrAl
aTB/C3f2zmHpp4UkMplawpQftx7fqDImgNEgbwRvHimPEbVVnLRdTY5JqnSBX/ktFBXgML/Dt0X0
ZFnT1E/lWUhF45g6VbJI3g467bSoup9hjFy0I+hj4KlgUa30/ozJKJSU+5b57vTYhjNtDSZ0+gEU
nK9Sx2xgXlmZvTp0YNzXLnkH0s4gEoGrEmZJD5/4H7qLxDn6vYghKU7rmVenJGjDW3OaK+MYIiKf
OBzdz+YeQcapriFKIus4n81UqoGlR+VMt0d0fCoGBP9lJizT3iLWs5RHPvuFV6Xccp7bQGfk2YjH
HKRZwbEFKtHLwvoZxGgZu/5HOQ/b+sw3nVnPN3hRkBaEwHyDiA9tbzOLhjx3oOHAfZsz+Ix9WDIF
4YnszxcV/KogG3Bk38DEvRT/rOIBRv0V6zl0D+zH4eRi7sJuz07w2+S8B1BtPL8bSFEtNik+cgD/
ewKH5ftsr0kd94hC8Afxs+wsY4QxV7tu5/K5mwQL9NQg4Sq24TGaz6QJxajSj37csDhi3e3z35Oc
cZEdvIoKA+KU8oROGSrVHESDRorp09kixapslx6uQ59bQ16SBzZUKLhSaR+eULzScXz58gr4ggfk
WvSuQTOuMnupJwDXcRA6xb56bRQp4MrDRK61VCT114k5dYYoN4XycSwx2L/o2BJfeTvB9b4XSKut
vcLtRFPF5S18Yy8vlGmEIvBDeM0JOrzvxK7ohzw0swXdmgp2re1gf35vadNRME2E9vyFt4V2Swsw
pViWZCOWaCWbA8oYLqgl7vMPEof/fHpZa6DiUfRLLMRD6PsUov4K3ZE5KiVnk+tKuONRokkFqmxr
I+7eH6id7PE7+F11fEMCL8C6vVVce0ihVAVV/vM9kThmoNQ0PxAvuo2yCiGp4bA2iXDXMYtXpLQF
QbdEHX8yoacpkZPbjMT5cldKRUmQBSu7XA8uCugf3ya8exWJvvLKEZjL6/iPUc7YsdsrgNi6V6Ta
ZeXorzws+bLc7tlb0t2s4YxYQIMFt9Gta9VfC9b08y5Y++JXC6NPVfAxQVmO02PKhL3/xcTTGt4S
ryh7X7U4Mjw6ovsrUNe5yh9OqRxApsQpmmuT6L/h9uGKeQRLKWTh4cYacfPTxpCkNEYXxXZ9V3Dh
fdfaSRlvG/vl9CgJCFNSzwglOqKn+k1RS8SYHsAMv/tQX4DTttNldaXo3PXzjtRay1SAx11sCuz6
ygfNNltyvmgG4OX6uYE6SFUK93g4CW80vdTazzDJSZavDSQZH/JtYVfOXx0Cr3LtCrB9ajgbN+75
Xp+OiwqLog9+iuZZNLSv+ehi4vIYeYAg/NkwYB/1BB5Vj+ao1fUh4DEo0zCpZ9B8nlb2Ru3KXR3+
EMK1cEsGG4nZ69dZCb0NAexXp2bGMdpup6mhVAv7+UHdyTfuOVGC1BYl4mg9QR1oc7Gcx7rFnMzU
YdYkXaJSioA9WR8JoElU56/aKcXvMkmDee/f90c3gwKsSPb10goLpBFLQ3acAqoX8YRVBzhKifsV
sfvolxYftaYPt04lY7WijI+GFMnI0RmK9bJLIz29b369v0Zl+tkcovJM7k9vx2Mw3viUxWO8q8d6
emy5o6o3TNZ2wXuBJyCTLEld33znHH8RmScvDjEcy0KTQuU63VCVrV3ep3BnsQglG7cZ6ggILxT4
x6nJDIQZnZxN1xtyViC0Otb8aCJiR9fh3ohzYx1gFnr7bzNyP1zj7r3o4YaeJcRSprMqiif6IkEG
YZqhxQsQ4lbHBaSnzlWxVlCqWI6o2q0WOTRZWOIM50745g1zd7hHo/+Q98m/p5Tc361Q2rnFAOvz
nBrFoNTJmharSx28d6Glo8jABxycKwFOm+TWV59z/uJC/ENrdw2Y8RC8Iiu+TcB2mNaoJsUBvCvb
VFb3ek5ac+eypOeUhmj+Le+NsPlwy/rkJlfHLmtZQlU5woX4PM8Dyz8R3fVHlvixVosmcptn5V3p
nE4rnskIEJiYgyyDqI54rm6ZJ5oGZuxTRsVu1f6E1EttudRCNXo2lbENRds37JwpDUKng4VT9e9d
G8Vz6mTlR5QZTOaCaH744llxHz9CbUX4bp0ckJcUT+U2UmdQ2sbnYolE3a1Waj4rhK265DPusdu2
b821YMCbCTNxeTZeh6WyxY2Bcm+TFLcZXhO2JTqLN30ZNmiHAgJjpNYM1yqci7i6ZipR7wfVL4Ij
rFFoPE0A9IQn1r7erThzV2SbDEmO0Qi3ObXddS9RiOGFRNtc3kU6vpaG10YIRhSJi+cO7e1ayznt
UjD2Q7TLJeWPIkVsYbLdL84ufghb2f0J/3vV/sJaw03TWHe75MB92RBdO3QSX7G6HaxAlIvxecaR
tuqhN7Yz7kMi+yRhmPNBxsSvm1lkxkM/aqyodXaQBmjhkg0uP2Dy0al+pc/AKaYvhv0BEqAxWnVT
SJ9JWdlZ7+q+r7mF1jtwddo7J347M0VDiz6GQgc1Yt1wKVO2xlssL0XFQ1sV25ATowhMd9sNchet
eT8Sg+ZtJ7gvuBYyGrTm/7JyJVoFnlYaGuqYmhxDQ9NipSj0SCpwfQ3OkD06ATHGMYITaWmiKokM
FBzt/eOPpbL6Zpsh1fzrsYFYPlJh4zUGr+p+O3eoxT1A9mYMvVTb4hZhqb4w8IpPZeCd8Jp0pkuT
AE4IWhymVaIb6q2FD1JXftVIYKNDsqKBCW4qYWj8wwvhO9Vs4ZylSdaS9txqDrU7tLr1LgfLQMVu
B9OTrSUYRGoP+HfrM5ugab66K8cfd3jP2FvSr6rUmtd8QdzrKMwtuhykXksjKS0IBDefGnpdPmY1
lF8j2cRRV5MdrLkpqQimFbacCQsa0FI6eN7/uPMvzT7b45i6oUaxV3Djwmiy46S2hGzo8BLxPxmM
VmQZq2zeWDWj+3PjWB1y4xOF+M8UBMeWp6E3m7c0J7OG0lFjmesIfJr8gG62pT0ROkyLp/E7iIaG
dFcUZxu1/lSRXbYcsy1ixWgj0byvszdoMtOX/uYjS4vRcbym3MiBgRBcYldxsZJ+3PAxjqnmQhVV
7fQLfZ2n0r15roLs0fI8NAteaOG2kpUetKKqtXv+hZeFQidPVR0cMJ/s6wPET9LVUn2FcWEFu2R0
NHrjXYFy0YZtrxdfgRE24V18kl5oxfVWWnQLZ/0IS7oc5SnJHKfRc99VzpSxlqFniunW/3HbUsWl
DuNPqfa/JX3w2XQQw3V7P5qOpprlZp4fqKVP3E60zigAZswhEkD6T+JKHBNQQA0m6YeiotzOi37a
HFdOXs2EuLGDQBAmJ/Af6coo4GudyznNtDe6d0wAKzuMMtzlnY/vpDlWu1ITdKJ06Ks0mhUtFlsp
ap8vYdVqX0qzQg4GH4OppMIh1H2Hv17gXRE+whUaTl98cdk3fOxASUQu3OexbN+PLpwJNp/CzkrF
A1l7cfEDQbBwR+osZfMi4vKg4SZZ/eAdyMIqtGCT3jicsyonDysZmAFl31LdVnOGq2t5R5nZ3QD8
GtQdaPd4dH/W2k0EpvE5JzOql3n6HL10+RwliPGY7IlfnRVRMAvJ4VV1AXEvqZTGgCMABhTyAoQl
DYaorlbVXb5JmRAWDtAWIkihRhNeiViRmSSinXltfq6Ee3/zV2iWLavJPmod57460DqX0i4G/OyA
P5BLgCHmAtmgnRVY7y7iW9WxkRXgUtKE7b2gQFWgb3/ZJ3HH2YHFiVpp6PkXVPjgWlslOGMR8f1s
LnZdyN5b+zym30WmsSpQpZfMIm1S5G2wvQcM/g3Xaake7b/FQ3MhZRspo3odUr0E6pgdL6p/97Q4
Ns60ERDubvnBgHWcmsCQy6PTW1Jookhc2rxw01Ho4tMvn+IYTUq5+Nr5kD7fAkWcymo07623N49M
/NqVveLocVyKHDNFH2xKQksXFUrMQk68sdj9uK8cT/p0hAuRT1+nsIipCVdYEaQISE7VsXfCxRlA
FOghPZmFRfAucQjepKFqJONOzVLqFw/x27PXR1MTmKlMeW+2TLzyXzONlGUTVzDmVVi71sLvtLSH
OuBHX2ho3ApdsrXSQua3AToO98YP1nWcKseEW1A5nMYif0CqFdYkTOKKDdRywKkpoH/PMTgz+k69
5TI49Pwh+VvC++p2N9iG2sf/CN/LpYjNkirm0i5pcQAcsQaWajNSb0mgAD2WXFJF9ovRL56QEaEM
rNJW7bqXhe7Oaviik6PMP9CRGiwBiAPZFXAU1xjRQaFZHczgDohSAhTjl5PUeIa5hxmCxU/yM+Z2
+xLb957Dcc989H4KAud4MOo94X7fuOiLRccxElwhOZmyivPNHtnBIzknSNkTSg1WPhpvmnFVQgOv
vFXyL47vjUD1nF6z8WuU5euD7ksQPTiCQ1BZuD9h2l3llfyjvmrwnFoqM8Nd1hzh748dzWaXZ7a9
zzy6gh7Acz3RhlKVhvUq7JUrg9bAAuYZe24KIoaxc+YimiaVjmVVYIu3N5ZxTCG4ozzyq4j580Y2
diVtVWLB6h7vupZCsRodMdP/FZDK2vgnfZSFKFvq5OwirjZ93FZRYWH3fF538Gm0/J3fOcdGLQ5V
ZkrWMcLdzT6B/AJkMJWXgKXCA2Vo6IU5PG0G5NJ97tn3t59sjvS1HkR8g927LREfwHRZum99tfvb
i4TOtEUiy2dUqrtRIAI7nEzF38ZtM8sgtvSgu0LicWtg0kwdRNY5CXUU0On8sNj+AkZXLiMmwL7T
ecYduKkAWTTI3ENI+ofBDknRsK1sf6/vR0wHppAOKe/u1y4aT/I2F9W3IWHwjzX4uL51adBpneAv
6iKU7aeCVZkw7df1B+9v/+AjWMA5JT7yNb1jQNaM3lfYDHFIv+VHc2HZLcVv/UYWfi+9MVSZ78xJ
Edkvxxy8ewTBg9v/VN+5IAZ9vFL1x11qj/YvnHpgJi7h8ksDDRl3QZI5fYKzBx8G/sYcicW/dUAv
8aWFtNa/SoR3F9XzZ0btl8oU/OmrKISHIU+lx2aQqXXl1mEij7vvFwYBoIrbhj1EJ/g5RNoXMDtY
d/WXseVY5T4aWANUR9FQ93AZ2ULW9NKW2b7nxK1PPqT/0E4XNkvLglFIhJt+WyZ3KOL+kdg3mLVk
OfRVuDCBczdZa21sbIGH5KdavxaP3R3X6Nlw0x/1qVwjOZ9BvCAsJtzBUI2YwON42PeiO7rAMhUr
hK6FNLgjQYd57DD0grjzdPwYlpqmbqaXR0n8/m3It5lfR63KeG7SWTCgcf95tkaD3cIfRhlBoOq3
5EdzBP763O0G+uer1UmlpBKKtSzju7s84zO1YTSIuNPWfcDtEuywcT4zzLaB1aJ1OfWgt0BQICHq
Cv6fdqv8F9AbdPQ+tfbDQNKDbSJUFm5WxHezFDcOSsRdJ6DFhCJPVAPrCBlcLvV2i9AD/YLps595
5OSAFUiJNAphU8PapbY2x8p/97ZCrwD+acA0nmp6spqFpF3WS7Cjm8LnvOelw2n7FFIZ/bP+/9eb
hqFloKhE3u0VV7uYq3c/491w6D/jshHEBNH6qsYdqaML++S4igb+TlJi/VrtV3an87HGnERXKiXN
oeYEEZ40Mc+6El/NeWbwoHHh9BJNM5rnmcn4BYiEba13mP3KRp3H+Sbqk8kIZb4PauTn8FCbscn6
MMDP2LpYJ0l7rvcy4PGFd87IpRCGwAuYNp1BrGS7DAG8O5Uvsk3/+8uNzUQNfYHBBAZqxtmMOSwZ
+NxJQFRu/Lky5fvJPsku+egLdotTXEei+f6hcb4EufrDz2BeMw0iLZmxrmfIV4f5roIUyK69jn+/
oeFTOecjWkeVaX7YSc8+rFC2Ap3Y5cBOuFG6Q1N82nJeZz26o0DqT+FHQ7MZcrC0vN7xXjlHXCO9
3SeGRFOVQ8uaOAz7RJBPCzvykrF0LAigKrT6tNjH2XBhaN2Ju2zZO0oyhP1H8mIgtg/mutTGJL/E
3tMS47++Rv4tUcF99t3G6xnJl1fJEmvzztTO5KTBunuoYQGUkZvHFQyVwYQIHpVgSR8OWeBUHiPw
9r01j4HMAORSiky1NLcjiR37ks7pdPf+fh7iQeZ7ef1bCRgvwqWU3fMKmTgtzewO7uN3H4VSOKXm
zo3R26ozlf1qMx3FNit/Ft42VVISBJLXkqXQTLWEV8r09rGo53mW/N4kEPaZHIfsrr/mpkrX9gyk
bYKQq6y1NeScX9mQay3Zdd6x6RSRoOQyZ4FZvDJiHEy5OMcbGqwrw9OUlAG8JQYmH9YylNtS7M+T
xO+r/6eLT5333jMuEz69i/94lJRk/2bV2gmahTuPeoLuV2sA5uKnEwMQpTd1Y2wAm8Q2zx6hnQZ7
yNpsvVpzzPTT9VKN1WVUXgtHw71Ztm2aaBCR29sxtlZ544cnmiyri5kw9HOp53Oxt8pv3XikkvKJ
SoIwM829F+53F9LVXVNcNBSf2Degj3LoA9xmO8he1bNB3g00joDfYKgZCAsA+HGSckPzjzVSw4Cv
yhVhNDYZ35xyDoGSLtM1EiozRWi673u8VfTqcogCWbMbYSZ8S0GFx5jNOA5FGYDN8qxfk5goN4RA
AFGuYSO4VV46S9OBiHa+deus9wff+X4r0flrQ4fVks81MzzTUbZLjRyB/cr0t7eBszj1xQ4BVzQV
se6YQEkqlF+JAJt+lClhnt/ulb3cYV0KomAJcig5c4N5jIPs4vIfzNk0Os9vx3U7CBg+guT7YRki
kvbpn2IBvm8RQC6VL4YX3kyUifiqRRYlbD0yqzwNTF70iAoGfyNo9bzazItkGP2o+xJK84MB7pJR
/542KX1WWhg8WDSrtNCMhCqpAGMHY34kyI3979JsmfTK5oUDIuAcA/vLLhOEVa7QI6AMD57b+mUf
vjGiZHU/c4vMW44SafZqDdEhTtimWQ1bINHQN2a1uvL7UEXw5rkf8+YJQJDIbr3AqU9bYV63iC81
Thm4Y1KxUrgJ3M1dNYbrazWF6d2QQE7bOOfk/NPMb5vErbm/DvBdlg07bZR5gVbM+J3vSH1OPyGi
a1aOFXrbsx7LbbrdNCyS9GwstwZFDi5qM0cnAAiFOppoHZFADEE8dkIbTh82jW8PC+N8SFmuK9mR
4mxpJxagePc2eX/gi3HjAmUJsEpbLLkW/+V5+FIsKM1HYRWct+sxr7COm9wm7wSAviGcbdDNdyRr
tcWeO0OvJYXwzJKkUqsQgut1yNO/+L1WcAFNraZIFj10+txj7NOJxDtCiJEQZaMxFY37DrCK0iWS
6Z8fvOp7Y7suNRQMQT4Oxfc3P046e7BfTXXbhSctaxbba4ZKv49wF3Isr0SBmIq3ZHdCzL3oN+gb
Ip4IT0V9LvOFFP0oNqRBx6ccxuQEVyWfIO0mpT8Q/8IMHeZ41Cd11lxNtN/WKipcOHFDoUU2RDYd
sOFZ44/WhtEqWhv/RNB+93Ip0Ikr9DUjBvYE6b8JDRgORJV4lAI//pdpmjl1oYEm8eaFvtKT5Ftl
II38aArKrW+u+gj3QmPDUqc3K3fRcGQ4cUszZfDth5uCl7aipgNJWhtKti3yJKzoeD6vvBKCO+ba
L3Pte0CmUz6xm0GG2iHKsNb6ZSk2cfgAPSUfhu8Jm27/jP+FhQvZYSq4fwgb4fQkddtpKtBhcikZ
nTAZXa2ysYR44yX2J5udeafSF+ppefckkkBj6OyFkzKEzhfksxrEC0ZLSMGTl48G+xo/uuon09t+
hfh1WhBuGfSR+PRDgdDtpObwzJURnsqBIfDWL3CUitrdCJ8Mfz3vs+aHJ4WxdNgCm2qNCGkOGFZ2
iEA75bUte6TAhBsvlpLQ5V5mxaglr970yu3VT6sZCjto1hdpdL99j0FCTOPbju4QDCdGXzExr/YY
iiM+KiGJGbKi2WnF4v6yRC/P1Ov6mnKW2+nYE4HnuX94Qb1XiJX0zsIETeeYsWead0O0r4u5lIGH
fTc+MU8Ad2xi7BxoBEdCJtlpkSUiFopruOxbSROhphh1oGPhzh/KCNO5o4tGJkew7XgT6TLl07O5
p9XL7Ma8vYXB8FJaE9jbt3i7GYgIBH0NL8h3chZj8DQvZ9LTS+Y3YoPpLqThoCt1aE30AHlY445I
BE8+QVVyohFdVaIefvDd7O59O3KXN0eo8CY2NUh1+jl/Y/FeUb5RC7WNdGH74KzkXflGTZmNoiFT
JRee7FWg49CnFYBQypcDNODm8OaCFougHMmyBkdKRRu1MmzpYQX3NR9CwVHKcb0/SsV7SDeAHLZE
lkCo+Nrc+jad2va+gSRWcQDwAOHXHvoc3tYL9tNmjcPszt7fYA201cVj2kKdANWpu70/jdXssAIY
T5xr7QktMd+hVIwkwjhA+d/+C0eKXACTnA71F9StRK+muM47T+9fUuccYuc80KWckgnlEa1GFOSN
o9STh9+pVjYG69RUkArkyOHMH8KntBndhVnNgtXTCGrQZ6Jxj9QlgghNPjP+FITKNfAAItLF3xPN
Vxj/CKxVKaAWYFZ4HTnsJBP2gFx6m4fvKtnyCqVFSiktiBzerPkEwQmOe9rT0Kodeajv9j3J1Z4f
R8K0un3sGS6T8jTpLOXqIKGgqkqkg9PmznHR4tMBY0xlRuoIrZC2YLlC6eT4dRjMhm3A+LE4ZYdI
2fbJQBZhLln40Tvd3t1nxrYT6edzL4QHYaZsVFF+YFgX2BAflRcL7FWF8wyhg02r8yKNbEjBdxdF
dqSCKWUZDSycuWDGjv+lRynRJHCWfzGgSO+Q6Oz0Z8jGKjxisELATapIFJHwGVrwd927b3rKyMqa
PCUtTIogJH8WsX0eWeJFf9euizv/VfzqnAdTjRV9Hueko3swcyodxhKMHlTYrRXZo4ANrVbkY+2k
3vTtkMa/GYH3H555SvI7U6HcuNhW7qAX33zj6iLu9ISheyLiHUVACA1zYr+34xpwHxcjTCnljyST
565B1sXsOSt6m1AIF6s3+06BfnI/ooE8H3BDWba1LWjsKmbS+6rh82mYCRTHqTt1fyqAHLprEwQt
CDwjCb6leyTqL3zl6qjWk/qrM54QsISf4+PJXslfAB15bnpPHX0iDSqriMfL03CRnfK3HX69Am5V
3OHQzAWFjqIMvnsl2P5DnYYGA3s13jS3ug3jOVxM5dMa92BcK99h3O+4OyaDGAG8/rdUK+5HhP0X
T5V+ecRNGGynAOmo9skKBIovyFFd/4Hq0Q8Ml3Y6OxqByaPiBfACOHFYvDBV2+dJkXcTebu7RAyV
x1I5jzWqN3IjLEqFHETJCEZcJKEoVPW4iFVilVCLO9WNB7Q6gGLZW9S73HfyOYlxGzT0BTxtKdeV
Ho5po4Akf9pRA3511jbVq81kbq+R0n8fQXJR7iIU5EhP9oFmTreTg6+ujBUWr9lMB8LJcrLWDCJC
0P18STC0uXU0O15VAR2mtKBBuGlTyoN20YARyQ4VTHxGr68YA1PYOGVfYQ76BsnZ8VyoM1kuWv+x
gJ2XjPS6yXYXKkDqS1YqEUj4JhbfDanvGrpiIXyDO6LYoisgeJ2IzeoInMXj0ur2CeHvH3vINWs9
16iLi2lpOpBQyNUXoPv6KkiJNpx5+d+Res/u9XSIYBCdGep2fgEgIchKZ2DLuGgFo5LuKeDXfxmi
nTTBcP5ZybSscbnrKkPG62l6T7H2AOsiWHVog4Ut72MRfxBX83Ei6KElgjzImBUjHIi/UrFjdaM3
5JPcynIe7PjRfmjPlKe98EVjB53d0p6qXlXGk2p6fUMsY9jmgnUhycugf5BojJhnIzERcbSEmCMH
11a5GI6RuYGehP8IgYUoX1MgK2jfos8TDX6Gy02LIVB9XxNcNKJt8SiDPdTmeRIX9Izqb59r4yT/
SHLO8uPpQFwJ3YCg1zjre0yiQ/OVFSHUs2zKs608FmL3NuhO0J0/XiI9UqmVqg+AnHGJ5uGQB5M8
7mOGvGUl/ZKx6Nu1J1lAvmwRRtHsIMoR8D1j/VIR40lOMseT3ZEH2qeNAA8QV275mquyvW4faulB
Muencs/3gtzG1/zZU0ImmFvJnnYLq5YfWMhHCv90WKyYaX9d1hqOEDCUbG9LbhQGVTK+QwfiVP4v
57wppOWqd1phjU/FuOrBdVAC/tgVkr5Us8ivEYNXnFlJUMlBkkkEhsg7XWTfZ0nDB5RA5ysbJ5kW
dRy2FNZ3aBPvguxcKGFs+sVH22S9xTAWlDFDSEH2be3zWzhuvgGszQ1leLnrWcWnK6P8tvBiMWKp
tclsrrASILSqVvFGOuGAP+lVB67wILF7S/g8wzKymbs49KxVAm1+0CecjQ+PfdM1zspu0f3aKf7X
/WGOFlzFogb8yOhn/hibwpuGkuBAHC29Hv9RUTYDH9b/IUwxliJptq9JtSRun8NVf4wSSS5ysymI
QD2sg8SFPw2A/WVPTbtbBuo7eRbmMEHHfj52RvlRbTUExNePXm1NK0CRk4492j0jODBtfW54OVQr
cuS/Lh9lDRvMCq19goXXk/8Bfmr383SmKhkw8A88XoAsvU3eRaucT5OCmsgmLyf3hTTJr9QLvkEf
yhY/cvUQvaRJFPLMdBnsCAldGpwCgpqB05WUILoGvgtojZoSBSsAjyCag4JElq0vuaOmY2iLXhzu
wEfgF3XcqKYTsVtB+G4aDmGD+xbOoA+/KGlYW2/CmImT4q2v49Z6Zzh5YHaFIPdtfxw03N4hYsbp
woPaJXaa83zVMp/VUICwSrm5CrF6oVon0aoXYipVudqJnk0Z/QPfgXgXGnSTEg/zHdBJbgdBIlL6
PmTMXcf0HZQhbc1QfFNGRldE6tliSePi4ZNT+1gOV3Gm6p94im0SzYaipuecJh9PUytU2JHY1+1H
BXXrE+3skWl7sABQPrVL6T/oCXspj9/iBzw4zeapoekITc9C0Npj/+HGDWnxHzK0ldyaMSjGb4y0
3+EVuDFCwpDAtZ4PgGBzmWyti842cnCgxpqn7nr+A77qcNArinX5zW1dPpdl1VMjGsxGV13oh3N3
mbX02KCwu3PNCxF9EVzArI1Ihz11mrSmdvyYPaDb6p92zksrL/NmcxHEP+en+Wml/YQKNRhELZ4v
ejT701lh9+g2NQ3iT7EmPY9gv6mqEx5Cyr33rTVGXt72vgLjhep7tvVLT36Jq4B8WxpZC2fBuie+
f/GZ1jmAOlAnQjpvpLfUwdmcBhoAgbmfTB9X5Nj+Z0poBZrMZNXKfq/cYAaM3A1xu+fYd4+N8jHW
5gLXp19HDPDr2xZwrE5GAJKCg2oBIiT6PZbWzR7LrSuAk2B49Hf4i/4CD33IaSURVM7IhGghnVIv
2yAKsV7limsxK0q3YQ3Mqb4KgnFFko3kp+Ght6oDQ2wTw1fKlBNVPNqkIqGlgIoqmCpTv/nNyt+A
q9oeLq6SeqeN8in7/ky1sUGzjCWAIf/9zeixT04NE4CCNenz1Iw2hFIdnXRHghjIs/3MZxbxh87+
tPL0d57U6OFFFmHB9AbRlze7/yg2s9WyS46ULFzoNo9Ac/er0K/CdesVXLEXUUxZQDz+/MeEvICE
FW5eD57qJ7lPkBf06fbdTfHbiF5upWOvwqFPHdHgbExAUuZ1NnKu5NsOjdF0HLUFYXnl8hLLL6Yp
aiAnFmvHNyRIew/BBu9ZVm5HRUTGnz9gY+Lc6evR/wqg4hZsRvGzwSGX2pHXBWi/QPno0ioj5MJL
y/wyUl3bqQQayzvFhzEzvPyjCL9hZ4dweC+7qX31qHNegX5q5q1olA/KZKyHqE5f4RXOlq/HOCWr
v5LHNjLMShqSH1LMiyZXVPN/+pmAkHXatUhEgarwizbA/xnV8p6QLFRUN98uwMC8bDf+vetIaNZA
PrwajtgAvOLo+EkrxqklUxSSQDOp2mLaumiymvc0yCW3s1PTtFQM7DZe59915/bp/9mrKd07HXNM
PqT8xsCH4IM35IdTTJMARb5o4S2Q++t1QRCG3yj9yAbQTVvxsEn1ZBRG779L5XK2BrVaeRe/yPGt
jJ50cdChVXzgkSn1AI/EpyNbFS3xKZkk2YSz5GbhgBAhnz6CtcTvHod1hSxFPl6EAlSwSnEY/jhT
ZuIjrcwiEaEnZxoT1LFym3lQyrtEEAuYEnM1VxDEcYDyPe1OZSylT6RlS7kYvvpVj6gLZw+g3YIE
oSgJnj6Yb9HINAI2tRbUw8w62mFoYjHrG9M0HGynspl5WKL6n1UcRF8O9dSI1Q69zsOjzOr6Vcsl
LRFcT2/qH52gB8OlARDHgD4KAaovqacMyO/8gBTzubS+l/dZdwlgZedn+fL835+/say8pKTutUZC
9QedpK8uK+7HBSJxr/KK+16u9Wpc3OYZAnGq2C9kjqc8J9ZFuPHU/eoeuUwkyKW93NnuNKXds2+r
gNCgKjAqF5FNUFJWz+TrDvnA6rCPV4ndvqao+omRdjIAGSBQ0oUIwnjPYjvCjJ1zz1zvjFdcuIcS
KQAs6mAW78nKJJ+Ll5VLn5TyZNVqHdqmnt5WNjSbcYj9Rnqk1Le1r/tx87/tsXh6fU2fzHVh4ENV
pdwhXZN5xJ3SSuG1QaFddhqdLhT4lX/lJT/V3K4w3bCXFnO8jeuFregeGq0pzEphy2e6Od8C8wIw
u04ieOSF4tZtFxmFQzQyjdDvua8LII5fEAW71uohBjDRB/tXUV1zgQU4acin5PRRcFNtImnhGDQK
tPMjHE3yXTf8rGPaU/atiIVeQ7G5AF8WDypoqug4xKy27HNt2R3X7DzivG1aq0CQqjLbTmDRD9Hl
0QAWgHv+nyspyWTt/+bhuMONB9vWpXCK2s/2fvabhrGoMpFxj6A7TKBdJhimhwPqW+71bpKoIMzn
5zL4W+f9sdSWAiyIJi7dL8xZ94EA2pTFS9LtjaT3Uz30ze8Angt8ayeO7kyd6vECo/GacEfVk7MM
MbXki42JfCQLoA0OescBufgeSFcebS94f+O5yqogUDGU1etaOMkGWmcOWAwuRVQ/a5OIIBD+eLWE
7x/T9mSGNlmxXfF211bA9/8aVQrqCN/JUHAa0MiXlXjo/kflVwOZltE/fpkZodeXijpYvJ1RK93R
vNlJS23OEfYbogMq9lD02+7OCDePrIJmg5yq43KSAtxP+5YtasKS5P5TPamqLQHNrwN3q5hWRTGy
NlbuKik2r1t4DjYQsZysu5oGoDyAxlUvmWnBmYJwyXv47a3IAGRWL5WA9+shCQIDUTuLkQLS+bHq
ZsdsRPMwIf6H8voubZagO9OhIK8xES4Z4G4NdL591eyFK/Ti+/lflfMQ04gTXxOZ25mZ945qIlVc
3ad0sUmHp8wkuBlb+NiErAb56vaO2HXfRo8q9o5ucegJ0KqLaCxFa5UnzierhGAAgxpd3d+LHiVM
nDEH5ipmzB9RTYKUhdQ34qtZmAU9aiYAeV1uSysx4TlEHIahmkF/U9+jnyS3AkSAn5pHFgQaQf7Z
ethgIDitB16GEeO6T5g/je4Gp4d3TfRFEOvJs5BRhW0vnf9Ys6hUcFbdTBiR/puuNmN1nSKA/vf3
ao0gDnX/pCAYMUXAKVAYFAdHFNSF5JFMDy/N5Jt3fzQbE+R1iOIeky5CeSPMZhN+B1AJSGdrTnQD
f7Jr8xhqIYVmP8FArAjSgMzfamemY2fCqZbF90pyGBYvlp1iWH3nfo32ZN4kv7vHooY4BQELvM0J
cxpnWps2Meo7AkXE+SEDwSDv0atLWLo2+GTomsLZzmyvP020Tue21w3a9vhOuAIEqKHl/4juF3OO
1ndD+VzOobvMC8PY0q9e6ZJlcjYsrPAaMxMN2W2S3rHEYfieNaYWhcB1vOrEMyixgqKxBLW2MYwF
jaWVVN239AIgEIoRgo6KFaW+Q5C6NWdpxto/Nt4ZSBX7YEHWOmj9cBVxSyHAtoZrwVADXSEr/c+W
cGYlmkiCF+bYVWogWTwSOgh65tx9WSNWk6n0KtBgMv+OhNsE2f7UAZbl9JIIgPBqv8+k3qczO7Od
yiXOEwBGtv9v9GToSGvVd/ildOon1w1dqx+UrDGcNGUx8RXY2nWERn8FUQjywc/9ARFnWTwkh2VM
GPhdW17cmev33+ERt7CUekkO0lwVnf2vMfJlK1aIUXqgNBZrXYgHdB/pyhoKJVqo/9391bkb1rKR
M98U51TEi6NJGCTZe2b3VCPPtK3Pw5Z/E6Lhk+aegcoUtDMkLE1ATlIUsGrDVyh63fJXoCoo0bOH
cxbJhhD/+/bnPOWMNMsCFeHnBQnbyK2ueOy+SrL6Ob5kPouvJ1zcFitaz/OuCGcIbvNOkeIPpiy6
1RuZ8WelccVGT5DAKtpgWM+pL9bzq1wgS3L+0vGs2mEVh4EB68SY7R7948sQo5vl7Qno3sfzJuVI
iAVEoxLfEldxsdICdLwkni37QyaQ8JS/ZpUdYHuh1Cd80sAlykk7wEphKAzUWY8f5YtFaZRGI1jK
xqFFV22HHLqsALzvdx3j0vVqY1DVxP37QflAnoOo7sjku298m9XtsXSrx0+eP0qXXvYtIt2t4XIy
0wChP+Ui7qi+a9M3Ywmu1b1Pk5uQap6Ocs37XGelOeY3r6/D9ytrGt2YBL/OKaedeiPQTQ40phL3
MjpXLD1VhzlxK6xaUzWxl0NHpj6q95k3FKdmUaaURmzF6vlWlu55m8ELe9+9jnyKLF71FigXJnzT
sHv8932oYVG1hfs/D3huwQ/bwrD7XwPh6x/kO0apg7Tn2ZI6CmkrGri9sf5iBK1HDDAaR7Z48pyk
2JvRMMcBWXzsdw/+reKK86YlzwsKAzokeY1PUBKfrss3QuByx2oJqn+FhqPO83Q7XBkH6dyRUbKV
SL3zFR7Dkl+PsmUEWB4MOzgzh+uoCDsuP0VZBy+7Yzz45kZ+MnUCgdxysuW0wbPofCqgXw21p4+C
6tdk6Ev1feOMrG6R5MWIgDxrXScH+5xOImMCcP3M6qgspAiyiupwwiRKJu/yJysu+nLyAV5bje91
fhUCjVQCPBCBEq0N5Uq3k0jQgCpAKvRGttZ9ASkT902oOQetjRosQ1Xh8J5Et/v8gFTJa3UJHz7V
ovS+JTbtzlgh3JxZCl87PKOn+JrqyNsYlNdHQDMWbky/9+gUR3ARYsdkOIvi/KICeHG/zOSXj+Rf
l2X912o6Fzs+t0j3a2l+CU6XIfxXe632Qtn5Fm0n4F6N7UxcatVM9K8Q7/XxoNcA+bcPV607JOoW
A86RtmfdWyaURA+iHwZ0TjKyXeZBclsGqoDgwaBQ0242z9TXe6+fpiC8TSkv17SnYAzQZ5mHcBEh
lVDXSr1QqRYSIv9NVe/WHPZlmd6C+bRjZbI8g+/w2triLJV8zHC2HfSwyjrNc1ShlJtXPXK08rmq
bSd151bgdtR1qG07UBhNPBDa8opliRPp7l1YXXJBx80NodUdiUF7LxjrMr2zYibyaOrY4+9myJSY
OsWTFHguMxMmS1CK3/rqWVG1d4M5qgBlt5swgNI+3yTSok/LqIVp2QEryjo4W9FZtLljD5SzIy0F
Y7kO8yxeHy/QfRF1rYC/WqVjrfacDpPZZ7NGnv+MerIplQv5sIh56aZOlsCNWuovuzj2U00XIgeN
Yf9Q+Q6xaGsFXysJenZCHafPF8grEZ0oA0dS2PpXav6uHuRs80FXhvNWnyOj4IO4yd2Z2tFKK6CA
EyinEd/G+fuWZUQAb6EHS16e9UD7bID9PRsGzWW5jz4kXvCLi6eYk94K8RVbYf9Zpnvwc86RivtR
zE4FkarFbgtJYtgKmJi38ISl3FDnkHafmot/bV9cScfbHFkeXO4WyF9wo0o0IGufGQwh6fSujRpU
UH2VlhRsWkoAD/YSO17oQX+SN+QX6ld+vxjLg03vmsS/imhvfwtn1CKaxyz3LAxZ8/BR8PIMd8wQ
OGx8uuxQ/GqOdYUEmgioqKlmTTLCStfcEJvZuALiiAgn3CcSjQKZzx3sy2rgk3fLgoOa3ZyomtZo
3/AvLNbaFOM3rPGIFu/RruuU2XlOQRHJ/Hm7dn77XExGz8BN1gvq68fb+Rx2yUoG4ZPYXe9TFMD9
BdpVcpKCJ0cuQGUMUA438YvzLIyed2z+9sxOXGo12IiAx6N+QrJV/eyYlWZXvCkCSL/CCdrUqt6x
AJy1QpUmYx6ploMHFSQWKbJvW91441CGl1Dv6726QxMBJTOW4rNKUbJ+ytre8recJssQz8F3t481
v6hQ0vVIpASzzdyZeZ51pp666imzSbxGl7a+gTNxKjkxCX0VnvTCRpsyI4J0qNsRtGR8wE7KccxE
z508HfvSrgGf8nKRP0L6CfcyIsYCEAsKi2L7ARYh+Ocg1BgI/WKY5QYQbpLo5PXw/u++JbYtWBV/
ts4i+5U+BdQaj1mttl2kJPruqvH6D8rUG+LYtls5P2iAJxdJaxBnCBuggt/p2UJGPnX1urPx/qjj
7MuB2ltpZly0oq4MEIENxk1Wfa8DhxmFMAv+jDPpT1ZYmDulGmQl2Kq/pIdUxsUrUVMrdxDqhzUn
Bkj8bvoe236siqzFK+b5KasUq2ViE7c5IshiiR4bMIFZBaK9pRyNw9cNv7MDa1A21+V101hVIVtn
6BUandVk/2Qnua33T5VVnKF5QvelDwkadoLceWxiOCWjZqIO/DBI66gLgE3YVlxuEn6hvw808jIe
R+8glileXj7JHd0/jy0x6pSju592OTH8YkzLyMOzkvVEkng2qZO2e5eKrYf1OaYUnqZet1Nb1Jwh
tAevY4ql/IsFW19dhuZ62Mpdx7bNRrB3LmmU0pC+itYiLdnO+MTKjY8/NYQ+ens5f0iGNC7nW0oL
PoZy/yMuOzTGlrkDekuY5LyhrIgXaRsuhHas4cVkEKTV6UaCazqAZaeFv3rv66q9/5Pjf//arU1h
6jKsEvRNaQM00mpdXUqyE4hTFEkjTrUBGmdewRz1fFVDIuxxPz7QS8PkdYQ68LIXQLtkilcJH4sI
dknmxmvPsOyFBBhsKDkIfyhrso4ZegVzMkDpTI6QfNELjiiKJ/2ArwFMd4/DLYBpuc4zPtkmT06V
PZi2WlHV+Py99YoynQkZ6j0W7mW/STVVzWIcx3sJNQQVftX+8t+9Wrz5TTWrQlfanv1kT3k/1Tom
FwI9oPSYitCs0jbzzX7oizifkmt2f2CUvyXVPxG2D/NzRiiQOorBoBTL06lKVszzkhPn3QwxCRtn
jk6flioSw4dwhwTBV94yreWUVcAiXraeU/DCQ934z0MD+XEmcFHP70uUV5qg2s4gLLe78MO3fV0O
SZeMKoq20DmwCtVMMQsIgmqMbxEWS3nCFSX0ge4T1TQqKm8fpS7yjbGj92h+gbL0d0oaheSlM74Y
QlwpbimdLvCJem4xoL1uU5A8hiCBSAuIchy/4Zu3/GILR0skdatNQi6nMQUQQ1klg5LgVckGrLx4
3NKxxWlovoCB595vU0ZRAfQaT0n+CyFOUjX0WAtpkurWBp12j4rIKofr2ZyAlYYqRhB/IjjbD2US
iE+14X2jhuPYgpu++hrAEviGUNmmnxaTo1a4pNj7pG/xxSnElHZMo47HYSbB+L7tfZeZxD3DP5up
Ao16+8LpfZqbi1mxj9ZBvEtf2mzxMsIqPLyX47vYFJK9mazrVBS41v+2yRza5AGpjaeobif6yRSg
4KE8C0ZlTVwIDNNE1AcApNg/uEefTeBx4Tgcl9K+nO+7+lza/v/j1pAaBxE0eiJlH/GLHmP0C3Ew
Swb7Y1skq76Czwiy5uJmmm2Pgg7LW+HzUAWgwQWa+t56eHVveudX8T5dvZCyPTO0xmfRkpEJGWbR
i1z+dC+xAvkzQ8TAt4NjAmCyGHCLHSWcAAONZl34bda11n4Eikrpsa7N+vA67bfQP2eoBf5G1ZoS
aJvcF8OEfpAvb0wyQefvROiQyUYQvX5uZQoDh7PV96kb8InLIUh/pVbpzJV9gteN17g7nvTS4YSS
rbNAZEN183Cw4gES4GODGgKXo//4boGFpoFTIRuSfT2CHSSDBk9Cu87tte0QuA372BJ9e6tn+ZtX
fA6PzXAh8PKnsUhYcdnmB/dda5Xc91B1Z4YrFc1QSOLGhfGXKK/DbOCtFVtYb+m9AbqCtHnpZGeO
EKe1VMFzJfMI2ePXpmiPrA1/JW9RZ/Furq4pOnCnQ3hLriK9LrN6Ah9XTHjOJpwH9YpFTfk+dsnt
Uw7bmRvTZatretG9YqyUXhj/bufdIYxOHeJ/HDNR1ldQaSK/jmJaXIOOIlcp9oPXd3JyrVbIy0W3
pfPyqPuNxnvUvcvQdp+DGCrZD7vdgSqx2zTJdV07CLk6vRd67vEa0TrwEePS7zW2ZxnanoZtaFSQ
Z+33Pue6GzSXqx/ZxUczHyzcf5sEyszu/fbfCeIKsY6RcpBpq2WIClyzOec/Dz3voa54PXPs6xwg
Duzg90r2VgESh7/vx4vrIwe3up2Sa9gfHG5AhIAHp/pFVc0k5VOkIJyyoyrEq97Ls7c4A2FP2+IN
r+ll0KoGK6qwdbfrbJbIg74NvhGxMD3j2sr+Q46hha4eIwfEJxmyX7LHFNXqoWe+BjluOf1GRMiN
cWgKp8t/JJwwOkza87qJIt6kKh1r5+a7qkhUupmAdKeFh1kQboB6mfBER7C1pPYtQBeKP9+MR5sg
Pg6bLeN45VTFSFlM99mYNltZZqkZTPruWLyQB54M0yejG0nTAaKrrwYXxDky7IivW8T5QGt6KBls
IXkHYrroPV7cvCPUxZfKB/X073PcrEMhH57krqp7zZ9w1aal5yTbt1zY04hg4adzr6BNgQhIi0Ck
dAP7sqdsSh1BJppVRziL3lNcEwwoKzewtZ5JCOopKWLw+tz/hfqoeRR2b1ny439sJ4qz/imJqvvB
1mRyBbDtsiYCyP5H0o3ZUffbBUDmqy7yWCGgpfr4n/jYKUEPtrC0pT58kVoJKJuFrSKvTwm87+mB
y4xKfCXbOGNRbEtfKTicCLjiYKtEMf8cSyjimCWf4ydJxkIssol3O8KdFKW2mmaVxJnP4Y3CrKz+
jfLkYv1m2snjhY2oU5lmAl3+zg1NAdkgmXyWEQmR5nS4ku0w+yk5ipUlS7ZQFF3tKGuISkSyPm1p
TGQ8h5hyfsAvm2RdEAEku3rttC9XtItIIinHVsIK6LTIbalgzPSdIOm7hnvSItvFhaQLxEGv2HoJ
dnZClkNbXsCNZ8MJW4uj+khw+kQH4rPd2cEar+sN61OXFBXb+5c/q1Dx1HmhFcsJfKygq/SXNs0h
l/tREhS+91Im1w/PL224ITcA/wQ4j3Yc0cai8wyOQgt0CuI4x03Fylb5Hqgi3zSXj9e60Kvf67qW
rZyVATSrED6UoLTztag7OjsgUXmjYeHMXipNDm1iCbwjXFjmDlPTdssYh1tYdcJmfoZj6Cs8ocp5
U3EP8nlb0CNmX0smTqWCjaYLd3XzbAEM4oLFInDcsiLAhcH13C9ph0yfja206XUdESejqaXhf7i1
wvejBRZt3HccSEAUyfgDytPHfp45qRlt/qYIvbpi/ZWSz8VCx1Vwkp2ZuJqHb+ioX27O75AYkhdc
FutSDoZil1vCyoBjk/dMohZc6R/gg7PmbZalCcqLw/0tk7jFtfsmtw866PuVfkpwmjCXNRxpKKpo
qhWV1UEJ+TU/8QejstUMWeEkxsRpMWrJKWkxcOSAdO4h4bI/Udnwr5meNcwecinI83GzyIYDTb7r
4P5RFDwLouuNB98Te+D2j/U7upmY3ZjVI06G3M0Wnh7zMOJXmerTkBIK0Yplcwddp8vrF12RNNt7
PaXVsJ/XETL+82WNsese/YRh6xKbjADNTiHmSBdcyGE3qT3YTMBhw4kpgGjnmmw853EhIeHNdKVO
ck6NIkDU///5hONhJ6NUrLwKNQCh0qPQA6Bk/fL/qHAyFMTuptQ4sbgzlVkS45nRr3CxkJi8IwjX
d6V4ftLVCu4d9jqrFQ0f6zYbUxOed+iDQLbv9/CTojzKjQSGufRvtzF0dpCLIvsA2ZKywZBis/JU
nNk6F0mv5KVQNH2ShUm7VlYtLnwnINNQsLLroSYaNg9o50ufwhx/7yC2tem205eH9t85fW9dfHSZ
PZ10Aa5Q9vfRSdkQyH88vcN3MOB3UB1FzMJECBa2VT/O7Zll8zd2PdyKQqDvv4QGsGaZO7ZpLJfU
UsbsvkZhoezilr5aHq4WSSEQQL/8GfnpiFB5qzcgmrKcdP+jsSH+lwCyaX22wCrv2gLZfRqXlqXg
//hJV26loKKSqOkYE0ckBQzJjnrAt20g7kaGJ8hYDdzjc6avcadshh0+F0CTn7LzlWvNI3mwhiOE
dBdpGTgEVy8lo1JvCWF85A3uHqrCsbyWo6fB2yQ4WDpafmzp0/Q/Wva6cqC+F85SD3fxl/7HjoPj
hQojSEewp+vejP9+xd0sfJo8LNnO61ZGL0vweIIGog2W/MWXEUodnCsS1PlMDsCMK2FNfJeVx3QH
1l/6BWKE5AEqALk/kW8ySkwakACZg1q3KnCAbbIhXilinUjgqFNcQuijdnNPzfD73XIRPKDY3j4I
IS5HpLn3yeW0lms4negaGV7ABPGUKp/s2bnJ/nH72OZz8J82d9q2tA2X1mWmUxYLXjplSd9od5zp
xCimJjW5YQ0oPI9bCDYio5PINbBdy4tdVuqENFC3GLhLPG+MTi3S8XhTcaoqxwEWChIN99AYgz9s
+iUQJM7da0+2RtugRkRVDrYcxGqDw9oi5afTJEI77dBkzWOWUAekn6KBaCNsvmTpdQNZO4VEKnYm
UbtWTBbY8S+Jg/i5P4uVwHdXOa7CPj0aeJTdFY88osR8k5qcEcOo/UlF3CYw0nG4NL8dUXeRGgaE
5PqH3rlKuMhcNfiLUU4tiO8YvBveQ/113YBa74p2XqiR/bJnUjer/O8+2sc/tmOAtMRE0Xn0xEM7
56yPzVuHRUaSG6XZg0tLMt/+o13A67PRmnjRA11d5xl5AJcWE8Tq+0S9kaVVOpIxX42ZoqK/x5hw
iIBuFhejr9lIpD0aM+xA4bsTozuLoCzBvorK5CfDGc7xFLO/0hxJhmeV6Jj2Ld/MPyBn1e1OViQa
DkjEU2ypkWkmv26LdgnHz8bYtrFOMeDBZu17F+l4XRlojI3g5oZxvFRi1liApZJFuHNuw1FPiuRG
UBkEM5PJDpRzFAkpu5wjxmRiVXZruFt9KaxSje0unBn85opo3iXwR+8A4avomPMI5+ph57raKe4a
RHNdf72BEFP/JxEN1pHlZ+GimuXG1KWsP9d7qZLgYLH353i+rji+AJrKkkZg1oLlPHo7wLEG3XRR
5n/zBnhEpgptsQeGQ4Q3mJwtkLu+FS7/w3D8RGOc2MyD5P1kmKSBuvYRMpq7wXYXKaid8GgbumJh
yH87vdmiAF+YfyvKfH4kfUPlxN8UY7A3f9twu4UBAd6096FMc8FDxPcmQtJS88Ej0dL7fBNMhOnU
FTlJNUsBUkCqyQPrX73jjKv3KW0TPehxOU8uLxHwzGne6b0TUc70GukxxalSVcSAnt5hNTEveCxu
O1lMwjIIlo6HzeAIF49vjF0BIx2/8N5GmqO1cS8GpOci332rbVh4F1eDtgHeE3s7BD1EdNfi4tsX
muOU1drPML3gaSyHALuU5CNX7LXfFszLIuPA8hgXwbr30w/lqcBSVfXXmJe+qe0Wu+o316ihS9Ii
arxK5F+EzC3WXmbGZk98Zbe/SAkm0YRHqXZ0S5BsKWhglo7UQX5WbYp+6C8+K/uYa+0UOEZy/N2F
/oC6JjPACuAe5z8XtQhaCcNAcsj1AioxIBbVaBv5rPLy0dNiLM9vwfFRY+AdJJZfTZwvJ3lzxIvV
z3Vph8rtdH17sKQKQfVtpk1FPcCdGRxLjRGJye/Q0OjzSbIqExJWg1724jLd1YBxsFDDnHvnd42C
mZhSqMXeBfBAE/GWHRXOVZ+VDFrGLIdvv6uLjlTVbG+GvAqu5VgIn2AxPr00xwsvyWHzRyffxMbR
IzqtiDK9lxTz/7Yeb9zPHB8ti/T8F82mGXLqOfp6106NbxaJ20gX8d3y72OLXhC62aZNeaiMyY/J
sPPpjTAALFThv2+TBiNSW/RQrUSVUT7uR4QoRZu6TJce8h0q2JN1ptExa3f6WKdasn5XpdE9/6Yu
YwTtdhGtrtkkbTV8nJwaNRMJAbQpfcO1uyoXYaZUaWoSDE9yL4NRd8kzUrpNmVfdL6+HPdbCCYrY
yYIkPnufRqOo6vgHmvixGmxd/P/8P3YMs+xTzBgaxmruuPwPxAzPe18+MtOyDvtEjjSX2NwL0iEL
/BtHc4gOGT9nMudcERYhMikOSSJL8LVVQUSiYFDq70mqmx+87HxNLNMJn/SsF80/dwl1uZwzQndJ
5ywxNc/59xodZeCPYhD3plSFt/MuD6Ius0yR44E/SsuMnlvjzIJOByyUNWxYAQouVvY89DLzzWkW
rnAAuet0AVh1YSalE7FTgTSSXhqITFZigxKvK2mVgHFohCQHx0EQAnyzchhJCvwRy+9famSENNFD
1RVYG2FR6SuFlrIefu3EA8ClNZZrcf5hvPafhDxIfV/ZlEZWYyiej2dbSDJSB8jWWfhYm8pYw6e6
I0a8GrUhzWU0I8Vr2XokM/dXTFzm2D+SZMDYZ0VkbsM0JS4o7yBAu8ElZA6W5YzvV/RLQNvC6SLu
4KF2ypjl5chdXiasS7NTcRC6aNWP4cQIaz4fjg/H5eRJcMKsOnuCuky1LcSicCZSX6tRRcadmvpC
eSGlC6Jqm7fMzywC5h19WSpaQaxsWBE2xjJDgsDFoUhDQZvdlCPF2qd5rGcKXgMoILuiFef3XFKw
2WSPZhgddyLjsdu/ntAedjLJUMO7bfoOCZxsqI6owfR8f8d10MT3+jCwhdtw/3mN014hXXo0SWFm
P0TY48qgPcAGRSEmf1i3Q6UdpS1zBSJBOQd3DAk9hOzHbmRjpJLTPHScIfrbFFLNHOrwdvphckrR
M5kJ74qtU8pYFjhNXsbT35bqYaZ2K4hby1bJl56tC70uUe7lWBK8d59nLvge9JBn5bzM3414wZez
yaiKYnvcGRs+1OWV4OyKeNbi5aW7MXh5rBLbtFml/n+vhDFtsRJeMltTwxMY3jkHUg8nkkCUxVJI
r8pqaO9PM3dsVaFdR9b/aqeOMzNG30Poqkw2cnQMf7B8wnkBd19ZP/cX6GRNPScpQamGaBecmEgb
enJ/F9KM5abpHEdrkzL5eh2xPgIXTE/X37d2cfv641OsJVgmyxU1vhIHHaJtmXvz5lCM9omZz4BP
TEBRvOmgxCjunaU+Ckpjguc6CkStjkSJOUDuWRXRl+UYsaMrYpxY0Qpz6Fj+hv6EcHc6rEPrTjMc
PCRTdNh0w7TqzI8xq+fxK5x1LxwYlUSjMxqvNtUfwDaUqQGHq/f2Ei7t6SCrZZgJT5ABteHSi6Ej
fCMeH30QO9TNw4bZhpdIRCQpG8+UdGYUDmfvHiikZRQSr8xDNdFkgLCKeeRykDrNqQjQivPc/n5e
+fpbARJqeGWLxS3vapkwlYMQaTt/leMjpZEPoqRcYVhxcJvhafsjDxJ1/DkAGCC/xSwV78pNuF4u
nWptY8ZYnqBcWuTUfmEwSukRIBCbcY67csSoTBj5PkxaJ08UZ9zv116uVL44KVeHn5ac0+qvcgTq
x6Zg7nF3bTNC3vp804G4aASmPyoS3ijn32yc/wvl68s6iQwlMYGcW/JlYURduO4wc3IlDQRegTi0
jUBIk0OCIjLZZviyP5VOyulqpxQvKAutXPCRDcxl421OHOWETaC9p/ZUoyiUYZTQ+WCrORfRrnmx
2z8B07Pz/WCdwMIeITGvqVFmgbpdC03WBf/H2ZCxwBnkSvATOnU9Mbi/1/j+2zyYnhbcH1t/UmeR
wSOle2aJcuQdRtmfcXexA60hrjKhOPUoi8XPWK+AX2Lt7CFjdjn4maGz91kpPqODLTmkS6QPXNme
XOtGn90FoGMFTn0YVko2uTOUjnYiBCCY/AZkDqwOf4LvNwTVEPyiXyVK/zpnyx3uAZtauUW1v05S
8euImYCi4PN2ga/89O2xeLDgVKZcAq4FW28v53urNMOl7vdCH2g+bgjOsaeOYKlAuZiXx3RS6ym1
RbOgUwwhdRtW8kPMEsAUvkaHh+eXuV4NzYv7AYJAIhjd0Hvd6l6OK4sQ1USuEBJCgksp0krvDbWI
diPLMl+tR4nLT45H9AVig/82RYU6C9jHWmbEQQrJ2h6XmF5PH0JskTZ1VXVrsR7CXcaN74eelyyd
HFQfKQ/Kbq+cCqp+dX7RCbBQBSlzE+H4L8FzI9HoJXmEJ7w8iPYkb5PNohNKgPk1LNVT6hQ6rYkH
WMITIs+5ui4H9FSr9U1ZYYWlpCFYfZ7kmVCXyigI4iOGh/Jv7tC1C6o/Spv71A3kbu7M3d5M3nLC
B105MfSjubKCzPmlxrdLgW/s6IZhlNdkCC8GgigOdVuptXDml/MbqKuiyoTfk/fliwSUhQ7pbg5q
IZAl8uIeawcBPyvCsC3ZwztVyHHmXgow27d380Vr4NFWJ95cbbJ3bbHynZi0XDEA6O11HuIQqGxq
2SCb6QKlI4v6flP/7Uwbf3hnrIaGf3dn3TGONn0FbWMoASN8qZnGxCKHWnxEgEFDIFzftOqyV5jt
TWJb22iAXnPm6lZz1zc+PEIacoY+CiXVztCzdZKIsyO+KiA0tSTQOugRrqZ7byg7yf90m5Rp28/t
/hAJnXNCmdwS3I2hIECvrbYEL38919Nx9r6GJ8O70ZlqvZvc8r7hOcFQINIqBpH2T47UGag+8b0B
/MK/vlt6LRhmH63LraKE28OL0aa57t8NteqEkf3qazcXu3Msp1RL5hBFUX2TuYAWtD1V1prNDkol
chvtuD2ljIB2/gZQy2d/VA7t3Ez916wQR/noFsuDYZLg7JpLS+EbLLdQSXI5CFxaDB62Z0pCYGLH
tN4i1RrRo5GBNsdtZtUXNe2Xi63rxueu6Wwc8VF6TkME6wtWQ1fGw7PPMkMPUeP0HUlsz5kiwTWs
MEa1cEB9id3RfZ13+cnE6opdqhh8pvCBqonAcWwvxv35zDUMM2YNiBYXkQwKrU6VDIGWQAMLgAy1
DP5rI/2XS47du22FmeRyVCskdiriIfZ1eBQBa9YaHwFj6YJFyplYWir42Ii1QbFRLQ9v1x9CP2FI
P3ieVxKWd2iefe4HbrI4SjOcBWrDLySzuKPs4b+PgcR/o/OYX1pxf3CWauH75Qc7ol0gDTZ5lKdk
YDmzJbv/JFxdZyvcQvVcTNC2fEFVewJHGnpWQY+pGPwHbpF0U2WFqn5HO0ISQeJVj/RdDPHzO/Pp
31CYxZ9OwBE2cAti+LuzFDunH+Xeac62wXy3vSUotbk6ypYTIOaRARu9y+mReuK1u3ai9QnTaVNi
c+oHUJ+7QfT5zMd6he5rtabt06GuFtxBHfwe+CmBLWdNAQTb0yZgiau6K9JljQSme6Eua1e69DJX
LvRYmjFqMP3uLGsw7rcaht7qq6Pk5Ju90805LZs7sJmqsU2vaKMA8O30t82lsCchuIEJuu68tk07
KZPGOxp/LGIYejH7JeNZe5hTAjsFwopzd7Z/zNHyFww21GuU0jkzggVu9KwyQ0QyVMIWPlTzUF0T
07q67CDOoupuTznYo0P4nNqrMHtgiybWMmXPcV4b4biSPPEVd9GuJfpHgkIMorvHFFgSBXrckCic
BaUETR5EuB8+0QqpFeWFNMygQXqMXYZCikSBc7uOQAepzHuD80TLWlNJ85xkVn/HtOtQeMn0P1Is
YvuFJSbBBb3rQSwOD4WlgoAQ2Q6c/Rb5En+qUGXH9auIuheG3oqHrX8Q9HN3NvEzjwv0znVLyIQ1
leOvTzj+iDHFwkRrQ17FH1xW+5sYEy9t+NC4dpfxEj+fTb0V68WnMSXfs9X7Bju6XIwhSHBp2hSv
eN+348HXFKXJ4e2NUSebbuYay3aE0WDIXHN481VcmPbikNKk2fForRuuA8tMYt7gECPSsFz0UtXG
usTPnGbyKazrUCHExFZay/5PpXgyY9WMhKp6CXTlnQiOCjdUsr0u0QHm5cqJ39Nxfvh/0r35iMjk
7FYAiurvR/lP+d4rImjyBxtzSFhC2dLiOFiMB+3936gaVcJ7a1f0VBoZ7NL5zrlQTgcuhHR+6qLn
rVmSiy7z++MESj9qXHn43NQtPb3jpDLH9uVsNyZ8O7wjL7F048PaejFkrpgycaQDyoiSg8CVa2Y2
fzTxzJuLqKdopedvLGnwLAm7H8z2VmbPUnNKRMzDq0bwjvAyjINoaookOrZ8+W4DmUeYh3T6RV0Q
lzu64a8a35IJzc2Hm1nJieHg2lngUs3eesCRkWDQR30enHX5pEk9s/36ckqJZm5J90sdyENLTxvx
9DAgaD7vxecs0n8edaEB7rOgAmpihEBcGdkWyLp2387PjvUyl/VsyKyxcSb1RVt7oZg4L2I7LNMa
r+/CgY0uiRchgpQgfXOgwL4MQWeN1VmZrDz+XZCzouJtV5WJvY6N0zwbIXa/yTp0aVSza77CRP2z
QQkeCDBXst+FwKQFvmlfvaWe+tiWTwgq4/B8XP1tKZyaMBQjg20ksnkKdpnMRERMFhPS4UAfUyix
AvRZEjisAAxK0yLHRkt22nZJ1EJUKNsgoHmgB7poqgtIEHXMkrkbUw0GO6JtxcCnJMSKPncnlOtj
xl6cVfzIJw9LuLSlqCAYEjfu6aAqbmYot1rO7uonQ9l+47Q4JBScMzjHkL3jB1Ok7HPzB4GcUExa
E+gyQDxRV3vKADEbbggyArLrjlwEcy7Y589CZ98RS9eYsZlJIYKfIkRa2GMoJbNOmP4jM0dEkjaB
LkNUqYouSHG12E2Z+DWCmwP0AxzoZOuXDYW2NoSihxDnS4znhoF0jeUmRru+jN/Hc9vjCk17DGeq
0C/6q4hIcwiAsjmnOa7Buf9qsKVoYsITWxTHOY+57eJQysQaJ1w8jk+ptHIu5qlxz0Fr3uLNja/C
OMgvvOq5AOyq7a/7k/f+57+dAUFeykIJFyk6WcHteLRTmj6Wq3C3NVzsVG7RgHrbdbalmj1v9v7p
JIz14mZm31GhxoVXNOL8ngtOQePrI+NPnOTrxsncrEil/uuzGvR+N/mv/IEU32mUH2AAJqriRBms
qipgSUPHM9bBYZJaWiahQ4EYj9bVfrIXESX9+dF3FBXgdAPIJrt9JlVthqdaG+nHmTtdA7FBh7+0
vekb1Nv1h5uD+mdeMQiM8wdfZ30nymr5N7D9WAGvvUBg5w587d5M4FnbA8RLgIYjuOK46To6Q4nO
Cxljw/A3p7ajzdi0CRohkFIAWc+1g1hQfKyfh88b+f0KwckuNvnPPtQVVcDpnpNRBrk6qioe8/Ho
yQg0niVJTOUFo2lwvap2zm/MOPSNMv+2gkjR+08NjQ6Tc3QTStx8W1AtflsQ1pCbyWJrQrgiIChJ
K6p0f8uyZ6bPCvbO6FkSZuZVN5Gwiu9CPjeTw/Z+FDDxtWji5APVZiGVg9nL6mga1SiPo+crcIew
9HuJ3TEnu2Sc2FwMSH5+4lAs7yryvMgbxGY7uxxEKxskaIq17/Lg9WwJgtjrLEWfG5B+FWY2v/o9
Vq2DKZNo1qtUEFULL5O7uUWmgnpXPttJeaeUebX1WwySelPxb1LoJ5HjW/DAUg0CoUc1I2ppjVnB
0AIOoTvuJT8FYTM5XlD96jEZBJGIjwoLR/fY+GhtnAixVaa8V41VpJufbZOSiX3xiBv5Cxy5AYNv
Og67haA2F3rRGcj4z3eBgSu35SsUl0If4OtEtlJ19kKaYkBj7esFRADCqcd/B2n9Vd4nKcFXhz4R
9ERvf7OV1yhBLv+OPUY827NAlstYIWBVph3khk8710ggUSgUEmycEuQHDO0+6WlhnQal++l8DUag
9KL4mUmv8nWyH33g7Kmcf38LPpwQMXWswq6JnIlvnZyONt7wcs5EQaP43C/GJfRISjetL88sYXM7
NRC1zXfcz2lp0ZIrOSd/uRbSAnh28y4rq01DIS1ksbnzfJNQoqQPUL/2bWYJ28jM5aIIhcxQiJgl
eDtntBbEPrBhIPRPmB3OhUXjcJZqnDozFJ1088dDeQOz1WkOx2G9C5SZkXQv74glyZ1FruhvK+Qo
sFMQQeHDdqiCmhAhtLHjZJ4IqADEdWD5zFUfxbLwdJOg85FTGJLj5T0R98cQ/iFu3YOUvHHyH0jO
3vLSlTuckM8cJwMmHWsC6BajD4955R3/WrZyLAJFtyDKVApMCBcAx//zfnPt4XGghrKtVsE68Xta
lpmwud5fiscQ86XQqzC/gA/MlFfssiLDOFvUQnaWzk6y3CVVKq5536su2GNcNeXc+7+E8XnYtsnz
i3DaK8vnzC6DNHSZu9TjZlqIMF6ksRMsAhiT4VmxuTAHQAhMHQMyMsdv3VO/fc8AJTMhS3OObFQl
E8NMvdkC8GFx+qdfQUlWZu/Itsc/Ks5+EHvBU+TnL+M9OMBdT4rN9gHhyJbyrSYL+CuiAFdR9Ixu
ca3272RqTEfhSUhZdDo+ZDZ5q73q6wGkQY456HHLJ1m5dOul7zayyfF2+H4WQrd78jdU+yWhjm7p
ImdeLr8AtOJkq+iG/TFr8hcS7soCXXX9690HNOp+idmlcjjJ4flUWjcFf4hIkzetSprHfkXd54kT
PB14UYDpo3OOOsLMAu6M3voLkTVIwkiOsJ2sxZD7Z8g9vIqmPxnHN6r8AWtz8Cay9ccdH+gegyeX
zucYLCaz9NyX2ffV8/WNfacUDe+tblc5EkohnsMxvqSSzUiMW9VFVyEzKFjezXi5ZBUX6+eXuUgZ
a0J/67BKtJtihO0lLhUGrj+tQ9TcMmQIWjIsnbJXp7lrcqSya2XbB8j1MnjROju7bHYhemOuX2h3
7aJq4AyTvu0enlt+U2zkk9FjfdLMUcw4PAt2vQKlC8BIHwbzLUqV4v1Xg+DNvLV9ktj3u0HRWxBK
f2XkCD6zJ908uxbfuRnIEJF6g/NsxCOlXgyGkKtRjtRC7Fe2OXTRXkPtr2M8gJxL7UT34yjOc1dY
kHu+k7tmrZLoynlgBaIiIDLLB0K/HQYtH20kQvcW6bFyNESIOS+JEYLGpZLax4yoJiaN7WzSXN5M
YeBKoH08UsEQtAK4HAh1r/a1ulNZk0mZtfb5pQlYHnvAGJH+yjquu+rZ5bA/6pb5EBpHoSMrZ6fa
boGI16u7d7UzMAlyiS0vOQ8TDesTofmj/f8cf1DMUVfss0TQrd4mOsOqfqCxT5Rx0DS5dEhfooJU
IC2WKe8zxBZ0Krgi8KboVLZOkNAMjNZVeRQBWtwZ3yy1M+wrmwhROkCTgVM+bXJIQLh4ePYW4rk1
qd5TGzqhHcJc/Rq7TO6Nj219f2NaRETFrAkwXxG2WrV1kaWFNyitniB8jk0ou8oWyQ+TVHyvf4SI
BMIJHJsRx95SG/iEbdidqLk9yuOchO1rInIKO8nQ5VHs2HRDZCi+0pRBcT9mXuQDZypw7o/kc2Qu
Kg/jaKgMgmlPHtRdzDpKTVoXufl9y8Vuq0rGA8uGUiGiW+zzWxYiTKQ/QaLuZLUwu+hlI+REBMxa
fzl+hArmACVmnE7Y4F+prJfJo4CEfOS322iK6ljdlzM/o38z0cxRhCK4W+e3hIn//I30hkDvWMrf
/1spdUDgq17F5Off6s38NV04asBRm+GNUBXKrFh904Gj1idcDUexTmrnCoL+zXaQ+NbV4XjCggj8
qSWFr0bKP4MtcJmiVoKDdFXc3y45dv0NC6tJBRuLJr8g2wSx5i3mU7KPwD3Jx2AbM6P6epX3Fd/H
t3qgsRpc4W5E8sHmFkAVr0IWysC3f90q7vRphSytgfmr9Z8wk8ZcLYGehr3zJH7302kIdM6Os8xF
7fr0L7Nmdnq+ZTkI/Kha289MnqI9WBE/gNZ2TUi1bSvR3+02wTPUGc3Ie7dYDa7jykV5pwXFLoci
Oi012lNQ4YcDn+JmhcHdQ9vjpkN4JnMCIPfAx4WW7pP8BUX5jE5em3je6x7ux1RINTkh7ARc+qLM
+kBB0KZEkKbEoBAgrB31Wg6pT2CFEMFvxJNkgE5BDKCyPr+99Pr0tleuLZ4dNjl9ch2u+Fa4QCzN
lNi3GI7gte5m8YUKSok3yTa5kJUzEvgYqs0S2Ay7Hd6elQn09k/abk9/L3hgUR5FvScEFbhfc/Q2
PlZ4w43CHZjIEn/NzQ5CKcoYt2T5GMLjkzkJAc3FNKImJwU/fCB0TzF1+R4QQ74N6Sdxm9rIwhrX
iNmVuyOXaxDrOf6UGVKkIRvEf9tW1mpv/iOBgvlEEnMUxEm7+BochwT+DgypWVMUTGPlWv8YoF0y
WbHdJ9i6tQ5xUfpHcLtkRCTYsj7bCg4covXLKC4exd2hS052qeU9YeuT3f1RDjbBGcy5dWYwsBqq
hkurX0AVsWqMSbcroP/C09vGDuiLXuGh/JE0Ww1y8QET1AIF7R7q6SH+wc/g9PzwDhDdJuE5dJhD
3gCgll/HOgxk+3fZo3+qJVT4+7Xc4/rAsMpbgDGVSAbt37fCzHjx/Xanjjs2gjaAgrFNzvM540oI
zOxI+TUKvQWh0K61iB+hgUlRJ8jHZLUndaX/mVmFcxuevf8Z2CfTpRB8YWYIY52ykz5OBGkc8XLc
eyOd71LnD1xFrWZwE9p4PR8l3jZ5h8l+CSWf18rE6+1aHSe9wjWYvY+NSqp+km3Uqk+1/RhwdRCz
CbK1b9C/0OrrnurkBpyPzKkIDoeNqgMoM6xwkCw0xox2yo9h/INKWpg1TeQajDrUY+6Agvu5Km4B
EXzXG55SKt6KyhlrF4GRcspFdwZG560YeAFlgg6gqfPQI0ow+eXmVMqo4pNAvhh1BzPktnAF5wCN
dbskgFnytdkiFTZWLOBGF94OJa3ClA1t2tlHvI54MAjypJuCpkjHa/azHr8uNV0fYBe7XDNLeOfp
oWOUaAJmvGTRWh5kLVAH4TFWMGbznmt0yjdiMZDpB4k8jqc9FqEhz4noSvgr+xmwNmZaSX3mT8ck
tYc+YQKXkrZeySjLpOceBMDOpZd1Tqcitewp4KS2c/Bihc5Xk0jUZJ+w3KgO7pX0SL8Odbd48Cxh
nr8/jb9/T6Htb/IN4K1HrtqLR82Yucc5Km96Mkd0dmkrbYCGHt75c5Cc/VZcbmGy4JcgxpAxYkBb
kJHlSyQiqAwAeb7zITFH87r66LF+gEb5arMPDMvxk9kdbByrKA0QSp8RCIdxD7G427YloPaKwhBI
a44kbiXPPsYbMZrBPbiGmulzBsJ8Qcb0rkwEBTUU34RhxyaR/JPA7AY/SerYXmTGFs9vyziZOK0N
zDI5a94jwdjdqNLega3xVm4WpIgHfCgqvtQZwI2QU4HlPleDNbsKJFy06V6q8AeD1S0208pHoqHz
7OBqVAtgu/6WmjzRaO8+KjMrU9WZ3Sm4+eSVSvEB712+4tLKOmMjDU5Lffh3yqKrErfFw6WLuZbj
uxzmuXpXK+Fiqx63R48Bc+zenBREtm2S4frPl5a2r4n/lUyZWemN4ozMDbxLQt2wKT3nbsVu80Ge
EQKxE/DMQ3kRLkhGFsFxIP5ld99N8Lgts3a3zluhDnAeFyBFqdTHg2viFmV/FgQtPYdR7ED3xuIu
vto0nqu4+WTZHa48hvz4N4BoPJaxPWX3uaMtEHfb6nQOS523FhvULyoomgedj3AFXZZbD2QBVXkS
6OjPtoQZvCt5pVI8Cy3YXjHFDGaDY/2vByIxm3WZYOaR65BOpD82qye4ovCwUQfUHHtdgfMm1x99
e+pfuQ53oY3ENBLfoVe6vU48xrs9VvJn7HfJNTtIqJqTYIX5Cu2viw9EOzkLJPlrosHFKwGYzWYh
SmQNTWJIFzLjwFthq0hdC7hBS/X21KzshdVElYhBP3L6YvPtyGXDUiFH79iak4bRKlCovh8XBsVt
eLTpy+b3ocIgHLA+uoGGXTOk0wSLy1O6ijOGFkccA88ZkzMc+ZSIY2YT7c8CjRxiMVrZ/EUnOG85
ghA+4Sv0SuZP9CTeYL0pRFl8RQ1YeX5+j2AeJJ6y/qC+4ZfSdAWZkTsqwkKVvoHPL8wMfvRWe/Tq
frSDn82xuWMJSpSEV5sMQGPf+zU/rFsTFP3u5MvR/51dM/hIWX6fPV6Gexmb2x//e8yl2DVGLcQA
4tsboDfvH14UBOyBkUwSUa6IjvlMDeFSJJ7XYU2EOY0LPrBlZahyDNI7bJ5BIVOGfrPMBistQpBI
Db5Snmk+JUXAtYBKpflKHwDbT7fD2QYv4H2YwqyEGzd080P3DSJma5I1zvzSuZKdjsgxm1jYk3NN
GFDVxEHpWYkavAaMhSssgJEKEIgdOOljx9nhSShrPRn9vxXScL1qKWlmel1mu+3QNrhTHPaoLd46
WtD0GtuRRjphej0hpz28Eiyse83VvYkY2DKwpvGmzo7ECVexMAPv2CUpclyK9CFVU481XYZ/K2WS
Wny3XB5q9p+INrFJqxZ63hBShG8NBVdUv1bXNKZ9ww+blOjEi1YwWuNUl4oJh3k5qC++JpLjNSdi
B7+G8HbjSuCeZfXxGbvEvHcXfuqP5hnUuyxmYCxHj1vGSFtKuiCLfL1mrsBUv3M0D4JvKRilIdTs
IP4kFByqlrz8HXrqR5HhuNbQVGC/5DORoYEXvYHZ/0Vr/CalJT7wSn4ykJOU0hBzzjAlts+3p6R+
osJGRf/WNpDx5c0RA2QgIAeoqQgFVxCU4f9ZUBm/oTg7HEbJ0clGHbb4q/SlgpEin5tYRrkME42O
F/FX2j1GL6FseKQdHognJCr5pZr6X5f/1ejr/BI0gy+U4ph5ICxsBdDrcf8MyW3JamHPAP1vywGW
UKrRD2OGWDR9fBBMjhLVEC3x+lKNNKdPjN4fRartZdq3mzaZae81i3doBcm8jjwzJ9nDrpsRCQIw
qh4WFE63Y6oF/92zQqqLwm43SptjcZkvol2A0KE0NyMtFr+i2dwkYyCWn0Jz16yqgpVQB7cA52VQ
+1HxToZLRpJK8EGB88/cyg5TzHC/LEWe+SIVJ0b9lpBceoMkYknLlQKSvLQ/UWgnmwQlXyI36Arp
FXPQV9JnA3H45pVUxUZZj259FhHPoR1UJw9hNhZMUsvA5f/B3A69K/T5UYBNmPaMQVoqtYKepKNi
bpBJ2Fer+JyIiHjx/HjxhWYKTh4g6u833X2tc76etgyz6M3fcBgOIlUgVyiSPdULpFIIl1cvPrSi
LH0Q2oguGrPNxVHiKrRtR5g8LOIk9Aa0bfHzhai330A7pGBp/2Pa5r89V2lBqdnioRIkTthCwMA3
pzIIwn9EZr+cREYNX/1X2G3Zuie2Ab2G09d04iazxDjtvfdbl60J7vqDoAjC8h9Id7uzlfhnIT7O
MoTAkGSJ4nFVZAIFMG2geEqaWH5txw5oyvO4gzVANZKk7R5sCN9TWCD6MxSJI1IBNhhQdrpLBoQT
ZughNZ/Z40gh4uGtnV8NIAUV1g3au/7o0Ndbol+qB1QOxbwV8PlmLFRlpt6xQXvxuoFG0AqixAaH
W1dpxxN7AbrID8Lg+rDr01ZvqvVzqik3fMD8APaKviRp0VGUlOt8W3sX+dfbu/hX1crGxYAwx+Uh
ws+lAoxU6LpkKCQHPs6bUW5OSwqMTI+k388KNWGs/OC8FY0f2HFE1sTTDKfhRMW02BJqdxa7O8b0
K8pSkME8xQXomLxBx4fSyAiC0/nddKXTIB6qw3qVrzQBrzW5VfmbfyCYyA2tkjYjZBY+tq42ligF
ywOX2DE2Ifg+8HlbGs5awlvsO1fudk8CSguJMWhSwjO3ey00k45IM0CFkC7webSI7uuxgOs35ENi
zU5p+mBTIcqVXCjXPbxppXY5uG+99lN5vwJ0j7f3SOgrCUzVosjdfSuie8+Co72SbWQUiu/zjZhg
R16NHswaE27J9Vb8MjQxkobfzoy3d6luwG3I9jlEFVAb95tPsK7A0qTOws9COnigIgcMeR6zvK6O
7HW+vD9EvbppJ9AbdRBGG741zPQW7pwSVLmVnW6r5+DyIWKOUknXcN6p18tjAeun1yRi7ZrlSHts
rODXrQBLUigrfaiiVxjxYwS2mEidocUCeGLPEgX3UXT7/ePy2L2SqBUW3U4imfVcq1cDUQadxaO0
bT1lD7hDUM2dulHNfaPI+/0wkbi4YF1P0GYtxnog+YEhJZtIOPBmyis+rdNtpdvFEa66l/cDf9g/
5bGKHYBPPNzfeITXvoG0r08Imej1fogJHl9SOHPvMZNrXed/UlR6iqnydvkFrC8u7FiratL9hlhJ
3gcKrbE8glExNizs85E2UHcWdxqSIQEctBKkvj02Nb+Bu8qVbDaca15yOJRCJSmwaFEuy7kCKhnY
BcAhd5HZO3qcM1FOLoYEZ63uShgTscvv/UBDhmCj01yxUBNfRk9Tpk6f/xHt8StuMnAQXDqQrDs5
tUckywbqrYiG125qPXp3KIIjiDyjsKrzeVxdMtu06ardFwavDA5qPDIt9bj60roeEN9POrtcr5ze
X8V1al569DSUSrS3O32crDVo377ax9jH9aCMfT2do8x0lDIXNpoTJ507MUrKgdvxAcpSe+n1Gdap
YtxwkdhcMLr1no5ZTwob+5ffoSl1kWhZgXbMrkQGWn/WG/lhhWNHNNUg+53bR9fvagkesaulGIDu
+Hq/zzQEEgEuCs0N4brLn058F33OQcFb6G/D3U7v8Ki5QbHrMDnJcOCS1rBZu7IRgpF9W42NewbI
ZluhvINElqrJyjkIwRrwJ7c3COOo2yGG2GGj0mZSGslI+VcaJGvVs27DPbDbChfns5u7STaJsaN8
+dSWVLfJq/lNC7H0WDreWxv1u6kuOUc/MMzwJelV1KTaf9MNcV2yOcWLyr+7ipTeohePrO6jF7D5
gsyBu9kDcBqfENJ2VYNNLNA8l3O181rZkabqzbseXeCst6ieJyYRcb+cqpH/niAFx0+oy9v9weoV
mcH2NaLV4DUYS7CNSkfVzbgeGv4DWYB0tyOk6QUklSnyRHPJK5QfmEUbWVsuYoh53Dy5KdRWBon9
Dldnj0nOLdCjLioHmaIvITolCG0InvgwfSGEbsiMsxggwvgQNh7ZGELtl4Bscl5svdooWuN0v66K
nAiIKCZPiiV8/ecTiL6dYjvFfbl6veJt2BeUTfcC00V6S8tkrPHR1XFBffK+lVAnXoz8d1q3Yo06
UAkLEWuV/Xa1to904hXxrvNQnEa1mtSm/7bwIYD4/wbuUXJdsHZS8wTMjLybt9dCKn4RREuBLFPY
cWdTyjRAllEVHyAwlg/7aHl4JxdaM3pKYAFAZzhb0Nq6cfmukl7UdS3sZCGTraQ4M2oJp6x7bDTE
aCCj/RlzP65Z9guo8OGmbpFe9s/sHLdPNUq0oFM4f8aHEeA9Wp5WW2jDlRXNq/FBSFKtlLbzjdqV
/lSAcjf2uSIZaGVMpuEcJzVOYpN1Av0jyn+18VnlZ8gHcX0ezdzwYNbIvQ0fOjXTa5FH+t1HxJVT
ie6e2AcIc+SXBrAU4ltCzWu6NuPDCT8X/u6sixIZfV+ttvRzav6z5QGHz8axU+bonszhSMafilrC
APt8awuOh45+HnOy8ameI3XRgij95FS6lq7sf39e4tywZBhISaotWRpwLxvriz0nze7DHlag3/yp
i5vPT82Phl2D8aDooo+MQFF4LENpOipA5FrKKsPCAY9tgchNc+68RhAyjfI1AWqwsy6Oe9vRXPr0
/0Gcoz9EpI6FJS55NIUJXXptQFXM+x4EMxWt1H4pZEpEpYDHAB4yuR9ROs+aNAHe/Ptn+cf+RH2f
HT8rEzBOTGt+tYgu3yx0fGc7dXkgVzw0X99TIQjx3jKlmwnkADp6bMCBJc11HUIkbJo1+5F6kGWv
mebEQk+u+4TJwKE2jk78wzkE0FMDvsMWd/sKEdoa/LAc2M4CR78cvYp3jhw/44pgbwDEQyapINWE
WQk0hWn1K56SzjKCeh8cKAHi0U5zs2OjWaL0XqXBIvkudZmcKeEsymUhr+B4YkGS6eRxdiR9K1Fc
STimS17Y9FapPywsonOiYopunGqWhT7pLdRDKjVbEkS67yLdgORb2RYowVcVuAxsK/nbjyZMbL1Z
gf1pEpdITC0folq8VIhPaI714iQMAP9YdBAKoaAh3M350Ws44NQ8iUQsDOKUG6dNivO/GqGqZgE6
/sj/nKcYwK+5h9maWZJ2VUmqRGNW26lpJLGHc16D49jV5xpoV0xdsMVYnLxLlmYa+aeEsC7IM9ig
UjyOLVqHJWevflErsnaIKepCUJgKTrbhRPFzg3oFFYnqHwfrsK1SBti1ZIioO7eZ7QvZDux605v4
YUUmOaufHMWDNr/wZSp/kwTxeNj++sQaVDk885lk60Q8xjwsE+k70RK4ZrIQNPvFEFTBtjpqdyAt
UV0RQGGSMUmiFX5k7JZaln5nZH9Wv+5FEd+a1JfVBZMyrn1cjfJen7bWQGRhd1c90ntKMRH0Us9w
YwbyEis0WdhcgnL/FqfWn9fC6xSfugoh4mWyZMXuSgtSnmJgVgonVqgR9r6HY+ZwfX4jcitDdihu
1Q+qfMMc7+vgZI8G41y5KfTxRwLxrXEAl4oi4vvHJy1Vir0G/PrcArIwZN/sO7tGfDB9rLW67Z4r
ieCkd4EVFHyuQZQNr25YYL11xajtcf8C4j0alj5XoSzpDqAfVP4YpJhVsbmkLBS+hb1TUXv8TE18
uPR0D60GFAxfFRtacaWtDgOiJwdZyF8nS+3HSHW0OrLXZIeWIOJcFcFPyv5BRM2J1ffATcAf73/h
yd8WjcjboTmEtN2XKnnPk0/Lk71HrA1rVFqhlyMnFR9DiazIS+iBYMu1nKxJ4A4MFClCQk47DBVC
RNdRHBVDe8mgLkuMKJtCo6niGyseb1sjpVl+wKvsdz38NmM/VP7D80lOINPv1Sq7FHfrYAt3LuhV
+6KapfK3iEuu3VRwj1HFQJ2XOVWHlaeafhjwmj57va3OAmLGPvmjIit4CjTnotqtWjh5hJcv8YgH
28QYQTJc7fHCnL+6r+0eM/C3ZyneIXd5vvvR5Yr6Uls6ffXmE6RcjNTKUpMQOQbjji7xMvFfOXjF
FmepP2X12m8juORySMvMEhzb6NLVdaHMjCogs0XlGEhJS5b0j+ZsSmBaCxlnuwjq9x70/6EdAcbf
EmCesJr/RHCK7bcsUSsPjfGbYj7GW5i93/HdSjBRrZKJrHJZwsNC7UmkF1lIBdOkx+b+vaHiWSPN
0JnB3d7INRJ1N2iC5uPepw83Rq9Q2waV1BtLHAp7z3PhO2WH1lLpUK3SXdQFLNjS92VQfbGjDE6X
oOQSe+RcnghiTixVbim6v5JltWMiqKVUa5sunp46J8hLCPS3P9ydR3YxewvxL7k6k7h2lsee0SmO
ITr8UlnvSMauM4uMXGkP4iQmf+ExAeucpbpWrpkpJZ/vml9iZrvhMtgKUhoVGS2CS6w9xLm8qxxK
+ID7r6yfBWcDeL+o/Oa3gaxtB67kzluuxQcmUmypD3DMqVK+rK5Vp9zkGEU33ic8tuH0GbGUt1Ty
pWvCJQuKprJXeClxSFa/YJiWtL8vqJWg4FRAoEInpiC+sS9JKrTiCoaHdQMP3OaXsCgOMpjIBHj9
iIkPyFFV+P1E0MGbRwyQXx9i1j4f2tTWeACYXd93J67uZR4OTj5M/3ytxU+89CaJOEZtqkiYnY1U
/5thn+IDimEdSXpotjJuO70Yh60B3mY4MZvWOqBjlbW4ydXXeSJscZxbq5HA4Zi+uPzJFux8NESF
Hb4PzOqzbgDijTP6NXmHaXXmGR/UkRK76UO3cQJDamIiuygTvY6fN92mSgiobzUPAigDuh/EzBPF
Sz5suihQvfPJp4y9pMNO2zvSCltlTXY4+1sVlmRzpk/jDOP8MNi1fMlpemZ5jCZQOXKq4toWaqNf
VMUva0ukwXc8rdLfk4EkVZmtoyHKtgkCUz3UKdxhO/JOPCj+qZhy5kgg2qSwL8ZA6dMIHpnyMgBX
IwlvMajhQVgHvnDvZN3PsQJDDIbcOeueHr6srV3wPpymtqq8Iz5e019kSGMmYG+tEZlsdacu4yKL
MBZd63RAT3nQJMGVOYO5qtOmHx1fVrYfkQ7KV02mSFMXI28EQKWjLJ9PgbOaHMkrEWhuORMIwG/9
gbVPnfpjJoCIMyPRkOMpEONDAvPxzmOgWqO9o4pbNQcnU/c102PpPLiUg6l7Srvk/uQerrjm/gmY
2q8qjqpL/TZzwcX0K0vkXHVOhi28ZEeVnFPBMmb5vJhDcV0bzgMIvw+TNpW/aA0g0KKLXsk+SXdo
BgZkURMICLBUVXSEohdrrQdy2wuS6l9Gn5TH8bPWAn/dPwwD6FQzbX3QoRxJHs8QK3I/qSA0JJgM
HEnvmC4S74qA1T8fftjpQPhCDpqyVnEaA+r3/aqhxyJUe+m/Q10KLg4+zDCzr0FoV6Ujunavx36C
VaMRNyEZee1SSyCCTz46vqTCJQrUglTDFDuex9+TQQtS7L+JCochqBFnuUDBvzsSERaqfU6gjjJG
KC6yhzvdYttiYmAMjLa63HewCRiCbwj23y1yq5/krnNnCkOwidKXwSyDp7JPwQ/K1KLUxu5MZWlQ
QNU8yffDbpSZq6+Rw6jNBVVJbc6QMDBeDgPKNnLPMNxm8O8Z1Pag0IxnegGUjKMY5NGUbtQYZEii
8d39PxzfQLorFvwqcrBEqa9lNPPKajl9vRTXi44Lqa7Hu6KutURRxJom8kkAHh4EZinsZ9/xfQ5v
0FPIx20GnsblcTLtRu8Aik6Y6g9/rRECocF28W6HxtMPQS0yclDS0Pw8XP/AgiHOaYBVQbG3yAar
3XYQNgk3CXkdQaiGuNenY8euymHGG6IWOrT3eTbsJJw/16QNwtCGpG1pmhE7XmvcFPnyAfhBuPpH
x1kWPQHDWPPnS5NanebTYiDE1enztRLGds0GrgkcC3ytZLVSgDDZbgNnK/QoECDOKGrHRcZbVUqq
wAQ1jduqLQrT1+AkMLKhvPscKYaXQXUc0sVoO1B6c5QsI6+uLsNRxkVhMbqm0nj9TnpJkHVVo8dt
2PvYdNfRZEcxQ6F2M9CC24TAbZAv7AGoiUzJYNhvxv9uptksfMkKhYXnwkiP+vTcxTHzj9DAhcgB
lukbCzVRPIsMld7sND0ddnSA4R70/+GyonEubkWlIF+6uB+mT3XXl2o3sN7F23JZB4iIvGDqS6Bw
9ALcNXhMG2dKR9f/LkbDTWfa9HGAxVZkUQfLZE0jbryRt5MjuFHPYYnkO1SP8PDUZSd/fUYvdewu
PJc/mqSYWMfByksF6oObD+9oRjUzPfrom0aExnPZylbYSC5hXJi+yUZBPaiWHHwTY/0eugQbdwtI
bqrOLJQHNaoDFAnptm9JvLLzeNToWAbiIVa8lQTSyAoAbfYvhYkyBx+6Zok7f1P0pMaNDowOnTV8
b16srBQvxSdqju5ShFZr3hkZTZkyLNaIwEGRTHrxue3ptqrzYwerNqAGNsNdut1gttPCSR0d6lOJ
FDPRiEdoXWZUGkyMtpyojoYN5GjTgXbL6biP5aEzsRHLOHXbNailDIu2bnUZeQlqsuQchN7rWH6t
PyV8xd8uVIYw61/4vNf1zsAfMiVJWtcq82M92vBJ6ptAm27926lm9VPYEYOd6+f+3LMPt6t12TzS
l6hXN3X/nYB6wr17KfJLxEuZKdtKd3jO833F52f5mknnKdbyM7GoVG/mfVu3wolZE50VooTG2eb/
UBuuc5QkPwgDLJICq+iGL/HroQvX8sHiQOYw26r8E3H+1vdWIps7r+1rmhhjnoJkcE1fcHx8IcEw
V4XPIn6nsgZj2INc1Gd6SGoYhNAUZdby7z3A3aY3F58rWGZqzwD89TPsrIn1ttzqiH7Ug/Ipsuq3
7ihvEaot4b1SlVlZETl9sTNe4j0/iwireA/rJBRw73SsorSIV1sBSB7a6KIx7n8+t2dvqVEpSPaN
VqKobDpQKXTO5De+jVSCO7tPYnEgGarMMpwWbaUySeBdN+hcNWQA04tsrXw+pmTf2D4mebYB4Hsc
NZ8vSx1jr619jGzs74oFhDoHqw/bbqTDkeIH2Y1iR9iJS5HCXKVdy9n73kGsW/Brdoa05udVb3cZ
fIOdBggVjfKuya2Nb3l1EyzhSXc7tZyi2A0F64IAK5eTIvDNWUuDEPie5mCDP9NMsCzIfm9OWwkH
MCHHOFB6BQPT9JBpYfHMxDgnD0z123YmAA3x5RcUObfcXJGQkyZkbp452TO55ulBf98GwunA6W00
qbIiSlVtiLiWMqA1X5qKTKkro9xPw1Lpp72UKrT7vXLKDv+e1Dx+4Nd6yFlyy6K7S5C5epuUlO2z
M+oPSN5yk3TIziIWwL1JJT2fY8hDjhkZnNpVc3pZ0wfRGETJXEgOllUYGgPNWnehSyRkn3+iUdnt
RsJv1G9MFEf+oHCfyhW/Q3Xn0ETgipby8mYgz+kTwu+sKTxlo6zRY+W92XCOM20hUBn6sANBC7SY
AUNLZ8HMo80DcaBPrSU/lzcZGtW1tamNTGj96H6IwrQV+ZlGKE/q55EhEUXEUJgysuoRF6Ex+049
B0b/8SRgf8UbhVLFFZGDUT2DctXnLEgQrSqlq7iDetVn5n5vV7PQ3Rbiph0r1dpwy+4dOQDkGXDB
N5qL4JRjTS0RGe4mr+96E5G5RvZqQHd12slpXgCQ6tQgWncIHNWB6/E7wstwpmWYkc0OGSzTZTHn
kk3jrrhJMg5QxYyBpOFgK2yotubXA4YAnifz/CyLSjEBIoG2qas2PqLBgTt8t6syXCg1fi8/k7/W
2qteyy7yfrioCVz5eRbKKb336JkLJ4GVaVmc2keqqxJiTrjhIBI9wCME3kOdGKoxmm+uO/ViSjUA
UObjXoTvgaAdZiz+rEPSStvqzEwiR+A/ado4cBTiS9Adq8IUp2X5ZQjHRUXg+Rl7vDVuR0O+f57z
VCvrSjR0P+AiE8/C1DU7YzcCgVSbQImA3BlA4OPH+bzjk0mT57ih5zkv5v61MQsRyelDfPS4K30h
sDEqSaXHKCXsjp5uqCjKZkI7EBmAVzX6reXJ0Z1M+7G8Y64w5ku9SYO2AucOvnxzEi5V8YBBB1c6
LIIs5mQTmmbpKDaS9ygVH/IWxS+eue5gfu/+7q0z6K0uczkUL3e4aczWzvcXkWosN/DqlFdeevnP
FRJk4yoJEVCZXvTHGN6Jhl+6qMTbt3O50YROb1HiqFpoaiZ90gYE3g2KCVY1qvAKkdwN6t88UUsP
lP2Zd653SOB6b6VYt/JVU/KU7tajSgrgDEfUlRKA1E3N9pxm7SizU2zxjNdFyk54CHIgiYGJhNrZ
5TQrbfxnvj+m6cBtD7reyTwfYPJYALr9zAl0B5PilpEmvTuA2ls3RFRPiFTIThYUGJIWrWwK+Mpi
GK+6Zf7kAFoFJN5gS8U5M3Di2bJFUk2q4jBPlvq3N3QrEV2fDkGpq8MngItAS2EKSPzUu+huTv45
o/ygNbTTu/zw125iRkYf0pTh0hodk58TftwCWzxhFIbg12BOAnM11t3uO4usc2EQtWSolRV/bvp9
efN1e3VEopK9TbcM1AB1MOpuIGmAeliG2Nw4c3nnqVTPgc5bBIvhAhZkK4NTz/WIpoRePc4TaqQW
xKjqEexf0ss4qfEuPcJJ7F8mkpqZSK6aNaSuGB8KnlQVNQTZjWR4bCHTNyQjFOXVSfqAD6ttIfoh
E1tKePvls72LLZYRZgMGDfbv4Iufgt5nxRSiOZyjlWEnyoWdRXwMXMq35yCYiY6Czcm+X0YzhI3x
PxY17EZNdXXA+o53z5/VgZnYgJWJLiTkFmbsPWjrheGQyMLW1iaDDbZm+GPjscre5lHIqMfxrvNc
UaLleAa1oZRs0VWp6eHo6n6zY3xkTBQXYsH6hGFyv4W6OTMtmWV+W0OdfDIPXBmDZXSTZTvQlpdR
SVVgYIPnzB4dNT7ZSScdrQFJSjqvmmw2KsU92y4abSPLE14zc9RL0/82QpmqdZqQzd7lWtva01n2
Ijg9lXtLty6QnU2Lfxxu954voxKq/b/+glWm+t6HDhcJdgu7rr+i8GORL/6AFuC0678KLJsqLbYd
dTcGXCSNPLuR7CaQI9k6xmHg0gaTGKlDS4oYpdP/gfuLF9NVrTLKs536U2Pi7Uko3Eq8xRvsyAhz
vIaZisdPM2D7FeIFdg4Z865daK+ckrcs4G6H/MDaw7OMdgX0rQpMqqKQ/QqFnNKlf3QeY9rEdiH9
wImVTllGCGzX3sMymtYrGaNCPYqSzywzovkmYjJH2hVCoTX835PWI39tGuCCyWvgsRR8k9Yj4Rpa
GsFdbGutN+u/ws3NKbBhOTEKboPF/qVd70XwuDHZGIpEbpXK36DkTThrHZ6quOknzxs2YIYWDuLO
ksVacuC69ts8ZSya/LRTUIszKP7zafHKCZaiYZVnQCDyk1zXc0bebWkR9e4S2tKf+iGHHF+HAOnz
omKt3W0/zkPV+epbQbDaYIK9NgMm6J3XtGCNLEYGDHM2AB7onis8MlHMPYCpkV7q1ONdzAtedgAp
n9Ir/vIwZ5xaUdoiI07lec6s7f22BTYlvRbVygwvuF8Cr748B0p4hNuOxBvGg53/w8vh76shBW0I
nZXy9cvL1MF+wLycslKyQSPcU255kMRZtVvfaQcdzomNd4XeowVPu3K4yMr0y0rBBfVgMmxqjaF9
X8B1gA8nyCFjtHgu6lBaQFD9AbaRGoHEteGhcmpWqQHyyUoj/ZXlCad0UuJs/96YPiW9ztkLnfX8
svj9ozdnTwxmxJ3NtSZoq4nOjDfxnq7Qb2gs/C9tSWyOcXz1cH+oq5j31xjG/4beCDTUY9N8LLF8
Bs/3G8esXDj//xKb2OpvzV9mgQnjBgGz8DFSzfUqBsXypxkYHk/LMqAT27Vocrc+rgu5DTvDIpwU
QJBXiPeUA5IS13BBwLG8fSFbZq+2p7WLrew4l7mjgzF8gJnY3hNKKzdg26TfVMgpB/Aoo0g5QC/a
vruZY5YzesgxYdPg9SqLBG3WWtx1uz8+S4J8dyXmQo6oX1XesXlgDlCDDRLHfiNeFLJBYd4zlCs3
o3ApO0LrHpN2KdIUR84daCLAFuIP1c3KHc4tPGvQ9uVZ9VHIjM8W1oMO3UsPXoDse6LySt8KkkFz
NTB/GA4CwaouJoio0P/TpNoI24zC5NIhq6BMVGG2GXaoVHQtnCpshr9qTRbz7fQkfwdTYTzXQTdV
7jHkByT7HxbsdEpdcvLhPPkpwY3zA97IS598Ka4vwERWuST7Dpg+O5SlBHszNZylmvB7bFClBgvh
xNfzgJU3oEM/ZMfBSlE6v28yPIhMjkMTDthlX7bdYvWLmfNLhVZNYh227VjtEqktM8kF3ABkqU/y
z+I88d2yaGetf6bmn2mcV0P8+XeiqIsCKLouRCPiOouj7GmPT1RHNVipGhZrlqw07p4bpL5ZzS5/
Qeq8c7F2qRVylZPTTj3C5gYYIc89SsaP1igdZp/L125yV4Qkd2X47SHMe8EdftojvQxqUYP1lead
lmC5kCg3Rvd3R4z2fxwkUnIAiLEUIf52TIBvTWXjRS20ZRlxm+edXCQuvyVu1MHP4bskbJAGqQYn
N2cLfz9szfT6cDiqcm9U4IzuTZZh51jClHln9v6NUWmuJlMhJ96nrw2O4/7zIHIA4ahBSRc9DMIO
azRtelcjOXlcYZb3KXMEqANRb/8xSMzKY/wRT2jguJ5BIsMwuT8vyKtoIqZLpPKcef63lQjk5JvG
DKj6J+1uYLU+2m8mh2S/NO+iepJhYBkR7Qf25XJOmt3lECBXGgMG4TD9SY7vzoPaKOJ3GgZP4zW8
RO0DirRy6hcBkM/2ANYOtsn8R7/TjNSpkpu3C2+ha7zJijhatIZt5Lrc5CCF0ogNok/05p0J9IA7
+IFeZi9rFefyDy1y0jHTQl56VpPn4LOKC9Zbc4DNi1u14cTM5IzZSEs/OXLmA5IOr/sOs0UCu9uI
Kb5midcLPOGQt+RRHVbKjdmazfKY/1YvXHRioX58hzk0dIRnF+YSef3wRJgvGzNoI3cJDcDdMmlg
HHCHg5S71/AHRf1AFP/SG0GqJZqe3UeI8eEh6d4DtZbryAGHWBcEawY2PBQJ18q97pG2Aqd255/y
6Y/L76NZmp5qFi/m//Q76d3qxXMQyX4IZkqHXqcmOwRVMY8mD71THk1UFV+vGZ9MulDZ3ZHtrES8
zyQFX3mlbwtcs62PH428LkmSUZylHXndEkhAaldfVAkpZ/5M7Cuv/Yl/6EVo89/QK3j3jIMVUDM7
nWHkaaSRnI/+aU2kWGeRQTWueJpI9twuQe84DeWIZX8CVHTVEzeFd0tWOfzctAMPHpT9SGt8W1xb
4B7GUGab0rIXZt3CUjmTXy93/xyDa5ZGW1nKfkUg1DbRhUGDsMtjzbmO5L4ytLUw+oQQeBi8DxLe
WavrCOW1FjLcQYkmCbjf6zTAlMHRSZiymXIziqd+Du/nECshZs+CPrAzlEdLJ6/1A0tUhrsj5699
MUj/CO1VVU3i/Lj5EWFuqxyS8HHzElapTpZcRR5osUBydLv7JnVx+Ca9yl5TGYbt6q+PTXKqNsGu
m1BKbQm2CaCAiw59Lr1TbyZm1RU//iNtFdBSikw8UHbi+tE/Gx9KC0KuNKvJb71dOSO5qFa+q02T
hkL7efvP3plB0LN1Ma0epd1Uah13XC1g0g9nZwMep7ILIfAqTBG04hYwLwfxzVuVEgP4vTsH5YDk
3Th1JZ12XPRP7sx0AgVY3e5YtT2JP6ZiBv3XzsQn/lM+52txvM+tqXTgwvAPgMkm/Y7IfNvLgJpB
7LaMtYEdpj8If9hA1yzzrECnjR8FIW6J9WDCBnxQIRsapEJMMKnc1kQnPi4SXOCGYMu8WEapk2wW
Wn4VkXp4RMjjem23vjIpw0nd+X5dPBwwj6sQbAeTN2/6aZASqd6nfNXA5DQHorbBgM+HLDlRRZ9I
1QQ9Bg4LAdXfaQGJTaQ2o3mvT0KVU2grAgu2lm41Mlej/llPGeU6Oaed1F/9/5SyX3DsehjJRXzi
bcBxLxLD4oA/XqG30nIpU/kBjTqWB5tardt7rp3U+hWJiLFutDkQXeHP/p8GDFwFmxmI6eMUvsny
1n9LAfQz1NiJj9nY5aQhbrOnxsDGQ6jIgFCghr2UioBA5m0CZ/0jhAAD/876BjVo37YJyON1N4YL
2ZlY0fg3GOhq0hPzL82ybJCHx2n8naA/TT3dztB4N2sf+51YK6FuyBE59GXq0N1GNQv23GNkUlKd
7h0woFQv2dc4h1EnmXP6Ml/KKK+PVDhgZG6OlXAxxU1fi4tGKTaUzdtaiQCdJ1yHp+AocTC+UTqg
9s4jN8ID0ohhTc+lrd2qk6j6lUWUnNGmNKXZDg6EsCqzt/3mjM7ZiBVq32jQzYsY7zj8HW+LqrmK
s+FVoq2zYMz8vxtpBRhrNlgnwcRciMeEhbgyY3OedJGbeTr/HFVcLLcCLrDb0zGb0wAlzHX8o3Dm
g9f/YmzX1c6Ge6MA43CI+fu38XtscDasot4nk5n1wwSFq4X0brwmz/302DIiRZiRgFvoTrDuymIm
NU8rC4JbW7E2BmSA2Zkd96efU67FLOtV1YVMynReWPnpmrORvX0FM0NAylS+42Uo2x0hGItJwbiL
HymUdHO+ka4tnug9xuORkHn0TShmKe85WKxCuzjH4pqYREgXWcr1YlccnjP81Gz29SQrmyXaAXTg
zdMAzzlPRNNEQKlS1BWRtpxlkaGwsqk2mMr1Ev/INllsb1iIoOUA9S7+XO5szsLxEBF0P+AKU3Vt
6uvPRLfHD86VC2G33VdeH0SIhGZJ+aqTUVbDUbX0CtKJGYR0S21tGAT9chwE1lRl9fUW+eRJpLlM
39qtSAD/aZ4lOCkA0VzaCjZVjPJvEi+vVmGsvUS6eDFDR3jjFAablkoxyuwAwhNbm+4HT65A+4W5
Oi6sLmcYR5pchcJgKlaX/vSuknYKemVCJzGio2JnbGewKSOkqkN4MofWUSnMIyORKb5NJENKzZ56
LwJBSGzQ2EEeq1vrShH12c9eOjltpkRJ82VEWOAc5ASOHn+anCrDySIdF5tlZ/2+U9w1jNizOaNd
EDpl5ILb2fB2vu0dLYrxR6nLBrFcKeHADh1xoYm2qW9N5S7NFzbUM/omxI0ek7nx1exbCQPGUaJX
DEWfhMvYie2UFty5gT4l/bEeokiE3Inclzhua5nyKfuKpSRY+8O5VKf8rHfZ6dJwEwJ2bj8c+JE+
tNaYgvEZB4RKk32H1pVU27Q78JQNqfENZJhwlFLLfov0ST61UsFW19LUPX/+495ZNbq3rSNj6wVb
8Qgcfsq/7WxY+Dp5hb1revFdfbEKUBD9YXL3gN8svvgAHXYHMxoCwWYOC1Ff3wIR4+0DChxvPuql
uRhSF7tWzj6JGWcu0G4xf17Ie/cZhIa7n6OsQai+a1liF6QCJBohLWMIjaUeNo02jfsVrlgxbCDF
zz03OWEyqbpHAKuCroHxpumxOjq563cP/sBgjS4+Dn3nzxkejZ7XTbw2yQ/mJgktqNGvg+3cBPxO
tlo8U/CKnHH66O3zaeRrQgABntt99hbUjBL9cQa4BbIX21uOXH9Z3B04lN3MTlSAdQHWv/3FwBFX
kgytFEAXH5cK81Cmuf8DM/AsanMEURoqgkcpH5977se5tg+WZ63t7SAxV6eMR5krmPTb2yN4TwKF
MLp2c4a56ctGP6t6g2SQavxuDnpCjTvPgIcvQWqMxam/8HZ2bQncG59DcqITdr6M/zbho0iFOqL8
s1IZuSEj5oO0pj1NK70nilj+qFhrnfL7sUFI3UUmEQOsGx9Cb2MKbUGayl0RepuJLXSXwuqGlJ21
KmZxmrJuodRFwFhsLtgBjsaws5B/7nTxMLDkSszaR8rCBq6Z65jN7jrXxhSrWYUokdjGlXkS17mT
3xaMngSB/VSDy0oPHHhEF86xvKYSFt1XJY/NBpOAC+j/88doPMQyqqCHxZSxEyti9vn9EsuqsobL
pSXkDvu6SJs2O3vaJ355LUYyEL/u7UcbuqmjXRUohppgkXkeAuligThTFANpuKOcTcGVRQ8VxcH/
0BIfjNizQ9Bn4rcJ1FjMfYRGwyVGfMP22gMz8trj42krWcBaUwnr29jm/u6f5TZSvjQGe9XV6dtc
MSEoejI+1f3NCVdYBGeWJt1yc6Tsp60qPPJSqkKSEBM3krI/vm93jYmn/CiuqJeAtEOwJ5JXh8h+
+wHh8nztgtXIGD0zEk3PqJaGkxyn2uJP/2hFALY/+4Px6Ib4HdLQKitqc2ISCu5D4tZPvJv4RiKE
RQG2uxWMXjnYybZbwWZBnP7UuSBnCzUco0y3sNSS49pIKNndvznbo7pEzLHkfmvKPYjBcor+N97g
WiXriosh8PnBDh9s6NTSNc97gbBk23mCV7ExpGi2uQc2tg2SaboSIlpcdoIo+V/OwY675oxjbcge
uVuLsOG5XCVISL4yHBDrp+NH/7e0UbxhJwkenFB1lDt7jhzwDAMQb0y2d9Lt8GUjWVPqpTV8o35K
cGaxlJmt2vg4MJkjkLFwGHnwy/NZaC1nG23FBDkS5XKAszVdCHMoP07B478B3Uu/us+P8+3hU3Lp
2HOTsxkgR+GolxF+TbCMAXJ++vx3p0nlLO14uiEUA4qdInEw3ZI+RXbDe4aV9owvB/sfE1yGfhBd
filP0assuCKNtNy+XURk6KsxX8Nct2v8E7b2vlnHpfp/ybdiK94zX9KYGbHaM5H0Wv007PPiHs4q
bR3Pd7Y8AwHKKp1TjK2EAU38M8g9tho2PNUlD77SLQ2kzl7NwVDySbUW/04WgM70S71gVjexWIsn
3ycSsNsrYxslsU4o9cV5bXDMTfRMSvBJqE019N0rIJIvmUzEzvaPHgoknTwRuT1w0EGZ32G8JLGw
Q9IbLQ/fyWsu9s9wdSiAL2oRPb1t1RMHudJsKd17+SI75aFTE4elpvHMNAunEE88SNWvyVo311AU
BtOSd2YWGzuprLCTwsqxF1jXN1XhfttrmOnIJP+KOS4R4z6ElC/DCeHttbS2JwgIjZ35+lu4NE50
aonHit3rDA+AwHP3q3Q24x/XIOcztP0o0tUjBCb7uRjd+w8Fyy1Rvnn0ukeL5LJF9E7ijylwBYh2
csCLBvUnwPbTKqrn1K5ZQY5x++LPqy59IoMShS+5xRkvDNskH2lvk39adfue2CjT62gqp7E07kUm
wZD9e/TtextSRGHzyyVFYwbgVhOh+39aGlAlbxis20sACunv5XKcTe584PT9NXaSeDCCM+uMNjDT
TftSCmjJ8cYja7iaojlPWuVo4EkmyrfImI8iHwnf54EymkfjahhmSdbc8zN06BD6WAgFs5kym5Bq
LSMSajC9W3fQrQV7N6k/mY9fE9FZIW4zsDnhdu3Y9h90FjJxlnvHupeok1HgFHfq5d2WjyhLucoa
+BYh/4aw2o819Q/vKBj2RWZK/P4zQls4b+kO70WiSkAJKFkZokGMEGELePwIHIftVmvasljF3war
PqmDnbDz0T5B3VB5NV1B/3AIx6V4RysIPA6UFaHjiTll4ovSUBaHjC8VhENA/NOOh+kKvqnD4bdZ
c695f0OBgGDAzX6j5FMz2MR5L8Mimq1yxoJDkbDVX3BZe76eq7Nkp+PLnIkv50lr6RHEjhfv0Lkd
Kzblspqhp3sceBlLnWss4fk0GQXg7BJUS8FBpcqokarsiyEQlO06rxkuXlBO2W0EjH4TXjnTgiuB
/i8elQuIqkglFsAQcnlSTcI/yXlYpY+irG2ENvxC/ZfSn70wR/Rr4jw+dH9tDe1pE1qEurm6BTcM
46kLzIezZQANkaFgsdhmsjRTrTUa/4RRETbev4sNf0/dtPWA96PiEUfA+S7iYR4Y2h6wHmLWa/CS
WtaL7yA29gf85eElI8NXlkOMpypbqB2RoxN7ZeXvQ4wlS8N8ZVxCD82SMMQtf9H0qDUr86Ceqao1
EiNNJCvpZ+PFNgoVKtzC9WTWrsQiAQD7tyYjck3oThDIPM3/rdWSTkVVEOWufXvUpAXCcFgg7id2
jgU7RMNETjFjndC4pgWmYBqekGVsm3rfHXabbP4ddVMKV1NF2L75so87DJm+OIVrt/psXmDYIJ3n
YJ0CkawcjIdbLpcN5MQBE+9IjIROvWseCzqN2baN89sDh37HtL4pnI72p9HPm1nad9+RrfAkdNzx
K5RMs9mTnsIjIj2p+Sp350KUntqOw/1Qo86OEsUrf3uZf/FVBXqqPFUpBQ4sxeZxDypp/Jyv/HRd
pk38qX8uIbBUivSzq0yX+9ArJL+9sCFtlWHvn81EJZKr9U5NDq0L/+oRB2mIbxcLKRDag4PyR3+D
n9AGWAFqZ4ht+wmER6hOm8c+V9z/guNLtE3cl6upyqLxJDZU88M0vZEJYxt9BrkaJXymtArJRWgS
IVDDe7m/PpE9MXirx2o9Aoy+rG3mhR1rb8pDQ53LhFRecAl08GYNsJCGdXrKYji184bkV9I0zZzL
BUaCoV+27KN/cik4zQUWlZd2OKq45e40QiANy34ysJontolGVCnIs2D3If5JIAx2cH/ut8IaBWCl
gHW1EiNaspHbAtp7O6Oeoo1d2QAMrMCkWmX2F5Sc1uZI+89gsgYonJgNw2xat0awZRZ0IzSvunOl
NjBYXhPrJsezyFr9VvJ79qXmWkl8EK7OwWh5cu0IaCxslOth/wd3FHrJhu7E0otlB/VZ8Qg8eWf8
1ODUDZrGGgEYJvfIoBBbgnMfzdUrgmFIg2x0uKfUZdNug3XG2iTvM4ti9TqGMCBB4rsyeEHmC/iA
gS1NSyGxQweDrXkGQx74HeP+xcqrZ69GHTdPJseKthGinVWZTEok5XUzIUP4n1LFhBDd7TIOwUsx
XVBGML1JWq87YzXSYIJvcmO73/4DtN/OxNLRoAJpNQhwMMEC7ElvrLC2NqIzDot1quzBzkf08XCZ
HEL0RzFFZSQJBvdKKWsgJ8usjgif1bko+9pW/CTPTflFruTAOShJ6x7m1JJIsgc/Z6Kva/KQC4zZ
qHZNzji7tEpVB4K/1XR+Fz4ki6b12qcoxkRUEG3cgCV0y7fNtVZV+rEOrqSG7rcuXKbol1dM/WIr
Zu54CkQj+7dpjDLBhxNz4YxahD99HZBHO6wY5eyIr6UZ7txv5uor67dvMP/0rFc4Pc8dkgAPDyX+
ayIdi+Qxq3XiVwwYltts7wec9lN1tDJgHpt7DQOtr6Q7Nwf/uOWRps4q/WMjZm/sCcGmNc3R0rCk
LvvJ1cyExWIKVG8KbS39XYJ8+UEBZrwipfraC742ZZJFNLQyEilXXJ0cv3EOFNiCiDb2AFHriI/b
LbY8qjjMNGHmJYSmcovYc8RC7IFTV5CAML4v0aDSzZeHZJZElBEc0UApdUTgamGRRLZD+Xhmt/j1
YXuysXmDsx3q5AoEcZ0L06tVjJox+VDNoQuNv/KopuPV0aw6+hkfQmfPAgHd7TiFf9sP3BUr10P4
wdQujy30UYwO/Rgz8SNDdwV+wyZF8xUSDTHuD9GJbZqryfP38MTNVVlp/mbX4KxuawwCjMwcP2qs
rbxQka/dT757aU5ohA2Z5+ALIrmyup2kkYLfooGjb6NPZw+TpduvNzZlSEBepJhqKYZ3RSuKrpHY
Fz90iD+3AYc4YyLqQU/Wu6WwatPUshgTd74foQnyD6uas8cb52NWtpN3pL33hmXvoZWboswJAjVa
rQ07/bGrIBnYcUw5/2nC5L6tA5dDJU0oTE0lqRLyfLyuEZUKLaBfDHwpg/xL3IX8ERMXjDPVbhH6
wJnxEnMbHCdYF3/KxMDs2cClo+bdHOWPB2AR4Nxxi2A9udRzAunMaroVkdI5PKh7YHP8SjGZDHiA
fEebZfKIgtvGvge9yn74LquSsTuFi2FQDxBjIJ3/Yob9en8WmtLFhqbDo1q4C7CxsK6DI/UnS3xt
KQvQpPKf5AGnmlNCHoZlCUeH/fByvnKqZ3H/z+ZK9KU1uO6h5furwgijAbiOl966n3RFbsoPG42Q
v1Im1BV0/T14GNNZwzmrKTMGi81+sgyKfFNw6av+Lv5qrB687e2I/5awQsnSJT9R8U32sNXK/qZD
PhHErRTjuJHP4zTwL5mcDHRuCZkrbNaCtYo0oYew6ERERtuvGXAgDJ+MemFGzUjAPjjKCuK76Z7C
8RkQnDWfEE0BI3KpMAy5NbbB0ESaTgTf70YZkmPleHzAF/4pomD8eSsUTQp8oYTQnffTteJkZc+s
jJ7B+iMRwz/wgBpKZPollqnxr3hsrJbStkULQF+bx9mHjlnJ8V4PPbZTjTyCSjKgpSWOEZu0JuWr
Fmk+N7iim9e9wcLFyJtCmYAdTCWVJg2Im0XXXPRkAzmVH2RnrCp8x8sZw153w5Guz6kEjRvZJKjj
9+LlxZaS2O10V9yDQmzHUCkbuRGghiAFrCNdi59rbB+Vhe2UJh88jnMM4jK53gQAH5gEMgysPc7U
/sXvgBz0c4dwcx02LOrgdovWCrEtENt1zmy5hP3q/rLkCid7ATGTgFKLW+q8O01p9ZoD0Mb6Zzoy
fYPIKanWzowfCzeVSGDm6hdQSXzbg/F6vRQUxW+HadLKzGphk6eRoiDSFxx5a/6DMPW2rE4YPtS9
ugNhdxcZT5RdmQAjt4vmTGmoAMx8N5IsaTB76iwjrKdGjwOzLovSKKwMBQy/Tc+JebWtBfFmp3rE
uin2DdA79SmLR4TtJ/wBJ3eZvfAjmOMP+G1xQCFm9VHQWZsaLPVH20LbNW84XcOOnnpTqZ33KWM8
p0oxbvSlmYgHE2EnVSQF+b6e3WvEkAi5LfPLynpF51rPW4TrLRvxD1PA0KVrZPT0FU+qDzOHiZnW
nY20hpj81llxDnr1askV1cOyFX+U046euFJwtGyXoclRLea3mMcESfgW4xTqygTxrvtuLuKFkVUq
vFj/gjZd3SvO5PPGpYBLs1nnzrEM5OIbLqlcYjljPCCJ7kVcRWLVA/aWsosYKzK+t7uQfRedfQRq
NCNovOkel4xATqllp3gg0cxSzW1i6u5f026EcArRhHGrH/uCFTtC+POGSNjGJRbRKJbKnpDx+qwA
W3icWaQmXUJOUs0CRExx266c+AciPgig9g4VPoHTrnlkWVghyId9qFcVeNJoRQzZcYLjQ9JjfmBr
ii5Zrd4l72WKuiyYABkVMLKLRQJHeLfGc9Pmt+kM/iwLyI2u1dK10NxCpQnC/+5UNEwU1vwgoK2R
QAnlGoRRJsxXQEUyuytcs8RXNErjbQmMT7RhiVCKPKtpX+V0Yc2slVcvUj4F0/20jJKv/0ibSNe5
zhF1CJY2g6yK1kE2IfqAt0IovpagXg2M9ZjA3JOb1RnkDyvbexI+8jkRuSx+fPBtKNj/B84ORTjM
dtx4wW64YwpxO4C3YD3QFSFpyALNaHdRXO5JBLEAN2S//CL41PthsipbkzsyYwInR8oUD18y9qX2
yuSJBcEc1CXwruVrZ0cVMdSBtGgJg6P4I9O7mhBuN5d61n2C/Myk1naso8m2m2prsOYdE+0uWVDS
h2kzXaB5ngXmfnNeIObIJ5i0+Cf9d9gBsTYHJulnm1oH6+IiCyuLJ2liz1U4nxbLduPK2rPBWfr6
v1WOpnvS2XndayGYZ/CS7qrVGIUIcytJ7v5DPn1m2v+wB5LU+LZksjm72cwf181UYDFb3YLkrF+s
EKArwNpaeBsylaAvb2agHtludq3dz4CCewJ+eD+M2SL4F7J9xZi9m7CdqX0ANz6Cu2kmDNNVn8WX
oAgZQQVbYX3injK/30fhAfobRBo+arEJXzUZFUscL+7HXrZ3nh8KxWV9BoVBgFXJSB5wi5AfeRTy
MyEUmykKm42UJMLIiLZvQC33ug8Jyq9C25mogTVLYVqWYI5N7sNdv32HGLMF7NG8Nx3YB6aoWC6d
QJQWJXnLDK02l6Gxp8qw/04YWTDZ1z0CDowVfIMQG2wBnRvwg9FVxhx2O3w5bpVLhCzmClLUy1EU
VO6t6S8DBveRsO35ARQB2uCpOgZuBlZRgzNJBI6YtwBbyatvhCTyCKxAzoJkH2iJsYFdiL2VL5xg
4el5YBEye/C4CG/v6/HBEU3/QARBl2Vl+uu61wt/jxNlVdXu2X1vP/0mRPTGGTI3G7diWleDcy7W
G3et/iLXGYkyKcxVze7UDWMPCJ4MFScDt8G4wY23CfX0CReL8DXKmbAvpoFULkeE2PFFOmoXb8T5
RvlkyBJ/ue3Xg3mu+Od282DdD/La8wrluS13ZDQWCdFjHPbCKeBhdVAoqV/fS2LJATtlLSxXnTVI
FXLt+4UBhcwkSoX1TWOXFMKUcizKMhr4A2nBNeePtxqzkCy6gV8b0sRBLnBlKrO7T+UrlCPJ8dhd
0wYY8ReafCUo4uNbToFIH+E/xGI7Bt04QKYnLL+imFgT9Yapm9hmtHp3WZ/ynECRlewXq1romEJf
SZ95ANGn3GaTv0JyBEo/WKGs29ha1oHGncyrfDB/FMzLJivIjUQsS8u5zgXhgAIP0ZNgHZmVI4bg
AQOjOCSdNisxGDc+kvm5FD872+juYaCq6NhpMjbdhsSNsZ6ExQi7Af3XVT7KUBGhZtW8eWmCDAoc
5pC7OE/1LG84dhQe2ty25RWyBrSY/J1xzF1lEQtb7MxVtlzsVgKUXFkscHBntO+GH4Su+M1JJMLa
H3x5h5JtSSAiQi88JXxNbP1UyVTShuTOVV8G4Rw9i7aL01b+0u7rsQHevrjx3gUsXoPH5X5YvWds
ZpQyzXfqlCTpgraKa6jIZQ2H18lhL5A8OngNx7kYq63l8omfBoIcln77Wb2hgGXBRz3PD+SGUzbM
JozMo8bTqY+FI8Z/o2GBjbdXniXN8pV9/0tm/BnL9Edzs7pZ/oqtnhDZmn4F4Cgjmck9s+PMC08o
Hs5MQKXrt5oo0+HRxbBss+dNwEcWaBQtL2UfjQPICven6Xgg/g4MWEbNIe26/+I7vcys0gpHzYcV
hz5ipoacx147mN18eefr9ELtFWx64LOmbL7/bgQ7+SfGo24vZNsudizeTOoGGYhU1Nwp4ww3ZW3A
gOZNiUm002DaNv1F2GA0Blerhv1JP4fbSTW6E4FsZR4xKz7AbsVIAtol7jsaouKDez/ebiliypRF
idB2k95HN6wuv9LqYIjcaGBPIuTuY0OQ/oN3vnpF85EH30y7yaJh2u0DJpDoIvJGp6MVgXLjC0Lp
fPrjjljvd6/VyB403C92f7cCppDwf9mI7VAFcROYnnHIivjAahp7gLV1gcW+TyvRLTPWoVJDfOIH
5epETWJ2Y8e27LmP1gG2VB0gfEy9EX/Ca+GR7Y2DJxJHabs3pjefgOenMec0WTT45StGqJ235ofA
hBc45JOCdy7dZUMBEWzc2J7boVdglXjdyrhorMBo/eMoPHkjmlXBQoeGDqFaHBZ13GbqWBcYtSvl
vlUMSfYd0Xy3rUlXtK/TtsJUSJp4EGfMTY5AlGxqIuitfOp4nPXjK4QqOjJepDgYBpgnZCSdulWM
ifH5nYcneZUFkszteSJd0AKMg2r0up2EFUW61N4frOXEpG15qE5WKblpt97d1hECueulX3sTSPIk
DQ/F4nmzSkSGXeiPDmoHCo+iW3CEBAOPKHhaulPFy+eSLU5BK9QOv2HEhJ92pozC875b4Ui5uWqW
FXfFwN9y5A80EwpEDyJmOiVtOmdxOBH3Ye81sLqsNpqWz0/LhfUXrVKqaZoNZGpm5nOWo8jyMTR1
jML2dqwb+7IKWMAJ0vBSDE7ONnmEtlAnSBiBV+xH9SZBF+VDjLTD8D7wWPs9mrgvNK1g0Pau/LRR
IT1f6+rdONfjBwyQiOi/KM1QIOYi0/8TMoc3/hPPBY3nx2AC5aPdJLnSL0USmc6pyDM0Ugq4EyOw
decJmnm6x9MMMXDAayirr3mrA1vp9T6EhOTr8052F7kefV2M/Zc8VOtNnI6KdIxu23Z3lRtWzjgO
7Aog1csEGjohFyKD6Klr9CjHIMnoOO1hkCI/8hdLgObNDYoEA4lqiYbYM2i39DxV6xOK/QSt0sGy
lFEN0D+jMMKqIzKEqY/3udANuXG5F7zZGHcAQh+Ys6ya0AcaLsGzL0OQJ48Ey+Lk3ZJkQP6SMBv+
tvHoFeqZYWIodS7oYOptNaVINgwM2IzUyYvyBo9JLBN54qYmGfSCjrPw438WQ7hSIlVstglY3YOB
G6kVWmTNDcGYRWiEabEQMyZgzLD1Iyj6ZeeI6pU3vsU3cp96oXimafhmjXZzTQ1fr+Z25tEZwCKY
OAW8K7lf0G9N2yurTQws/wqmB0SZt/nWxEGdq9a0uszq1MgI2hbowfxINxeFKjxJg5CBHdv95bbI
MFgeCUzHiy8zrMYMB90FKOFh83uPpbRPbVDNjFiMv9VF+484EJtBbpHtn8U/aphy03Zg/fg63mZ4
SGvMd/om3yIDaIsu69q4e0nmRLbBFOZUefEEe8ew82g61H5lGfSU3Odd4hFIZqkOdRIc/0wKrWkW
cNGbJYFfDFIC4Gf3Q/oVZEj7KNqAtou/dhCWHsnViXYHiiKtYlMSQGEba39Gjw5SW48EpWBlF01I
9urwEQDikogKeQKEW8F1PeEdvYssxpVQV3WjBavcViGXKHZe0m4lJ9MSGHZj7ZSIlL3Z9yT0OoTC
OPnnADl2zle++eIaJ/k4G5qdZUJ+yvIT6B9Iivn4xYxOW9Bc7N5dlyHqWABNIo3/bZXojxPfXZ6R
94S9+QotUGu/PZkG/gM6VbiasPsSU6PTtxgLRJA6DjKcS+241N0+8+Mk+NoAcadYWZsYwU7Qs6xC
dmCLfs1oHpeDLJ2iTsA7WOdbtGwk2jgpM3JcfhyJc3+bNqQUy3QBFCNxAUNrPL0xw24xmpyADU99
D1AdSIIGD3QFIHS5Zq06wIuuS4U+llm/5nwD13QSNZDIoIFLzMyKkNzh77gtaalebsID1FofD3AW
0Re8HbBHzuX47wlIa3TfNXUL8ZcikwQoHlE5rkrFrwrf/qwA3n5MP68p/oBkdaNdyzk2pyCgRApP
s5z3fZtPtojxN0pS1ms7x4cCWRXFDU99mqkm7iJGJttrsjSTK1xS67BcCAHhgK4R1ZdThCKsYVbA
Y2QiknFqreF/ee5nAWJTXZ7La80cdKMHMPNDCbgKfe8obBDLVBT5W3lLV1JJAUsJO1Fd4FrGqK7D
Moz4AzaFKq9T7e47nXrMODrToox8IhCTgZSWsonVP2Hs1E75C0fCX0Bo5rf3RLIFlo26+4ashQjt
8k60m13cD8PcqfJ13vSo+q4OvX29usSFxn+3HJ4mWnG3Mf/3pyN0pAHS+Q5Biyx4cYxpRCYu9lhm
/ge15w5OcDrFj9yo0GifBvalatPpA03leQRnT48EHkUspE8KRMlIJqNQC3m4NTU3jCdd5sBcKE1H
vMbTykOaiAWCc0zub+XniT7BrLtz76cHNQC/qz4+ecbAOY9JeZWKQxd7zjMHh/vpSYB/BctOkKV7
JkXhdCb/Nrsyq3Ae/cwA2c5YERE1LsZFFs3YTpEUkOIa+1BvJjvWJ2h8WBE7oh/WaHhexZE2w8vD
/u237rVBOjnU5e1xsV/vO+iC7PLIUNDmtsqZ+fezLu3W9dgAznorz6CC4MlU4XmRmaAP+uKmFgns
9+oOPBuKq1xdROxdGgYfAI7y63HnrHM24b+WzZqB5K7ZuZInSNj/RqLjjcMO65zrI85C+RM4JRH4
rliJJ1PoqbPb7l0mvJkTM8B6crUfvUShrnbkTWhTNYJIJUAXZKLkCIRCNIIMUEpacaywxM9uEe1i
KaiqN1tI9Yzf2ZfHPhNmxuaBtmrRnE7YoHgzVlu20sw/ff9LBqPz8kBgzTMJaNajtOvdMZZtCinh
3GzGHjFfR8kxqTK92aLGLHox5wNAT8epq052flpOm+o3+HU6GnoNN96C0MjcvPa62ImoawwgFhvj
PW7zOEaLqMUwcMnpPZHZoqxlcjIICP1UiJePIGLbrkwDOD8uqQBbdnkZ+JLGrZRPKHzUuzyYEgne
UQ1CpoOKt6UfJT9z2k3QF05zePm3FZN4fw9iZXjUMHk+X/rRoMToM3jazDKqu2RIrwCuiQsK6MgJ
U0dxuIf2RiB5D2CdvmtDpY5cs46rXIdOJO5qyreNhtLd3eXj55NayVxayl+Juh1uXbMBPVC1faUv
egVFQBOols68xhHVOSD3UY6ZxiBRCJ9mvSRXTOZ8fWBHx6uYN/NKx+/HC5/AqnvlHZU2swGJhDeI
MWJ0+DNlbjoNuckLDgs78L4RSqr1jNONxMEMr+ExKQpZo9VgE9tdN9QZx4tYgE3Cl9Q+NWhQrrcu
jkiFits28l8gO9x6NKrbd28e4TxXbPTx2pGb7Tip43yCzPDDsktaMRJMsnkAOnXr/9XunmDpcFs1
wiI4Bzg2gd0PCduUFXS9mbA9KTUdCwxIQEVl9AtB2y6ZxhxJ1egP19B6xN8Vwd6kL8iyq8L5JcGf
ApqUkqx+WkAYATpYFN9lK1leQKtEnVvzfJ7gW4dcZCaOtKK7Lb6TQ2sGetCAtIF19ow7H4G7mcE8
+XnYKwCyhgL9kBuknfk266Ds/WIhPtyMnbI5xGUpSKJQSrhd3Pth3FbcKFKvnwto4KmxXd1WG3Dx
fJ1sQi+5pFo1NrHvo6ZMqpEHSNEIKzGNIQShkowOidDBNKVJD7OXuBbfIhWerrH9W/OIJXD+L6X6
qrR9tYx837f1+VQnKvqw8xYVwDJuxM3l7iAtSvazui/W28dn53gBWI7fmD2iVBm1lxD/trs63xhG
3JeqaJYNW5ocKFVVOxuFACU5LKatJI5aKdYVJFIY2HPT2lZOZrmHY/gIdVMEqFMUrthhqxu+BZfN
8fwsVURkhirubbMT6v6g2/2ja49Hb8uY518mPXrhDAGzefg/ZOiwpNoQN/aVr67uKdAdNzjuvMTr
UZ2VuM1fjzFpBHnoktxJTWWbQtY44Emb80a6E0kov9QXnXAkNca0GvlKKcd5Cnmhs+Ru8Q63FjVM
6g/zxEC6YeJqDvHyHORLnn0v6ZrRlquZ7IZg5vq0kVUOqU+9F7ECUfhQNqWx5tltD/zuz8wfwmOV
U+1hrklKNCh6SJE1EQj24mXq2kODPbgP7dv0ewFxiEpTF3XyIegIRyqcfv8x448ekfVWXLFfiUDR
S64pySjxKcydDZUoRbhtfXsO+hHiu4Mqc2+gSfHh50c3n9UlMw6b712xWM2yeJe5lbhjsvbCP6as
IGWeOWfDlFolsTnoo16l0dRb8A7t+Plrktf8eBn82o46Ss4ozFOvNX/XXckKjzY5sLcT/TSWtI4O
Q5fMj3A96cwV92BsMVol+L9Vu6ByJjkSTmR4c15TUP/RqHEghLQwiTV0MsjOhkO/HL5hw/f9WCfV
0RuTeS+iMz1Dt4ozJKwa53tC4lm2DRNen9CVJWqeSmNmtKvzEe1cunv/a+4B768mnhAHxQkIvep8
tO1kcIAdi/a/5JT43gFBLYA6YK7N5x7LSXOhziBmGPEP470TdvPMshGtIZk1l+Cf86aNNmsouTDm
fy4Bzq4KmfslIFpbm7voKy57JXBXxkiBhWE9MJ4XoPkOC3jXxuAG5RibJJAysEZtHx7iL/wcRsNo
v8gNouLQxUbQbW2l29sFzkN92keUShK0enjv8A7IsWmKM7SUkYUDw+gQgOy4jsD72NxXfceUSQmI
z3//V4kPG26PsvaxO+7cCDY+lqYYensusPJQj7MkegPk3G8+BzaxFsJqCFcHPszNUqUOSLVjcgK0
qgxUYp0HiCChdIbl6L3qsN7SXQ0sx5KYF/1RV8XLIdXOjwQvt5yYRQa8HwQ8PYcxREZsQ8KPTHKG
3DImWmRcjPcf/UMxjas4wV5ienxkHzNTycgRMEfitS7cZajdzjD9lOLYLVdJ0+/IJjPfN7bpBvcf
fxSFaI/hNB5DWVcelxH07Jc12u2dMLG60vJaKgWMM6MJIgQeusOg1vmAY7kBWba7vGq5h1m9n0LP
AIY1PKDDXJJmQ0aNNDyyII5NHCQvK3jK/JD7WZBDwIYqOdF0TL/tOPsvywK/dml56PLoyPguvfU3
/vqz5Kdf/uS3JJ3uJPXI9a7/99aFKmZ0XG6vL0g9mdPox0YQmM64908s+u+8UI1yPwYkYOEd7Guu
m6OskjKOYcEs83LI0wVdrXiLWeJq6XCxOTJqiGEjPEE8CLCsua4QLkTZN9rmbwF76XTzwe8aotPJ
JqdbMbCNOCa58U61tgZSc5qcPvjcxPV0d1qmKScCV6o9+A5zLfzz5Npg/o0i9VFPW/FwjorjJqR+
SJe454PqTpy0F3xeW14TYKi9GNXmx7Bb4UQm5eq4cN+E5HmheG5LXBAcFA6SPB+VWQ6XfIwoN66V
679L5SmLcjDPcas3gcQ3SF2IZl5qO67LXyto110k7EVdzHGNjMekRR4nihBdH5yg8JpAm9j9ISEi
scTLGJnCZtT2DUInyOf1wEvZwgOvND/1aWS2IJPEuNVhagDAmy14iAXL/5Wg9wbK0K5kcxnHijcy
63nw3uPky1AlBccANMDnIMNUhyfzf5MLH1wLj6X8QydihJK1d5fG4N7oV9NNbp3Dudqjtuf3E/Xu
1nyV0moXpN4x3CXGUn4lrj6IypdKTgdqpzL9zt0rgVpCQgciIQV02pQJxCs/YSiZKwLS9sHSsYxt
l/HYcn59y9WTLx+3TGnmSJ8k9gRG5FiTiyzcb/iTMy96ctE5YIEGjP3lJEFO2c6qGxSyAWR/2En0
Xe/rAfoaribFfghzYy4tD2UarBvtbDTJDLRHdjAV+ZuBe7C4KvI+OGKt4lkmXrmXj5QWd4P5D3bf
Eo9mABAniuaT8G4mAecy1cWIJR5Bj62NR77KpE1PWmaOw+wBF2M17J0e2fXOKsIdB7hu6gELmd4/
v3sJNcwzyqcWMSpNe/IFi6hGVqL7fmYMCZtPfkQxHtfyVJMV6otNXL7tk7Jpg8wZbG3FLEoYTEwr
LPj0mTIDeobL4jA1P6OIfWpGCBajaYdYI7HtCjrzKmjikXjaFYGEN5ygReOreAkAs85TZHUOHjF3
874UGeAaUCf2Jzq3vsAi7PJ+2h2G/NZUrpLgUCFNAhZseG5ODG/Yi/j632Oh7O3q88in1XfX8VOF
lKR2CWMHFX7Ucat2Nfa4DhoCTCsb2lgQpUT8/DWw51J4mGpFDrHb1Z5CDhlZK0F4O3Yam8rLdPpr
ZLQCOxjPCjHUvc5izAWgKRo1N7U59DB48gmbdP8QqZgS5dc6w1aW/hvse/gY8GgK0lnLVirenauQ
u4n4VOq2bFPaJ1Qpic0Ho5vm5SxldidN0wp14ZDck1jzpW6CgnzS2FZ/2UAFkVdoCaxOTvPo2bF6
SaAzp4bBIjJTHj6VJATYtnJ6kWMpvalF9H7L4eI+rG5UxfUac3YGQY6SIAaOezZT4jItcya/Lxha
M3L2+abewgNwi7HVmvXcdLfWWzemTaq3TwT++O0N/eJ9qdo07M9Uw77ebhV0d/W9N/LmabUWlR5G
hSQ/YKUvYGQ21Fv8zWjaZdXbXtu8B04oW4yCwoLApF7CEshT01Y+joeI/DPIdbatVFYnOCatpJ3R
kPD2VwdYtP4yWoVbsuz2NSPD/lVlRtfTPXZBmR2vqdfy6NnkPmXCWgMPJAVE15hhw9ocqde208ZI
1DQH65dciDKmq8WRUgYd+GaEs0lfICrAmFCAzgPrXR8YUvU0whH+u5asfE2vc+oPmUW4tNFh9WDG
qH0rmDS/u5LU8unEiRL/vws8WBN4FW+KETVtFXcpzqZbfykJyWO2BXdSCekNb7kd60+DZBWrObKn
0x8VQV2QrRqszajS4zucFptj6HAns9VklsQSq+yvo+T/DtI1j/nhOwVqc6h2lQXmLoKjUGqV17Ab
sFumIQTx+rKSD6P23pFJUkP8YYzMmaYcWJbSiCvmlzSGoJ1rNL8ge0rrMaHZOQHn9+9h0DU+lv+R
aMx6kOtmKQsTFzAlGabvWj1y0Y/YBlq0JidWeR4tLl/ullT6gLrROPjv5nNyAEYkuxHfxi25FC4c
DqIRoXWMQmKatb9EtK8tzRKU2tRgwdwzoVHpiZRTjYddk4TelbACvvGpoQADnQOwA4YC5JZ9y5ax
NdVplPPLuBl5gYDkN4HqMInTUnP7HmudRQKCd+ha/bkmj1SM4L6kF5xfyXHZfUnGBO8DQCyM3nCD
VkGSnO4gglU9EnQ4vNlx7gQGCOFwBn9p8lGzXX507WAjcCL1rfT5usYSZdWvTITtqR//hKwtXDT3
lfaweCn3qU64kl8Z4kOM0ZsVz+Kr6sHQLXse22bBDxxBpXsrpIFK2QVyhCGS0irCAkIm4RutlBc2
TgvhrxT3WqrSDEmp5dxSdhZqHP0MZm3Mktg5EwSYRSOuc2cRTNDbDu46rkPDIM7YsBVY6NoLAQtE
tf4zZh5kybI2ZOC/iHiqOamh5ECUprnORTy19a48zaQSOIHkUJM13kFX3sC7kXvowKIdZTJvuWXA
8jjdEZmYIlL99BFb4jdj3GI/u2GUtQUJOaGSM4dQGB6XtrMra/WggamxUsdLtMo/NrzDby/MTUb2
R1EEq04dU4Mpo3HESRhhjg6tbeQxQK5hnrZpyecEvyksuMAZK7i5ZcknXJo78JnCefhIB0Egfcvs
P5yVQaIYocCKOE540ay1k+3e9qkw7TVkujR/ZFEkgNHsdr3xG5se0bHKByewDKvgIvnVQag8omCm
gTRJ5V68MYcUHdAzUzynqchL5pKC7BCMg6F56wDsoz3zxI03g/yH2Jp6s7TmRI85O4BKSdVkfdoE
zTXVj8PzLmva67Ci6N+uFbxD8Dt4y/mvEzolTAUbYrQGGHJwmNV40Bi4sDDgH+3ioZOpHg++XRKc
I4fOZV7SOZsp4gjrx/9MqFiEBzh5dikS2cVw/iK+XC1R15mKCLdYRnV6lrFbQlNqdYgx0V+rr5dw
aKF4p8IryHar2I9r6k8gl6/PP/OZezhQInyB7ZJuCn4s8vRA7e40Arl84wSFWBfZSeq+p74zNWbH
dOREiqogCagfgz4xNblmoGB4VnQMpUuZgCFPzRmuKee3gqX6ehZab7GH+kKW2TLwE5ncpefr2fXK
RxQKMfO3/36pOqEMnthqPZawwTLxE0Vb1pKhBjQUYPB83fSPnavm0+FGyfQuxiDsVyWZY15eC0hu
mxtIvO1Sa8G1hR7wUEcRD5brlwMaB9psO+0ZqqfLaCEUK1s92aGFgmnq59iHrgq91QNJ9UYkxGjW
lVXKcaAB0suDeEZrc7OUzVZdZox8hGo4wXJmcFqxIuinrn3KDqo0vz4BkeRX0nlcPqf0aiEPS9Pj
1uA4x0B0BX9TaYMx+ZEBSNoRXqmkXNOsjO3wG2+jKIpX8lF8j0T40bMG6fjcO4otpMomJcTssMgB
GlPKUBI1kPEOdIGaueN2ldbwVyrl7gzPNE9tb2dta+BOwZPxesKP8eiZ/xRltQY835NGofjK0SvW
Ou82VUA6hzI/MNSbpFGXyYpzO/IWVFOVhE4YkWv3AyIobg2zys6AsLnj7YzHr1lc1rl9jmzaIXC1
sCoq6e0nYKAM1zBWo9hgH/fDjsjFAyMtptl2qnMZZgeBN60/PnlzzkuT57oe2NV7aYeM5FYWk4dQ
b2mIBFnDkbioNlGihI/igI+6Q8srUDcXlXiRpjPCWPwnpxh+We7m8GxpW5Jj3FXusNG8gCpwhFGd
/mSCD0W95zbZO48VVaobxzBju+ywjR0NAv4kVZLWMdbMY29qEmKznC8RlIUs0c9Rp1CkrcsX28DE
uDtLHtB1Js0oyWcSZ/ift0FmYDIEgvl5kd1KmQcxbXdLgNMC51vpFZUHiCKSVw3AKXIJPOhB0eOY
aH+oIGlU6/owvHUP4uJjwSxg/w69UFm4edVZhnpT8yDpsC+YZ0KN//kFugh5kQ3Q37DU37U659uB
MwCGVdalrAywG63Hc1jrf/CnbyZRD/W7cBziWo4Oyldsp/ejAFZjSnlqpbO7y4gSa/Q/kA91/hMa
gHaCB9E3y1SnDgXLO+Ic5UZdx1PTRtRIZEr+tVufu+YCOeExWAHupLv4B0DLNdJLjOZnGgO3jXK9
93IUDXJDwtpsHZZXAP3QIh6howf65bT6EoiY8kkFsEWXmJVUrL/69cpZsSuIm3hUn9tCYi8zAhQV
H3RWDKqYT4zZrtImzugW8v45ynhE9zm0OHqmQJPQOI7zPUZvLMRRdhx4n0GhPI6zEZU5Dbj04TtQ
ZWj36gKRSQjBRvhOUw8HA9jKHKLv3NBGMBFOh4MIt2TcImVliEI6GB45Wvkgmc/u1MsrGmB9hjuG
aNS405x1ob/M/xnPyb6WI9Msu/D3Va14OA/Sy5WWFLWpqj/AjuVPjzihKFwUVIrxePu+2J6aP5wj
IKwxWH3GU54jxmSg1KKMbAPpl0E7s1FeAfoRhRECNTzp0IZ7T83ol759mXGVV8gjqgYIgnI0L48M
cVXDILZBqZhViFSgOTfR/i7wH4SgkUquw3pxFCs8wkMsO79EZRS14t+IHXwSXIfXTZhEcmqEXbVS
CpakE/sNIz+2P8QeouEyDtxnVDQ/+ZNuGkX2bij42gjA1enScxrDQw9+lfaGCMbS5Ws0MWY2frkV
lt88p3tBnmOWM9X0xWfFkIUKTgAH8F0IBCP0DNpb57S7vN+XpunhTfBzUJztlZyHfTHbPvz7lW0M
W5Nqea1VoRaJNKR2vbFmkSzhiFLRgKhLVrh3pZ7iLY3TopMt3rdgEm9MC91kf21HvXol1Sl72HOq
A4AVqlbK5A+DRF3uIPIJJa5LkGjP3DcGE9RUcQ6ox1EgQuxOsP/nm/g5tToQu2McE8Hcm/h273sO
0+TKvcu9x9uOlTnHkwqxey0I4qr7nfTU/hbuOfXkfNxvuYP7nlt9TufspTvSLBg2FeH+pkJKZ4ai
SllXoddmZaZjkIjYawRsnJLmBBdjJv40fOFYMisu/PpZX73dv5oxkCLU14Xc9r1spnfAmiwb3n7z
T/Dxyma2oibVe5ifK5tvF0BaBHJB9CrqNpsBlcld9CLEOntS0pJEcNaiT9dFfHoaHg7SqO4mLiZt
gr7/2YQ/WwrK+INGsBYFT6n+XeHEZdjW565p+yATJQgnxy84WIgMZrkh+kJvraIuATqYfJz6Vyqq
pGHxupruKm0osCSXdXhQxqELvV64zrFT5LCAWGoTB+bZ1+KISdE6sQzBLMhTvGvrnZuGF58g3N1m
im2G2XZTgiCLRLf1nUqAT9/NY4+HCfjJiqCpAxmg9aonGxeEQSw6HefBY1meG7e609Rz3IBqZR+y
7wre0H8dL1ATjoX8ujNoYE2saueQ2QUfm9VsNeThxpcV8vBtOpj9RNXK5NY+82prrliTiRvol02s
Ti4iYqkhG9UXeyA1cKbdZOnGkP/oGM5AwgMDcefTWG1z1qiu5f9UtT/Dg9JUNZhf3divbegxEWhv
w+ipSICGXSpN7NlvpMUvfZzlgpvLXwxuJvpNOlN2iuLJSLd0RTyBifeZ/9iycObZ1D95hFKxHFEh
Kisz7DBUODZQLPlwItg65teKUJAgEbODC6VPBWc0CxLcBASVw27LlLshCLBW6/0XnnI0hc0fFW57
yGLl08r+Mr51sDU9B6jGullgELeDoEfnj0r64wmL4pw5UcttGwoJxV9T487CGcKVmBU6hLIlK1am
NnVv1D/yyI9AAmIQv08U9U0XDPBKhV6U/6l/4w+PwGK4KanNBymF8ZXcsClCtkahlVuVlOGJD5R9
A20PaMf5v15pd3JdN7cKwOhsuJVYuUKxMFKCPMwPm+7fhHF1VLngrQDVxxbe9kDWsYMQ5/4nglTD
+7p4hdS7LC+OhFJAr5rCklsTqtKY47Oi9LKazERH4qxVybZ2xv6KRqDAmTVTe6JXYnYP/bffcIvt
9o5w2CUmk1UnYwLdQ2GimV2qmHQ0Qqe1Wc+S/gQ9zCOEhS3chiVFKCUAtRbM7KI3bA+I6xxoy/ZM
ZhlEm5bg2zHSjWZpiWvMdmfxT4YbCsM0IbLwXLLRoK9oFJ7YpWHjRKiXFZPFS1cGrUQjA65I5v65
/MyOu/0dw9oEO2Ujs3wUdUnM5RK5sr0I0UqFgK9rQnT6s5TLPEgOZEJ3CtvXLBipiTrjcv1gyC2e
/3J7Q9tM8FghT9mXKj79lkuF04fSmvMVHWGr6SUNoclMrtSyM2jGbgpzLwvogy1GgCshdVtzmj4d
xnwMjAqASy/Wo+kHUErh9W/iwUyRHHYuoUpzWbhKwiF1z6d7Yb6gu7pF2R0upgsbR9gOeqKM789K
OnC73KzHqeIQfnHciDnMr3sMfP4oYflFldnkkK22zU0WgrOX9exdpdgCSwH2xMEshoyQ9f/SCy4b
u0BWEbBucKUxCCfV231u3EilnFplcGVOMroFB9IKW/6AlSyCHyL9/ceSU7QSXFx/uWe0yPHJqqWi
xjOo0lwkMkryQrDCkH1x1FsOqjRtm+XB4c7IoAgyvbpHFyEAgIygGY269u3LMn7WpkXky9VywZXN
iYeeJa+ta734hV5QC5w7muaacSGjRriNmhR4njvcdSOKD9Nhrevi2hlFaYbCimwmkiLlSXGghqnE
1jm8yLRZhQaXPXKa6Hhy/NIEgRQvnUnhizPynBPZEtlHy3Dx1GPqg2cg6xfWEQ7VMF4GmJ7XEa1X
/icRQV1hpNBHyn6Emrf1vLhppvQGX0HpJHDgbCGAPO0z1wDEBKSASirEa61sHUpf6Tf+6DLhcsuH
0+9qIxU3uby9HNR+Gf0vxKwNdkH2GkjUxOfAaMtsc3W/B3ODhycmV+f7jowk+pBGKciODMgVF9W4
HUWlfJoq4YE7QsYI2SDrif9+TeFlPw5+aoNaCsRfJa8FHqom19QJAeGbXqj/q1jFX6bE4ofRBvOQ
bkcn6Wu+OInMgCSY7dKfaF1CCsebNOgDNkTRw481bPmEf/DKUw41ib8VMT+m9DSyTeXeXuS9jFg4
PFbVxDCMwXHd+aXQtEKE1Xt+SlZoWYDfHwYlj3+Qe7dfDSE87nssj4O1w0RRG4LHrzZ95nHORPir
nanq7NButxnSznMPokrY+lwggtdBTL88Sh3GVV50RtSTTL2GMzdo9wzUwlZiGVzcm7UYx5dwfUtY
530s8xmoDLRIL7idDJnOx3/j4OefHamM48PkYDEdvU+W9O42Vd0Gdq18w1cgBFSts7UmfpiKGvJF
kOksO6HfPV0WRviKdc2sqBgx8p/SxEDasFYq9zJsvgb/mlog39EWbngIaJYjJZPulXgtdhS4Xmfj
dgfiLl5NUR0sM33jI/xqRIoIYv1nF0V1+5aHlAac7VZyJIdi1uaStE365OSMSPgNu1R7/ZnRG7nH
AQpD1/RzDicx2geXYYREoGZl5870xoExGDyeCQBqWVRpRu8Be6t2jdGeXmCGJy6ft37Z3MCRBrD8
Z/8K//s0fiOc1xdNDUMbic6xTq8JoaFiZplU1veqhztjcAYWwzVtZBICVHtP2+whLZHbjNoOyQvT
YMJ9IGWYFLPJegGE+mFD9qxQB/2y7ka/H0MuOcMLFYxuRcXBbHe1WAlTvsKzII8k3jUQvCGIzuG9
x6NO4ZB/Iw69Ic1R4fwwZq0DbCW2NeW7Ctbk6WqT/RvAnL8lIIRmcjjKTDYMacGazQtMW3PiDtTU
FMfq0hGE3T5L1+yqbI0N7/AB418sIN3dyuHpXKFwNidISc93eN+qITXUpC1ZNEYGlzIRbPcrKJbV
960DeuTdZOgym/BSU4p84V32Qdj5A6kh4KNSi8xhLfYGYwJuWNZ6W5LNbdDKog346D6AItDkr+CB
8HyMQ/yTrb9Xwplu5oDHXOAf9mh/tyLBm2icnvu1zoTdbrW484lPCvShOpxapxNqPJ2gUiqZvJnH
XHTUjipZM/ee0bggpV5ob/U16EDeMUCQ+Awj9dYAMaTUJBYShwuRDbrmvcVE+TRkMpqOF0aXIvnw
uLUA2DajJBEKnnwsRtCeKTeohtCOkhUy94Y0lzAY18wipHKCAPonnERxkcl+EZ+N4gA8WMb1VXd0
wRx4QbcvLWF3nXFv0Ll6prMsbiL+e0mfnbxnv2TEQ8WXVvtjYdZc/6UBHIxxIPqDXK8RfEx+THwf
e9lAZJwBYiL1MBhhu3cq9F5zqybA5LMBc8dYpAg+LaqeQlR/rMOkOOJweVtI0EEzaXOZCuODAQgr
RVKtegwv5HchkDRb6yPD1RmHP4c8M3KmWiIHYUlNFQIh2TPiclzJqJgpsNRgMGkdtbSV73crtw/D
z3yeEevh0AXVCVCGBsultf9AQVywB1VAvTyNXz7Kl6q/fh+E/j9PlecKbrH0cxx0V4l7PU2VhAVw
1rCiG+hs3FR+lXB6jdxOZEaDheAXkiPcslek4Wzmq8U0ImXP4tBzs39p2LtoUKVrwn1dg+KLgUyW
saxYPQXI/ahCiJPHrP9EVtbuwi8yP6/65dXyLAf9ld0ZTsMUm5aSl7ecuz7oW+T7cCV8nZT7f9nL
gkZh4MfWK2BAozc2rRnHkzCVE0+Xvu5VilWoe4ihkpanzrVyLowAlBhJejUUbUoaZOjyUnu6CiJL
OnPtvBJoQjL/eydeCtaAufYumdeUnpRy9KkUs70dCNwZHJltUCS6Mk4uJZ35Tbx+a5fmxvbGH+90
8eag7vDrDpqE7NnDFK7hCTwE77tkDBNOyFPwkyxVVi5yvMD+tajGULjNcVi3XRrZbpclxz1693V3
BVWgjHeO/lyQRFjVdZwom0Azvh77wcRADZk+VnLOzYR7DkoXT7+J2gktVnXYVBlSOlQ35ZjObgRF
iJUyFm0Hh3yH3sRZot1TUmlip1Q2SUdXADuZOUVIDurVBGfJy2OotIf1ZHmnK5tMPqMLoOfBy9iI
u1aV9ByviOpIYaGyJ9DvUzREyqt1KduFi/wvzv1dZkRRKHa7wBycXqd/5m1q37fZ62er+7UrUWvN
wLfI1mx3QIwMM9rAHZVWgc2UppWf8W3LwVs4enzEJthOXVzZLiNyO0eqKdXY1kh/ZUJsY77SywZd
z/LvdKihuQdsELRKqdXLfAwI5aTJKZTFoTu0x465AfltbjPnaH7M1ItZkDBO+G8WAFRKCSXEEOMQ
A8FNjzTJh39G686Nzv0sdqyA9m/35sqe8AY0QsPvDrLTblSfjNU+rVWc2iNQEwZw2T+y1lJf8jDV
qcQ7PRnmBOoXMUBjZuwPvUTsFAQNM4D3qrCJCe5SjIJ3X0B3C1P38Pif9bIGh/srmgfuAJVp1hY/
HZDkk0w0++ncW1eGIXpcIUyNlH9nqlvakbMu6qGGUvtXOdyw/BdqfSBFh2Hdy1u+KFo0+MinAw1o
V/D69YQ2kEzOJtWcsqlkU4TkfzEWtVTCACI53dRTIQ7Oa3NSVmt9vJtye+RfXg2x9YfTRk/IUtxV
PgYR410SpzlRqh0x2PTHzvI4pmKCWM+gq6rADWuy0VPnb9y05qwuDW7YJqoxZ2TYcKazynf9z3K4
3xCjHbLjHlIUdmRDZEbpFeIZH6jzFm5jb637wxTvFICZonCdoUX3n+T+VkwTclTqewBEqCVA83HV
l9EAM9LfR8Vu67pMFqVg7R4FwwmCH8Kbmqu2+2Wp8eK66p95CXaEvwEYCeDBqaQS7uBOizRQMGwS
X+876IlTJEfPi6a4F9kMuyjJXxr8DbxxqWstb/LkT6SxKPBTomP3gMJwxw1VesCoQYNPn6LtF/Cz
59RHy9CniltmPQPM6lw3rTQXhH7DYlzA14Q0QKLT9ua/ZhKuHL3KQvQIe7IOb7hnSePO5AfG3PLO
wV9IHaGEY/OQ0xVC8Y0fN+H+V8uKbqdrwOYT7xTtb9n/GxkvVgr7Q7tf3LiU4l4eIFJpfIufVGVE
Ju4QExLgy316GepZe64NO/H4bLT1fz3nebLpPl4+3g5Pf4hoxSWX72I93u49GOCkmUdnngyy/mFS
JE0wSyIpTICr+Zlb0/WrUdrdcycD5PIdIVMmB+LDWuqYBkKgHW+a5XGjk9C0+Kso4ciA8SVC1JQO
qizWIfpMah8usWkvPoTIaPsDbg4aPFC4JF2nZma9zQU/uDwXhu59xcXJOz9OKency3+xdo/NecOe
ezA8Q8VaWLxjukeIAjYCGPWyDL4+eqyTpiglV2mXs0YMjO5HPIc3ry9quXfXnbfzwFq4FanuXe5z
rx7hgsqiWCB0e2aEWd/Wgi/KJrASRE/CaoF9NAINC+xi7vGl5Nw6hD1I+scGVAldVbLutbtUvqBE
+ViRF5Q1X6WIOqkAYhtL0cdJxIfK7Ln6Rvg5tuiujU3v7u/t5xfmkZlb3HC+okp0d4b5WPDxhNy2
RXB+FZbD9n7X3UO5/mI8ylzA2PiwCQ2UcNZtP95pX2H5iWd46Fm+iyCvyxv6PdOe5Siqjf4MmfTK
li7V5zSEnvw7MP2rE579KG2PaCSPXaHs3sOxRRZ76a8n6hslfNHkN5x7VuuwYNCtmnl7TD5Ag6CA
HyfalhzcnPGetFsJXj9trhFi2bXIsqmxsLvmDPQSuGYYAP0+fOxVvtl+YH++e1kTxe7VH7v6CAc4
TTmTYJIoTw08nR9bzsPHeaKg2tAIMxdd974fg3jaBN/985g0FzBcl7Hg0NQkJFfnNP+vESCCzWSO
uDEdJCkSHyzK7x5pVNjLRpEujveZtg4Au2pzFPjdn3AlbKf1X+sEuNp0/EW3mZBwdWuzJV3uL5dl
hK4DNNy+kISyNV5NhARZwx724wZ188f8eSkGtQFwA2sKOBoQc+uonBTfp6pJbmiqX3c4xvSYVyh8
5iF7LyG8jfcg6z6rtLgnjyIKOSeCwA+yaAuzsP2c2G7o9xpiEu9EAomHgWqiS7ky11B2dEjuJgqp
wcWuoMDEyvGUU4RS52jrgzmzvrmf4RLvyy8oCV8Jz2KMmd2WyUmCmS9+zWvivrulxAY0DYENV8Pj
WbcWvf72rCRZkutanFuX/4IzFILL0UOZHvE2MFYt70g9RCzFZ/SWKX/6VGYD9UR0sUK2+YlBoASt
zb4iMMxKoveKyrJ47iSaYP9ElmQ/CRU6wihuUjvXV83uiobNVzBG8J+oegUGvWkVQ2vRfs8f8Obg
dQG9S3l4FyqH+ZkOmvpTpNBY9KtZncX+x9vYFJaAqZEWAaU5nHL8t1i56w11wweeldyFeAXbSDpl
iwffMEK4+nbqJxFbcoH0NKytXdOqbdty6LVvBPagwFrpOm8L2uUDnNBcIYbt0SCIhncLy9jJQfPU
O8SR9rsxAXhIsCZKmWzuyN/pzVb/7lorMnDT2QoErfXCyvXB5R1vYKFmaLEZgX4u/FQi6/pAZ0po
OzfJpkmMmwbG4c8E8ObiLQkzM3Hh/aH+qh6oftqbedQYkIHH/WEzcSAQklGdjO4vVOzH+q+anXoS
NUIm9NiWlO/HzFES/QCIT/lwjFdXMTbjJ3OjMkIu7MYaX2VOZZAeJ/jrEhQlC8SnGuoYecCCiB0Z
O6TbxTsLNM3nSNhtj3H261ddB+m0eEdL93/+QF+pPwsmeWto+0us0KNBQCtmxiUSN+B0RAh8KuyF
FP1Andakit5ZYx2rd/bf2bse6ROgda5fm8vUv0RhnrbBgN4YeQBzXVEBOvsxtSHOau8QHCwwlKN/
+6ougLuFf0hL+GO0SnfeeeL/xG2nL4xsgZaqXQx7ONwyhIkDkGhe3983FtdnqXamhi6bo1wFusBD
b1Jnt2udRa0vXk4m7RIAmGEgH8IGXmNVwv1zR73yCwAK8JnPKWMlcV/w46l4AQlwwxfK8JGCJGki
ioqtTwdaQkezegAUL44LB5G9dlKkoEkfO0ZtdT52kbSXenvpAEVckjtQsTS6cJzUPFCXBI5GbVHQ
p4OWA1WwX2464Xhb9PbS/9z/DDS4kABB1oSUMQQsWzAXE8c+SU7RdHy13ycuIQ2DsQ/6NdXPcHJk
iu3fwJfZs4Mv2pJUnV7QrvE0UPwvXK9xqv9cdN76Aq0Gbm1FO6xsqOGOm2cY68xRQouYc1/O9a3l
rGVFz2Wz40wwTtMcTTtnNo7S7gkPuNErIdh1H7j8UmYhnyPa4f8/Qz5jXSltIU9pFrJk/D87c5lv
P60e3tdvIneivMUtTbcnptVHCOiy8qMGPvs0c/EamIJSFLwBk5dE5YvjD/Apg7vckg2JgICTSE2V
uf+RU6pD6X2o/u49beW96F5c0mbKS2Z8dG7k9do/8RqG717oQcKi1EKV6nF2v2tQjJveyfQuviu8
9MdRWRxGTHKCmRDTS9uOKOrYZfPh9D43kYQIT9KG5Oo2uHUT1g+elXor87Sd6s7GtL+ooLUl8qAc
D0q57o0QixhsqEwfOGKlBfAmZKMZ4oLzOoHuhEBg4tLuoK+Vr/MNRdACMfgwU1QhuMCNHEuhMTiB
384k18H73sX2L9BQbcQ+G2zJQTuXcLmlGr8ypJp8lolw9LxELUt6h5vpvwx9wxerkuG2DBIBLI9s
hHRLynvwXfAAqzJNFFcHutEiXSR11TXOdZ/00KZs3xvIXcJvuL6STyJpBrqHjjTaJznpwIHeVbDz
FVZCK/EBDkHhPoP0Xi+BTewGm0mge/uEAg0cx649LoI0yRJf7rcYGykT6oWMuY7c/RDYcr05J/vs
PciSLrYX9gEK3aKV5/B1wJ7TATPjx3neKgzb6t/TUUiypouxblk74Fgh3d/U4+80WiH+CNL2P+k3
7xo1CsssptQ39FmZ4H4MdOlUapQKO4m8VTgLfE+PKjGoebALOF5GBDrojHUz++NfQpl+tqcuv4r7
+X0UbD+CMFlvZGpAdme7sLwwHAx96m1L6rzSEyPXOKF9xbo8wz7E0aHzwd646DmwC4gOA8thtx6W
ai7eUxk7a4GALfOwvbsEK9inGXRxtLogtc3Gm1/0J6+TY57e2EC4tUHIXmZWHBHTnecXWryfW0u7
2r7IDso0A8RMjuEGP0EvEUpC7VEeqF+rcmEWzlMubQzsgSV0Cyt3D2fSL8mVd0SyRG0zHtsWHgZ2
+b4T97tK1NvnT7F8dQ7rZe3bSXP6JIcOxAEpS9UTAUaJjLuxAU+6xTp/AdVRBtx2MyC5toyp7dEy
aK2ELrzmeqvd3Kgb1493gzuX2OCttDNfdlRlAx5ZnXWrFYBmceuYbMnvrhvFWA8lPbSoxN+MnQrx
aV1aEFfwPLHF3hETJb1AIYOxiPfgpuBM46wuEYaN02mFPyTOwrC8hKbodmfK9rlrCUzl6/KUoIu5
kvtj5xy1n6BRuVHge9bhafCx1dhJELFaV5U0fzXfJE7rtJ0aYsmqXngKOKPvyhx7+gxW97dPfxHC
zPqST3I+7SmF2X6pimktl32ukgq4ec3ecWZOrHcTz7D3ai6Joz/Qeobhyx9ffFU+5hVJui+JpPX0
jxlvZpTtMLQexFOPkJUuB5s/6pWQ1fGcWb6VI0IFYPR9NEfp+1gQ7izzyusrY+XQo+GMsUb4CPWo
xGgy9MwB5VxLsCeZym4t2h5ZKAdRhkNEl/sw27P5NePyWnnbRL4bXIl/XHTLGz+g1y8db5EJswJC
8TEw1FdGGMBCnRxCrCqXxqgof+ilsv9EJOjOynwHhXwAPo5jlR1EPsemyDEz19ocba8Ln5QlEurg
L8EwWW8u+ZGJxfXH3X/D7/indkGna3CfFnDPmIBVvAxecjnEh5NrS4SD7JnGAu9uyr9qo3iY2oiw
mjQQFDQAcbsMI2mf1La9E18PIeP/hgLQ7IG29US+NGEHIB+s/GwVxTwJNeKZYOe0ayRE2wlvU5Vu
csvX1LILqMNYGWEgR9trUFDh8E7Kak+/XPRhpOmWLprXayKwA/jDesmhLNbk6oK3RrkIZ9W6MtAd
fB+R3/jUnz+m0TPUVXQGMD4v9wnuTrAAxrSbRyCQUz6ovY/DqOHVGFmrTHmbHA0XGW8zUHu6SgKy
J6FOeAzQOAvohs9u3VOIlHz1l2+3Q9ETfy4E4ZqOdIlFpP/wxYgh8E1TLkWDvEQ7Zg08ePnOz1dR
5cFcTVZUYB0PlZ0NborLKE9TSLD2b8y80OxUmZvM5oy2xkPyEp7Y/1KJZCmHN/yYuAh52NUe9RHz
A48lCIdzBTedMOEd84sKwfXAMMF4ebJXJz8h5MiAssTycfcqDyXYC/pqUjVDNzgWePmGK5TGjbd2
E6mgB3cR8TmLVKhYbizRYxt/66RsQJTKMqXcXkAvLbYSilPrBflzYMFTuJAhJxVzBahiCZXC1bsR
gS5kHMfj1FMJLSkX/BuXRSB+9d5uYNaNszTU5ooyZWHU1TO0roHkh3G/nz0v8T26jgNGVrjvTr2B
epSPwECVrbJOlnKsTcz50yrWCLnG1P6Kkmavru40Yyvn0HAzz5dKTn2upM79a4qoGdKAvCQwsopU
GykYE9NCBdjpU4TmdguKsQzZqRD+1sbGw710CxfpV5X3XeIUAxQAOGyWy0L8GOZrISo1ns0FRya2
vCSIDAZOKUD8LKV+BCFcmH3FY4Ez2bQeXt65D2V496Z6iD2MTAprHdGjYiz1Tkh8TG3yMat8dUNe
pPH9PMhWufAnZMIyJmOu8qDNwnhgMSSGWk5BUuEPinqPvdnEfCVSYAJ+0x99UKE3hUILgw6VdiHo
QI/yVO1lxGNPY1obewLc9RccfEiOvD8QydNqywkkIcl3sEFp3M0TzICx2ohUNwwhp7X5nVF20wUM
KdFiHPPrXWDaxJJ32zu2MIJMs9g/qmTEOlk5nxH/iuj9G9tHJ0+FpFz6x0mvIJXtoMbjmgu5dQ8J
P0m+I76923slcUssZ0Gd/iAXZMmCPqIsUiV3pJkiblClfeu8EZkVfHjabwfYAVwDY8vTQCkQCKfc
1m2hdsbgnfdLmRWu+DMxFMzDxs7NUssDkxuqu1J2s+2LvcbSW5tRQCUKg9u6ElgNHKRyI5M3dftI
981cLi0G709rBkbRuMzE6+Chz9PdiOruDG0PdNIPzVT6a9JD7sXXaS2k+xHsJBqr8pDQ+ezcbG99
mNCUy8Rb+DcryC1Och/oZUy8faR+N8POJG3LfjQ3U4Ko5NYFnP57SAgLshcPP287nvynRqYXV5io
gIm7qLU4gwgAdjQZXBRSIi4KfslyLfaSfUAvT+pSTXoLvqL5LoUdQobKJ01yH7p+/j2DecEA2PNU
E+AffiEB446cWQsGrPiuW3TS2ZYZgfVcH97WwAl5DKayv25qL0h3nFPruv/qwkj4IlyGEd1jEkzY
fKn7BmKMj//Nt7uFSEgsOk/HMoI93BPXYtk1iyTrWR4II8cX6WoX08J+XMOp8pLmPiK0/7pwO7uZ
9Tr8ohBFgiEs6UdTJwcC6CBKsgWoclspLnck695omn/JX5ORdsS+1ucvsLJm6o6TqvvFRpb+nB1H
RlXQHYvlgPvUUMTyjXlvWaiJMwkaTOw0A9cz0h/5fjdLv2LazKRLyTj+PIvBTdW6fu77jOlmEJq/
bMLM9yh842XGvkKVxaKHPJtUvGGOuKr2fqZbKlxcchekevLB/9KoVnxxJlfeJYGqvOC22IUv+ghU
9nJpQ/W7HMBU1W7E5jWhjtndIk3a+J+wjxNUDo7IAlRbbwlpoMsPCV2y3RqFosaxjgaDcvt+5Bfn
L8FT3FjhptNR5TGEmsO1LMEKyz9gEs8BpeFws8iYNtnxeEkzZ+aB5el8otKk1fKJc/JX3WEQDcru
G5XCp1PZbl/+0bbWGHdW/PzAwFpkpZ/1pJ4J9rYBETA1TVZp3TC7Xx42rZ03LDXRn5+bs/HDjDoc
Q6Q6uUP1XHD20MuhxDCaiktA7y+TujGrhMdH8Qii0y9PBYcUg+jtgGcgNnedL0EK8W/1gTLh+1BA
17wQynCd1fJYFD4PiQ43wmVRPKaUUzGp6Ms2y3ksk43KfsxNoZwNI3QyftsUWitE8qjL9xoTJJ8c
EAW8smW3txXz7HOSChZ8Ps3+w+4zm74G/6q5oxkpKce703cL5ilX5+7D4l49SonimqZMihsZ63sj
GzLQCUy0Ssw1ye34Q6pZJe0x0eHlpNHSj/tkhnpmaZQuMo69x8zIcdV6iJ29bXsaFxRzIyWunVmr
gmtYzdWkr+KB8Sq9G6Pz+41/QiyJj2eeTtb+9Z2NsiVVwU9DCwWmN35rQXKtXjjNFr9QHZQlIzhD
B4zJAtCawEGt1QZ229SfvnP5YrRtHMgcEoGYucV0xAzXgtOdlPDd7STvZpOwH6/6vow91UShLUbE
1dJFVOl0yFIFuxq2HzQYUkkjxzrHIxOPjCgZig/J+qt1GM5g39QxSdyiUjKvd7YgMnZTjYWZQdPK
h+89HoITSHFlUg8VdhiCgko8O4otiGp6YOaL3BroQb8MufEO6yOgjWPT9dD3cRXPv7lCqkrCTtWN
F92tWZFR372pSh4uwTA1KL7PyL1aoNqHofOdZPjjtZuyoXvh5sv8K3NO/eS9nAWbY27ikLU/k10/
K8fSP7y4BmhlQ2xs84huUJwkY7Ks7IGOVgQYGXffCC5atpV3stkhnSnJwl9JWU8KMRK7NU6m8s/t
5jC5fv8QZM43PLjovxbEBJBIimhzn6TLCxh/oC1wE0ECYaN+zY5DIptLSXZNO2MZvJDa76Q7mmcb
N6JBPZXFiOy3tuhbMjY/LvKdDeCv0jkIbUBUwdK2Ok007AKsnbE7KnRxTlm9tIYG9GRKXL68NMZZ
8lgYBTUaL7nR4/HV0KQma9XBRT4/MtQg+WcY136whV1Tc1NGV/I2orQZ5JgTvfYVemc+fnou9D0m
EVqdDVfaE0pPi5GWakWZVs6wDqTst4ILhknHp7fsv1SD5024tThLsg28+F0SIYv13uHDz/SLYvUw
5esec7WfUAyuaULTN6/LEvAiDkYRwDX4PVTpkPYPBcZYMe8o6tAep7OqN2LMSNyPTD54BgRayzC1
h9YQ9bte6LvJgqDRDwi/Zeq7byyADXkBV85rlmdPfQ2m1N/cT97sQxloPwccfL4Xp8drIMUKVpyI
lRBeTwA2KOCWQF25QyWy6VoAJdocjkhFObxGUK8fo4ISpv0cMwgc/vHoFb3eLZUPRvxshPOwJNaB
KmWATPoLBYxYW4vpDNFnANsFqxxM0RcfqlcJGAqutA11S+TlMKfmrkQVMHuSj5jzYVvVa69vCerB
OulWZrb/iCLYfA8r9jkRrz4jlKGecHe8X2TCM67xGcJziqQjZB6iyQHhKksdCKWg2U2j83yHu5g/
8iDEHRxqNULdVrBKK8a9FhPWlKZBTz0QMNBjQF/0/4SMqZ8zOH8UfghkMcduEDtmWj/FnV8FATv2
9V80rdeikDq14hayxQ54pyiXw8b1OPipQ+Qq2etCC0NxvGY4EnYjO4iKyXI5RsXxEk980gi1dMHx
bbnAegVdKP1awciWS8zPGCB1kLjmGqmjCF3/TwKaGTZmwuQ5y+Q04+YJdFUrHLm+iUVWnFoSiOUH
xVB3GYgDQlcmNdW24cSoG+Cjpw4BVccM+vbLakqW3Bl+YdSRMuyX4xbW6GXxUZ7RXMDm9wF7CvrC
yuu79zQ2gc5jfP5nk2qradt5LpDyTAEHnoYh/YFDwPIg1oMmHbeZll66goNSF2LnEBEqu4YWpSJM
DOwrXofGf0n9MxrVkJAi1LpfYRg4Bjlq4MxwaL1QRNVvHOkNlbIj5geq4ydsykfGp1aDfXsGV0HQ
ngqG0yMiSL75zeRmsZZc/1BcCFAUwV0N9TtlLhaA1uzFeJExh3tSXP+N7i1r2UutHPBUgweZ2QJ/
MTIsA0ELZxdsEkhEmlolsbRWk0U6Vnb0UU6daN7roU1QtVGNBFmYEi6I8uxeFRmXPMGiujBQhjX/
zOlnK84zzvfizmHdLqpP8qL2F3Xaz1At+FixlH8v/YrHDyobq8erpa0GDQtJnmsYjXOrOBejmOwL
S/6wKHgIuqGUOtC22FvcEDoY6FFL9GpiW1EuUzgYQhVwhC2gXjZmYUvQF9XU2bDPIPWAA2IhvCwK
60HvcxGxmVPlk6lRnUgCacQacr7MYokrcmKaP0/5aJWAVpEgWRlkBFH5/hhxchoe3VLrb29Xqg2l
+n0LOK0MrHZvQXnj/LviMV5SEWCyigGBuCYr/6pYDZUSYyCkpPChIovR/SCGF2TGITWpDBj/N5jf
VDX81kANWZRK8kSwqxTRgqvj5iBQDuDbQAFBXvUAfeKUXYwKFZS1OG++ylwTuYYxcrGQn4xg4ylr
cNo0oJUyRLTCGZ4MkP974S6kn5U7WJv96K5HgD4zH4RM+IEWBhdF0Sbgzpv1VwFjsioeNmfsCKzo
i4JoUUpA1eGFH/Da5Tj8fw8ZqzSdTgLem5D0wQVTPYD72ulfyENUJiTz9vEFfGwUysOjc4e25LGI
FmkiLbpIdbMhFA+vTG5T1R8xT2zKuOcZA1Llu6cmM4HX/oxHDtMV2xBEEh+9iZjOiBb8OdcGZjp7
aa14WGhUBINOgF3RrzNKWIKdPijX7Wi4po+pEeVaeKjxVLbH5Erk8pYA6uLeG2kfsvVOc9Lo2uOP
DRyO699FfcMsyf/I4DMIKvGiu79yMjYOAyTcjWidBC/OWiqtJjvE036/ebepS+Oz5FaNpkdnOWT7
nyp5CuTghfiNgKdjHBWi6+Gaw6RfR8XMqaiFi1hnrCp4aIGR8zfZkLq32q/QqEJhJW1nOFKemNL8
X64qswWVVW1VE727H2y3Kh1MB/x6e7NmIhI5UjhCT7Gtl+1s4lxbPCVJlSejOILI6qjzehDzn8Oo
8eMAeg+XOBY45e9Rc3QvdoiXI+qutDGMRppAH2J5cQg3nBbismD9yCkP5nLIrKNgt4e569kdcE7N
lQc6mVAN9wiiJqXBS7DviGx/muvETW1wtHR2I51Z/LLljlkoeaqs0t121r/IJ0/6bXfgEvrekRA2
1y3O05yzB7gubpEYX78IvGpXaSdSkTh+2Po4gx7asY5H7hJfKUhKLCljoYXoNLTsZDWlpxZM9pp+
JHYVM/lNAXxCvcGNlSuxgCiqmm4nhEGkvPolENguVO2HJuSnxH62w/CbsPMzfxOaU7d8I5z8B3Tw
1vhtzv8oOqZW8Kc2LU/Xhc2u1pU2djnLBEXOvbDrUxlKkEBuLxAw/bAbv1LIILi/pn0Y0Vwd8/27
qpeKQqDDLmYRzDgvyI5A1/JNPJucOfY27lyYWoGD0Cextaiq11D07Ej6MAM3G5/MQCkx+o/s+6ZP
WxJagq490F+xiVX/bUxbvU5gNkmK+ocRWuzj4v0NZFZeppvUsk900LcWUKzEEMxAwjv1PcsBMV/n
K/OjxKOW33qCh6tLyiYoOX/w1c4WBVbL67+L61NjTbAFJ2k6F3/YrpLajtR1ENvJu+iP5Jdm5THy
MARbEN4Rk5+D2J5rFkRaiSAA5uZPPDzx7gGHW+RfRh5O/DMXfS0OJgtihJcssb+Ur+SrQSaarVDi
MpseXLMXW+tHnZ28KRh5XLXuIKiQ1h7F7wSS14K1+W0f1lK73et+2AO3JAwss68J49GFLT6ssXhf
TxQnHlLOPcnDTK9atdgEY8Xj+cYn3pU0aGG0XQ8K8xQLlUlrOOhT4CIf+jZ8MO834Y0Aj83lSaHT
qwXHBHnj5bRxdhTdknHE99uQoopqxhweNWmNC5CbPahWSiqcLGWnIQVEkCtGXVn/pYkHg+jX38lo
bj56FVJ5DWaAb8OdlZ1sq73RDsaYnU1nGSecQjUCRoAoZ+0zZmqMR+80NaipV5iTFGGbHIaxGEw9
ebQ8cWkzbgf9fqwW7Cu87xDMoDXb7nUW05yIazOVp91j+cph9e5CVORAK6B0/LD5OxNduW5zINTw
XdtbyOYxDbEtRekV1v+Ei8y6p3xOe6pPsFRj+zKM1HbH77iw/deK8nDvHtUItYuph93V6kCbfGa6
HO4PklqFmKskPmQ/de29ptQhLIdMPQYIFpzKJZF8wjbiH5UYbQ5DeOzGOD9rUuIzZzE1m3W1jFv0
Vu95HlfwfG6qZoQGH15cM+WqnpkAy14MXH7ohVknvapDioD4GN1fZ4z5At/AGc2vHNJ0ZdTNk03K
LW7MbMsa/x+wlZmnLeAr6NLtNUn5oNg9jXgc+ZroT7vkA54/uvZ0iEJe9VkM4qIG3pID+uL8S/nO
UpB83qO7nJy1T5VVmuz5qy9ZZpczMJoayDEEd9SEGK0E3OkYiNAXe4VxB2m0BJwu06x/CDYfPj/M
/6KobvTg+hrvvZoVFa5Rdkdm5NjcjvvyWcFnsC3glBRhIadenjoKvnrPKPvVwlpbs0MDdajPVtw/
6Zz+H18L8shMS8xINmH3RuWgvALbluTRu96o+0lOcObKidYwL1DurrHVt+3ixaj21bst5cKY7sc7
V3jYo/fFTM6AvolTDAc6M1UjgDD1LV8s4Vlkopj14yT/iyFYgYMrXd4ajdAXbwLCqAefoNjPUrdE
hIxKuaIDH3o15+ckZf+31glU7PDCrnhhMSAubIQAVsH6YTsGaCIMTZPjiSi/+b6dV/g6GzqBx9Og
gYfc3nho4Y1fjJ+wR4Y4nEsKiUN2lOxHW6e2izI5LCODuSRvmUmwiJwwEeVfSvWgnHrLP4DYkY13
W98PiE93Gc64lb79O5OCeoDTo4jTGfRfyUXdUSpIck1USQ2wlAXJ5jS6vjq0jwuyYp++rIcV0Ec/
G2rG11qhi12rWG3jKePEv62cXv8P+1b7J8umOer+2kvtnkAaulKGTxq7Za0Ww32SO+TSJth8nojS
6Azqw/PTyFYvB0OepK4rekAG4op9QPA6fbA9kjwoQvG7lt2GYjdAs1ubD6SqJsA1KRuDuOTeW247
Kwwhw/0IpBPEW8CLbMFXEgZUgvPysHVhjOLBnFkTvNVz9vxj3d5IcEGQL1oRb27wcd2uiP6SwpnK
O2QZvJzwvjgVaSUQET6KV7/cDOL+rl52aOZ+RKGSvcoSSmcg8gZ4Vgo2Fcg3NtQdV8tFPG+T4BuY
rpOs/uScpAJyqjYkAA8EIadWJcqhkYQm/mNAQl5+lmyuEx5rqMGgfxdWV2wJ95oSvnPg6mD4QfSn
05NWjquErM8+36t9uTcmKo+ZAfH305r92dBZhBYDlB8uy9gfe4rB+Fx7NWpvw+syenjDqNcrQwA1
V6u0YUwczW2apfjAC0eFZsL81xmgVZkf0D3CTe/V4vLPZV1z17Egj7JlhPCf0M6XfzSTU+5oz08v
qxZJG40iWs4+q1vjMJ+W2wU5eXqn/xwo85JG/Oa6dKhtbkTidYRMRu8xvCb6WL3d/rL9kGq1UjKd
sXIpqXSuNVxbT8kkQJ8gAu46XQ00Ostt/w60/Tuy1Tsy9mcmWezRv0ZISxaCVTr5naaYSXrYB8qU
yQjEGg8R+5HTEDhe2Fr3H5tiv7fDMQqOWoOHtrqi/PqTbMTa9yE1GUTyaMhX7yki69vSQjRos58X
9bJBn7znrhw5bMFF0TRp+a+HeWRftC4fvMbH4YomcBgQ3YMkujsJH52n8s1VAYMRm5wp70pRErah
toX9LgcRbwrgYXBYjoMXx82ORwTW1fTjeuHZlbmAq3hZwWYo5MDRduR7pcy1sGj5byvQeNQ1zMjJ
edtMQ+R8gLBGlNv7L9jcgLNx8Btju4y3ZC2b1hPG8A2DtT2SlEauxYB58WPsspGHalhdFzHxntOy
IAz/KxXRIsDD1ZDxbKi9pU17FuyVSw16xBRtEL6j6AlURzCza+P6TmlXSQXWDfU/QIZt5NGUHFX4
TkbYsq2Qc18q7SoL+da380WIlXkyJj3/BqDtW1KvWafpKrXwJTYGFNpsRAOZqziRrcWeDKuhuOx7
7tvExmql+j9qfOahh9yqjQKA+w60ISBdteCX0L3OB7oIKoVnHE16UGfrMENJjVveiKDo6PBGvkUL
A9QI8+BWf66p2qC7gzikwIDGjLyc3iPpzAhoJaEwDFEt8RObXFLK/+A8fq+xhy0/AjoDOoHXJ8DW
YMpTKI0mOl13fx+u52BU+neV4UPna6IQ3ZWOv/RaHN5R/Bz1eg0FVAkhRJ++tu8pKrJHXQ7WSS+p
SY/YCY1KQev6E4V8SDfvGb/whqaBWw8Fo4P3o3OcGVLFnD9GWaSNuFh/p0pOJXD9k9PZNYc/H5UN
Demsl5AS0TL2fi9S1JRpkSC7NKbSo7lu7l2U9RRFQl+hyfph5jH2SMDZrzCLXDa7yPulnKXjtd12
0493x/+ly4Ussnn/YDoaYHcxg766msBWxGw47eWAPnBlU4s3VAFyOyti6ReLLnUflSecP43WFgWO
JIhPWi/faXmhobSV4NpkUoZdbfsoiYh9XvNNmIDwK/UP3EQnrXm+Pw7Qmh9uZst/6YypmBoY05zD
n7uVOylzemLG2/0i5j+XXVmA5DTyjiM4b0bF6KaDk5ow06yExz8pCD91rL2h1Y3w65CLJzOFbHGE
h//9O8T/d7B9anjtTa+UyRe7jhgDoTHXzSaTgtbuUjKVF7+EuastAeUmaXaf70mAOkfWBTOdVByj
bPz8XF67bTF/9ybXrBbdhEcxUV+UjPI2ZFoweP2ltiBDjIEM1jkCVmZCwFXTu2ehcxK4R1eCnaj/
jpitMDuGEPWnKa29lTtm2C7NLezGjml57Ob6UsncwVfcEsth30fi9SXGOucChzUPIMwk/sELHWqe
4EQLhIQYDPhKBeVKIc8PCuQiqUbTwXX4WWwlALlUWad6fwBTvqR4QIwgGZ0pMqSIN3pqjPVODrcS
8/PfDCmw8MUK3mOhxyEy2xuJAPDClT8UOvVtfm7Zxw2JLxDQx3wUDuL4t17NN8L/Ww21SpsvpjzD
Xj4V8ELaiFeG2gATP14Xj9HXMmdObPKiw3S10K8oGA+je+eiZNzJd/ZnMx+6c8A653FTWcYjNZJO
sAngxFNjsUbJJxo7ZjGmg6oescgatBcxItOxHLeysdT7XzKsv5rZmRosJY68x8Mb/IIN/YisdFX6
lUPBJVDbIp+fpuvFNq6V0K4f/sd0XFhxm1cjYUFBnbE68roQoaolK3KvZgppxOKRf02FLHwLvqWf
aMy8bEoHDU4Bf/8jOmvI1f7lDC9nq3XA522JWnVb0PmStjdPOFSnl0gytT+vN1hfWZ79O1XpBZFw
kmCA4WqJB0bhr5MTUxRahhzBRw4G5W1FjTdia7ni2dl8rxScLDIhZ7rAPRBFBvZydOEVWC2l79FP
bHYtRy8a9SD+VbesSqWhVN9adH5BVHi2U1Jpw/33qUrrdjOSS1tx/h397kWkC0MOKOqBds/Z+1N5
GHM80ywWyyXkCIXxQC4c9FhlFzWNKnsOHCU9XzYNSYP/JsWFZhyp/LYS2ydRgnIUPYENN48MlsUb
OxL7NkTAJGFt/KCLKjLN1gjFOw5fgwmYYxybuJRKq9OcETsL3SgjXSsUS0xFF2dw4e7z1ESm+3pv
lgXnH/3/o/MTP4rzRlAEq1yspglb91hfJGvs/69sx0yenbcnISMruJrC0muaXjfhG51DOARRbRGd
dIcwz5MXwpXx1FapFRvm2Kv1W3qQlie3ZI/2dBxKrrAFGhGENmsDlufuSH/xM7fYQcwlAsPqqLTN
7EwlF9GDICH5TAmTbGpDT8sRUG2OW+eZTTT+iPjSVQvDXmSvB9he0s7LN2zosrjmGupjGhzkY0vO
2R0NsHb+X055WjI9FTFhYZlckRna2UxADjTgkCVK0++VnrAV6mErVhaOzTgUEvra0lA/00YgDTL/
8JmQffNxOXhtx9p5eQ5zifT3Sdv9YthJEBuhYYZlct1QMkJ6dbO/sSF+mqwi3G6K9QN8kEgLL002
FB3DXnKx+tN5u2XgEvTiybovI1blKUniFb+XhzxiLq1+FH34ZUMdHjX9tr9+2dAIAb+e2QL5QzBC
UVn1QgXiNMOycfHwPZueqTWUb6fJiN2s7sPKTcYMwHnNRVX28Xhb5ePTmx2lccsm4kj/4Nr31LSH
BVx9WBadTGrpywcNZBOBk4DEi521yhb1Y32BuT6UJfETLwzta5Z1xZGdDXiXXT47Yft6ds6oQ/R4
kAfQHt6lARt7uvcBsl2bZVYqnK08F7HhPuqrJJt0rWMmFeZPcEgyK9ALSkuZ+/IR08OorXOoBKUD
srsP6WFtDPyAw5tvucNwKKUCvWgK2j87XeM+NGa+MGwdvNP+hT3hp0UOW7pHlAT8PO0eIttgwR1/
Z47zB23Ys5dl6pDzG6dI5fyF4y850hFa4agngcXpFtUbVIi/Pl7cxVcc8IATHQQIgbBfGG3Tbu/d
hpeA2LIHeJ98bH1bW/XCoFryuaB/lvfAmL4SBjVTgDedbuuYaL6F7OZ+BqDhxu96VsBN8i43CKEJ
A/Abhdn0VjS+7IoSiXP1619WhEqTEeTrRriHtUOyFErrzWHhAD4UDsOzrfh9gW1ZoFZY68/bujq7
Svu6qCylyKsaim10/fOoHU9yUZly0A8f9WnnCwx28Gxj60XmdNxRFsD/ZPsnV69+V0kpYu6c+SP9
0pBR4z2/hJh4OTSg1AW7yBtoovtBDi/VsLM5StL5nHuo5D7zM75xD2U6cP32TSPQF9LZlf3SupQK
uJ37ONyw0Uoy+wj8JCjdkS5jayBzfqIyjGcI9NaHV5aipl+scwcO9kC8Vn5x2Z8hC/ByjesfI4uW
8vtDenw7iZujDPP5r2q7bSMH5y5mCKzc9/8HGO0tJjkCOf+hHYiEtq7s2fa+BgLL+6CkNXJNvLcy
TrKGOjTKduZnhrtOW5XnNm2SLrx8zxMv67UxNIQw0HRv7CZ2n0dWA0VOXtVKgCXiEFfDzYhROOd+
2mIqz9C4BY6de4D4SPRBQKGRQF69sZfw8HdsukKdABvupleTuGyrXkK4qM3guLvhrdbFosafGZaw
h7Z86QpWrsc2jlLysJKXDfMcItdUPccy1xBIpDN5pseJaFIIyImUoCEOybbob1/i19ttGVPFdNbX
HcKYar5rIjAXz2jfoItOQo3LndsW7hK+jh5LR6khDdj60ZmSdwVtAPwT3/WLu9qb1h0i98zJIpdW
SdthbYeub3qf3pYk1vhvGviWhgg95OVne1LEokdluWjPKc1Dcb0rWxoKs5nJ1XOEb9z3zQONWdpe
iTNdtn9nCC9NmRJIkGJ5iLcccv8j5dpXsmDqisk9ym/3pPXdXOsVlrA4rcjeP4VWcTUb5NRRPMuQ
e0+G6NzriuNDg2zJKKecCtA6jvT9ZY5ZVBfHNA4D9ExKsRogwIC1/I0jS9ertZBqP29QcfB6fLtL
ykMeGJUYXqf46pK0SXJrsrvkOnc9VMLQ5zsuh/qD0B+H4W9dB93pjiaRkhOWmM7CIhhao+nHm6uy
N+GWKEZY+2ZMu9k65lmZ3zaPL+ikD5z5ykZE36zOpbuvEGc4Ld6Z4Z9yx/IedopUsrcwCxg1N+OD
GczEDTKUCVaiq08U/h3EhS2WApi9c0zmlXsouA7+9wHFYooiuzmU4js/6xPqQgEbhOLeVWr4PusB
Fupied1jRpFcLyRlQAp9T2iWqB+YJ3Ndbg54UPkykf83DHyQw7kEFNZk4s3yfmzNfmHdDSb84EoE
OPJyW+NAf+vhPfh0dD+QTRTsugOrI4Q8gavtLxI6XnCB0oYIGR8IgpDjcmlcOSWGfIZ4EIfL9fe7
iUYpp2guR3cLGSQrCohUUYn7XYohgXP8TCI9I6ofrMMb2YpxyGMkrVm6RbZXcf1EWlDoSvkMvDSq
5SYuxN0a/au3vjx9BfeidMlFym7blHWPsuWV+WAcWm8SX7CipCXJWn1bP/pRsTyxh2T2wigETVzN
kBk+ghzL3KmNJ3X6Udmv1k9QUs1MFTmdfAJFPn4FhIquuDerTcjVMMmbuFThrpyn7cvQdAQedB5P
KjTJA+ijqHo1H3EPUWdatcAAUDscktEjRQNb4kopnM3dlMtB+UrxFBo3VNDvXlP9ybUKRUp4TEXd
VS+0dB8mjfmsyVU2HyuvEKD8mXdsMZX8RSc4bgkAcyJHNoUydUhUwGI3ipeIAyoEJKRzGj+ph0mj
ZnvD7n/+jRyQJUOhi6lfBjKzLTb3LwIEuKpHrv/SaWpi/DwCyydFlq4ntb2lFL+Qsqx/32WJzWo5
IB/IJ64XnDMRlBHFKTmM7CnyuXY0ba5AkFLjODRzyV1q+8LKNF/m331SYkyaRgsemAQ7cI9hHvRb
GPqPk+nJmdMhAkJywtclImmWUdBXWvWrp3FxMZPmq81lmq4zLg6VD84Ia/LspdypOZlwWtWcqB6u
1ZIUFvyoL607jL/c1q9J3AS/GcJC5QS23HFTqIFkha8iCR/q+l19EpEdt3fkO1DOHcqtsP/bY/Aa
uKVcQ/tgYEAzT+KNUya1RL4eOCC2HuBTYOgxfUWpRXUCWYJLo1rEFF+is1ABmpoy9pHz5NDaUrIl
lsxI23oRTHunXZQRtrq33KdLcSZwu2WgJ0Um5/7yUOpPtoTmKZO/v5dCpBUybH/6U65d1MCn/VTt
+zsVarjJlCAlmDU1iKPnemSgBu1R5zIP8oPyLlfmF0XFflOAoVqU2Kuc6ZcrHKhF2r9/zF+TlSTT
EM6KEy4tjgEqTAvBQGcFmKSUrp+es3ASfrRZYiqvGnycUVDnUaaLY8CHf+GCr6cKAkmiRpmkD3Ik
cKGcf+xTCo0fIRVcQ8uSrsBPDh2wHqQUK2Y652JR7/FQUCsaRXdVA5bwipOSi+kq6GkEbtd6HS7w
YFdZk751+w7DGuO+cQQiKzBLibCC6IrNQw6NlYkgd0U7U0vFOlbFHjLsmuRKtCOUkUARjwmotD85
lteCwhiktrRF65oNwQlx1V40aa5V6+hrApDfII1piTEr+czbqy8cxAvtLmJc+PWp2H5DeH8T+bhl
HilD7DLW8JJCePJxIzLmyMPk9TqPVtau8QEL6iK1FhkQJrm4WJr+Kn5KE3801oByS1UpNw8wNJtl
1r3lyclRY/xGqLG9uXZstHVzS4+LjnBOtPbYK1QVXJjtbjvVopGu10y9BPAO2f5lFRT2jSIqq3+M
vUaEx/p3dzM4E+ooS8aWFzQpdNBe1ngxtUA1diOTqRprp8ZaEHFI/OJLzuoSI6aVOnBDXZA3W07N
IelKRqvrWI+APsagygUPiYe3GGvVSkFMNdTY1KM9AvZz8hjNj7+1bXVrkR2fKvPj/+9Gu/BKsC5W
YECZB+BvYEtSOACISjbaZHrntqecCLYGmmtxTS0ykqUGJUNfxht+JxZkrsjAoRwOuLeXB08sjtqe
IweXRaG5EHJCCYJfdcteSDOrg4+vVa9O0guKHfCdjcARK75KTvnirESSVq3PlFAQNWYa+8f5wGUs
AwGi54MMvtczLQhVQaIRb9adWGg96DjraaFbC5rraeRjni/N2Ab0jD5ljx/OYclGsXBo0l/OoIQZ
a/ZEC6AZpogRN/NyAYydKnEE9K83KWwEaKosx08FVWcXRvoCewjIHPbOoUQiKMZSUAsGZVn2Z1sK
B8zgSZ67EQlAAl36EvUWFlB0cO5j/JGk36uxUAeUKI2X9Z1nAbXkDM+rDSzEBCRUOmqzKiqqYTUL
HOq3nL104uN3CFQU5DBnVUvMu5Xvnj4x8Qqi/R3UUbTqUmDNaWL7mY23bw4OUPLlbPHcciCAX0NZ
r4tCRHmmyooDwq6DdVMpUGNLREGg3hGj4owm2zC2Lj0R97CICplsEVeI4kjCHJV6Q2zRhUBvrTcB
C4tFs5txRpawccYd5BvVJd8zZ9vIPiirkkgFcWd4emf8lEI+YllKgtL4PUPl/FuaEZ2Myecp6S7C
+is+n8K7FvaI796VpTkcL0SrawE6HvZRKHS5fGDrxEDhNSbzZ6WyzFHXTy/eljG5JzGAMB1HfXQw
XVPUOIu/+pfJkAJgp+HGI6cWp5Zb8b746XBwIu6Qi9mSwkafbuzWA8/Uz7qz0aM/j5sVXPPe4NN1
2yiBO+JWZ5aEmZzQnuv03gEgKJheL48WYI3YFavKoZV5OEIhSYBSj1WUbIRmPCVgKCRweyjVUSUD
uHurT5/p1zERRVys+Wfz+HM3Wo3G7+VLz9CX5KcqVVEoabQ+0CuUmSIKYSBPqndqi7XRgJeLpCYS
bH6hm8fWzsOxysakNXW6yW63PrNEPCGTGCpBgYWeRca6YEMkwCAmkfWeHwYVZn1yShVfH4qquy85
oA5HQ6CBLvWbm/QFQrR4MLPIKlLY44lOw0yULxMRFcc/Zt03YbAbP0FB2XEOaurH+qiJZ6mWwD8j
WTBVtKDtrhpUIX91VQ/7AAam+/btdT4PGx+3RdU9DpRSXJmKdVZe0/qgYA+b2Qz4LhTT2QHhKMHf
uYXKatpnENJ73uxNL//jssp8BFZkYKAqDm/RVkcP3WBw4T6Qw8fwKPKq1hX+mW66sF5FOrW2Xum3
opYgInnIcJtj4V0VAwm/IEbXAIh6/M8vh0Sglrz5an0h5SqfQ+b1SEc8dHgylsauXaZGJkoy5efm
0cunX2Ntb3lzbm1TGua96XeNUeVwhQC/WQyhJtPoadfbjWH1UQZjveqLhTjdgyGMqt0KATjT+JbP
9Z4VTGSSYsr1QAo4+WqfH4r0ZDB3nrkk5/wXUnVwujzI3/rg0UeGlQVNAQoT9JxrGPqBJNpfC2S+
VAu0C9uL7atqvInsg5dKKEWBBaejn95KQemVRYmoDf611oHMMaqBtGS1VWbHexSOba02J9h7ndDu
qMelouFGc3Xj60jOjyz32jFGWIhOyNBozi4mZK7SPBL4PTypTqqdsKjnMttEMnXXbqU4lZ+oVPoX
JVllbbAAhvMvpXkxWkXENGFVKdX5TlEFyaJgVhQgPo+x1siUBSoIHRsTSSlmDOcioxadV0bBKUkn
lGvkVz3ALm6JW75+WFBbFYCzZqo7Lmh0WtEaherUWgkxyRg8RQbM/3j4qDB7dQSxyWjaD2XbPcDb
SqBxbj1hy/qdnYBr+ov922t7v/73poIyjj8w3i2/iKky1khMDz9qs6GToSxmlBrlVIVFieQIKmcX
pQDgs+F52lDyhmadTQHBYYHtRY6VaWUWEPzLfhg+jsDvIClMVnhggb4QUMs3OKyWEc1vFFYY4++e
Sy+oc/OmjiVFbiR3YD7Hi1Ep+v6gJO0rt1mAcfX6qCMPaDw/xOHQEVP1fzx6U0Kk2uCE/3qaRdND
aR2331/0LAFEZh0tqJ3O4ks+KvgGrga9VJdJom/6ToUQ/ywnoMb8itoe5+jgBhqAHBGNp9MA0Xe5
p5liYiavrt8VA75Uwa8eYpDVk7VTPon4WAiRPX1yrE/rDzRHMVU7jqTBASSxNwh/h+6WlLF8rpda
CQKzGTVpsrXvARYOVeyRfEN63AJiVJlfl92pqb/NkjKzSIA/qqkMZddWl40MvwY52ovRruIPybGb
GsS6cXE+m6M8Ouu9QgecVpdNFS6ZbzGscl9UnzP4GcUGvMkETl55CqxIsH0+An7cRIMUv6l3wgmG
b7FOVAbk1qFgsmCl7vXY8RQwWPwQsPiGsFZF8IN+oP/dJffeOA/AlYaZbjW+iwc4hZlEqSOhHpIz
xU0wQrHU5auBqJ0e9YH/+9VvMKfcKBRjMVGGd8QN/VgqI2tEaM9wdWDj3Q5LQeAwKzREzFkDCTM7
CLgBbETT9q387HwXrzwEYWIhbaCxRDyXr/kZ06KJ2wi9qWnR9PRksvU50E/dIX/c1RPeLz8qyRDw
/0EftqViexrXx595+MRjrTw8eMzdVIh0ZIjOnXXMoLLycDl2kjaCnu0eNP5+ggkHPTTmox3TbWoT
u2n+UTeSC5h2dOK/3yHNJPhmbfNaYGQvHklL+GuBLBcBIwTeN8IVAVWSdd+IMIwr7aO6AmvPo8am
QcigfNdFZsiJu2qKtfsYvcAd8g/SOAsa4HoGIuk3RG6xP6XokB4h0JRrqW/RE2cr6KSxnQ8/J+6x
wPqz77T0csRoN6QReXnBeiqTIw2ytqhRLjyEbnllgdevrD1xf24jLAM++t/a30gdn4WB0vLsMKiF
g0gPaV+f5/QUuIoAmxdMv1Bgwwmy0XWDIJEPHe4WI32HtybUsmZAF0bTeUF2qIAd3sHhD0g8nkOI
aIQNltc4cfl5qrvVvAM9JGdPWaLC37NfnxvjiloQs9zVG6LjGQCaQc7s6KvYlnKPgYYNPpJHwDfU
MX869SXan5kAeAR92kCegqHM7jIxFP9U8so/AAVmUED8bdBAnkVqmB/RhTZAJBKxSAPEpfvLuKY7
L/WyFjdt/rzXsyl2RIi9wmANHZtlhSzgyci+CvpocHRwHb85V495BsEuITnbdXxqA0JISjuugu7P
vOK2ElZeLmJRg+vq0kIBr8w1rzopw2Vl5gxwsOhy1npy4xkYozpOKgNIAUsNm84WjlrnegHzktvw
HU6VkZ9RuJMqXMsT7ANxfxptDIITNky9F0j9FIYFEmK+GnkTfIi4DLW0Q2xknn8Mc+zECD58/4SP
J19jhiEvQi6NwucmeRJw3/20FgLZfXwNg2y/CTf2WNLN6vFUof/NETHXgksQh55GYVMazcBsMkWV
pEWrJ2KFNOjiX/CI+G7fRZOX0XBKCOIoU2lCQ06M6YDI8sifbLYt9mDU6iTtwuKBAbRIDowT8W/Y
qi2BjwGQzm504dufNqOCMDRhIICxsrvmEEXcAXIEXkmNHnl63SpFuBTDLhrGVT7Zcj13QUflRtMp
i92QYlIdgImpA3Qytj68GmlMfMyNlN1ZIu6gHb6SOR2o+Q8eZuOs3eh49vdmXtSuFWcQOX09SzT+
jD9QAoPUDmIDgpeOrEarl60wpayB33ehYvWfBgt3TGlW1b21tKFbGSdNvi5OEPtMs7Fn7fwD4d2N
gfYTMZVoHHhoPCAlfBQcxsQDLC1qj9aMWw/EroSofUTq2orxo+22KFG71WuJlYhG6aV1MxCcS1Oj
gC2u+M+froVfirkadEjJcFBxDu5Qd2RmQ1OZIpSc2toccx7shtzlPJ4XdaExPMWwmBt9nyi+BKTa
+RjjbNHqAe/DRoYsFSBcK57OBwuNp+RjJ8bh+It9SarBEDBCkxUZSCk223rkdBUf5KB/v9cQ94W6
kmMASWeDzAPL9U1DPGcUjo9ItbiOkyY65oBP0z+lSZLjsQ98J17gLQ//lH1KYHqq1Tj09gTQLWdl
dFGihQIMOpj8YK2R29Dws6OQOSt1fNnOxYS6L/svqMsApTPo7NctSNRfQFpSZbT5kv9gE6WTgxUb
kRlKPxjDCShh5oQfWBtRJS2shxIUC6BgQhIVp1wZo9B+3G42YNOp/869OW/18+fCUkWnR86DNuFZ
VfTQNclrGoUaaqsW5rAXvNzBF6aWIcIa9opsAHEKqSG/fMd/9+6UQ/uuKCwVJHDlmsiF8uqOrTqv
uemB5g0D4FDklBuh/GZuZXpOCZoogmkBm6pdHXBncvQcWCN8lR1MKG4dsjSLmAH8chbLfDnGWX7L
dpsDW7m+oOINwiT4DZJMmDVrXVtJAbgLnIBNVgUMdDe02ibaoWh/wFjZteHbJ5uy/kwXHfKgtpcW
YdPE9WJMVQEqHU+cqR2wqq5oaPD6hKBh1iSNqOl8zQ+bwgBX3vJg9Uv/04RQvAFk3yLmx7DDN8Fy
6vivN3NOWxr45CVLux8uqlATCS3OwQhEnbrzAhW/PWd70PRLi2qxRgcsvQoOO0LQYMGCN/4jtYMP
6EPifegfmVusr4tN0WlIw73YmRszyFzcoLVqkeMFeJhnMY5OppnXXlg+k8N7FEKW6JhhFzvFax/4
KYFOlVxhhsOtlRMYRSFLmblfa4OCABLlEaPNeMZDQbfdzJvJXnNQxJzOwKRGEHkI4w/PS1UrpReY
Rlre19ojD6DHLMYkpkeih4EBig4oRX5d4SY7FkIW27203CU89hnltGUqtRE3qjzRpfybiN3VGj+R
8dykyfe1+ZyKjAnDMKWCYzCzl4zceOdfcqEhACt3K4GTGQUvoTN4sjZlkgOlJa2Nntq5hLoNrr4D
E3qL37T4sR2/cVJsjopCl+K5l2pOAVVjjGhWRDcT82ggYhEVLkCX1G0JPs75AzKk/WrZ8qtQEqFZ
3dkKniiUuLoIARVR7KjkMkm7D+d7oJZr4ZquhZGSZckaYQlYg8XF/oV2jem+O6zEwRrUf8pQOJ1F
+NS3U+q3FuAELuRLM4davK4tMwQqDgyE9oA5/pNekHd+ldrHkjYKfvPePYo2GBx0H2Qe0NZHPdUq
fdJ+zKAfVTzg2cHAazcuHezq7QJRqa1QoT/LrZYrT8PISdC3usJiLdc/fB7gkkQ9Y6xvDsgRgFKI
88DC7QzmM//YbvYCQwEOIapjG6CkDHPhpFMPWhSIzJ0ecCTEsuhjoi8AdRSeCMWLhibxWyx+esHq
gEpVy8ILtVh4dD6WL5520LnEmzOSCJ4nbtPxlQ4G4cklYeUlqTgTvi9j7zP6gmc4mYB7K0OvFbRJ
esSxCliPtuLeQ1x9wbyaZMBvkK+yrtEBf+brq5pqO+8Qff5oF9pGac4N5Tew3DHs9vZvlYWeUajK
eusWRRpTr4wjH+WvyorprPXdmomyYnK4KeEK00A2G8n2vpLEEdzzRJt0J4BwNXg5JVRKAZbFylnV
qg24agbIXF/gszIC3UK2UzjPkawnMmGVsSiNMuSMd7zTBHCaIJr6/f6grzT52VUvYHIUxyRDbgOd
gOFp16PmXVsWEhbgZsCotm8PkQv1WgsHlPkTCxKQ9n0Cm+zfKkccSNnUT4pXWn0FvUHq0VgnBvoX
RGHBJWgXtFpYm73OA+H8I82g5NtJe7JDqhapMiE9Bsx3V6ISlJestl20vMjSQSxL3L44WjPQHzgy
F0PzPmuTit3EPv3WodQyibOFfL4BNWlw3nwDrGWv4nqxttoZ5dAdxZt49HPOV+t/ln+fME31tP9M
+nqLbtj5uJ7mzJFm/LZOeffjmAk1163ZeL1x7l6JMJX0u1eNEpdi9P0Q6F8c3UToaQT/q+6TrG4k
OTtWAkhNAM5DgIwwxkf75f7Ngsl0uQgNah0N/kafmntjyjVfkf4AQjXAfpJLqz/6hhQRjxuAeSVA
DivbCWak+xYIW1dF1ZijvvnCcI2XfxZpxxXHq9avDKY+dKFJ3LWL2o/+XzWv9DhjO468Kyr1/I1w
cIZDUaGTztg8zhxpoz0MJzsTvnxWo4i+7SjsFUYFhVIFDojEM+59AqMvMbU/SqXP44YZiS3TAwYw
mBgsEafOc+920A4wB6EfN6uSCzTLlGmpqdXDIyI+2N4Q58+qjOMAMf3k2uoHnPGx5Y7l3WRmbs2e
RlMA1s856+KpGp9HiiCLhbZIIC2+dC9DfTg5VmEA4EdOGQxFRDwGmCc4TEukape+VjTOnyXtcSpU
8+otLCZ1/TfF0+znfxrpgFum+Ozv9eEd2Mo2q0AB5E1ccCJjTIqvb+ym3/x+dwqzjnaeotPBtFH4
KjHogc+Q1sBUVqAtz/VRYz2ApXKxrRbP9QzGImLkaO/+LCspckmspMKA+YgBLxuVluez0C5i8SiM
PcQn+nJBcaNqeioCPPU1DtcupgWdP7fmD3LnBvO/Sae96CsJdpiB9KGYPVIpYEl2ShndNfnTOve+
OV1VzU6oXI14CeKF/cXsLQsQ1+X5D5ymeBzK04ThSFNrlXFDHDyyqOtqlwvPSZe097hRT2jEjRW8
SHaDdLBxrU4ubsPthy0MUv6yRGFXsmvp3GAFxPtsWveYFuDJ3lbLxwf4HcTQdnfBQaltdWg9eWHn
NnzL7dGUjuKL2np2u3hbnvAUKQNZQPOAmGBqXQbs+9kC0ztkYj8u0EyWCn2fOSRYHeVB9KiEvc3G
d5qj/Hle5blll/AGRiKCz+p37IpcLdZb9qPlfP3i+kJCZmeHWFLDSUnPj4NpviuYVFLZNrf9CRFe
sR33aQrJRRVn0ZM/jyw672ugdD9dxUqAI1oyLcOC+GwhLVEAzrE4MJD5Wy5FDN/W1rdtl5afphQX
cap5QAV/RYu3IDPwcd0VmKGxKLDH92+EZtoJZBlPfZP/KnJYyY9yu+VGz1tFk8ibD2J1mLGApmSx
NVAUOcVxd+VlCFznnkWn8qKLELbkX1wizM14mWWB2Uk/ROhiDK0pK9qqgon4v44jSbRx1VhfQZCZ
vuhW+scWdgTtFjHBa/vdY+CbvvTNw70WC0pIplunhqy1ze1jjohtRiJ/IsLAE0o9Qf9fUcj/dLN+
ZlYU7oJvz1GuwtLOX0AFzzZKx1/dQX/r1+W3tSr7Wre7Hpl9G8k8mBzDhZAk/k0cYiZytCnsUkeV
N8Myi3imPw8EiwAHgn4EUXmFe5WxnKE/H77v3OeBP+T6eekktaC9+0tDrqBmnMAlIvbJzlp/3gfb
6KTI5mXLqsPCcX8FIHiOptdHoUsOm6HNNiActyo+FemJIUW/Ug5+096xl+59Ib/v0I++ncSNjSfR
IsgvDk6nJx2YDtXaLTRZxglMEo7zwMKXPmzgxKlqMzoye6tMXbNxW4qroBTwsbH6QHDI7Az4RMJ/
zRX8cyo6gOWj/FVjHWSlc8JzeVKM3THPfsoiAKBGHZ7iiIwNm7nn8RixFzOD8SQTYsI3oaXTdrsN
MoDRu0/VshYyUoH4EyEl/gU+nMc9wU7X/jRu/Z5X6RLgtoZnJsk2Gc6BpCNXXAsKsIbtYmj/WWlI
2/2LqExuMQldLvW8PKBh/vlJIH2mvU5mguT98WAz/ch7lXDaxqSIscabV7D4eTt3aosAm0xZpBxo
kEMJnXaiRMeij07GCaxtUaYbQrsh355WfiL1LFYaKCn2aT27eo8E4RnlQbUJSVtUnSVYnht/zuk0
SZJIMpF7/a7lKhjcUWkMPBtRt2KnnrTw9VcZUT1XAWojG6FkjQgG+tW00dnWcPK//cALQ8toVWhD
9iPL0fRXmIKM7FBvk6i8r+iTf4CMLeRk7FC590dmSn7kb+qXTyXkw5sGdiGMdHqFJnx7tGJF6PsC
MjZh5bYpcWAMMlf0g6Q03eccguKlYSz+xkumpNSvAXdzRLJ70KTW/XMSG9Fr1laXjbIHRmmmFqiz
8sRx80p6vqFXUnRTmWsJKx+ucf9aK19v3+GgaYEbNtikzlCxO3YozGl7DMpZnETYCEhBHGOpVmyW
IAc+AErrjhzXLyd+lhS0LAWk5H1cDaZ4OFU4S43/cg6aaBxJjGmHpEUOET8SMcRL/1T05POTFh8z
96ecfj2YT/30Fn2m+CpXOk8tWCdx0OGltpSdJGs4m2lskcSlVbCuP5KxRQX8S9jy8a8rf+/PdSvS
+U5aa3H3/pVBinyGy/NJCzwu+k6QNYlFAAEb/VqYS677sNxdJospFyJodltnfj7701+TnrhqKqFg
7vEJqt8OzkmJA9co6e4ULdeO0Z4/6/P/SPAPUAF1aslOPn/qa5FqhQadODFcHAryOe5Wklx3pxlm
f0JPItklDMw9uiO29OF0CwxWETLdNJRCrbMMAfBzHVf4eY7/0xzyNGVNbcjaa/+b8+20fcq0MEb5
o7izuPZWe+diUiwZoljohVlCEdHIbUDjCw+k1ikp42aZIVyB6P1i4O8jO6t5DF+LaL7mkUrwYGFV
y/MnBqI/CILLQuYYE6+iFDEZ95dkxYHmY/St0oyWFjm1IZxsKau53jeBsbyNo6THCSOmzNz3/6PJ
uB5+GEc1Cx+uErrPUnbhdG8O/lb34kgaLQU0kTcyqUnI05G3XKrJzoHasHbGvhAC79OdbVaKdc2g
C3eBRtuzG3x9a3apKb7wfdj5v5FbLB5ETojtGHs8SLJQ0dvcKIuu/SZkYJvJKXLezwMPydA7dfd1
Vdv3i6y53bwJ9ADWs0wvkcpicnnn8whhaqs1y8wvMELhR4SZ8WD1GZ3084N6G1xUuxe7LYI9BzbL
C+QTDtw8d4/swe+MVUx5axKCOM9J30VpoeFyD40GeQbx/uI5O+Th5XaygBAdNaYehP4jzdyyxXL7
6QYo0bdHYfatp29XDpvZ8e6w8TRUkB61OvJsdma7OKniRWshIrCwnjgO+zBiFvSRoQrctmUX7A+c
U6ubM7JVl65i3q/CKpsojeNI+kHyhpcvqtaGVub69Ekd2EF6l482kbzE2diJLCDZSTd7vmFKV2ly
iTI9v/ZMVgePemVtWr3p21JabvrnTSFjxWPfAMevG6MM3Ceud2hY4P01J9Dg1vhy/w+Rsln9agB+
BAbWit+wfhZKcLXPD6DCA3ey6myiJsvQQEj+b/g5eS++a8lQ6Db9lrzWiHWdPrWGe70/eSDsxCnz
RVbHuV8i5NkUWpDNa7IntjURy2VBET5bz6izratmMO5Igzu/t+dPSdmWqucc5ZU0lLLSv0Xx5uhy
V+lum4AHuyI56kqx6Qm057qhUEDguS63anyiKZSpWhkilRAaQXCsOPsMt7LT/MiOYnkG52d/BgA1
iOpzwDCEoDMHWTduFoaBNN/sJO/gWE0jVnpv7noMoYuhf1yY1YYcQiYhdGGOWadbiV/p5dtfPxC8
H7G3jTtlJ82V8O+rYufXW7SfTAMf4gNz9Zj6heXwG7imzjfnqzuGjB2PABxtGsniCH+RjhE5erNk
U51W8qtxRa9CAw4bU/g81hkf8HjaPqwy92zHX6ZQphbQQguDObtG28tS6QMLYJcsBWbokyHYjNxj
EyvNnooiRfKSattA9EwIUfpddA5+b17ewZYiyDpYtlrDLgk0FywSVXxPzLJo5NwcAWn7XVGwe3F8
3rIguVH9Jg4I8qjREVu3Nueh+g80mRHA+HbHwSWmOsgGH/gxIPxLfw7BCgq5EbrWBbC5+jFzxpmo
EGPXxYJE3U661o4g+AsIa6Mr2ic8S+Y/rH4ISdnvI5vTw6keoXkwmPpFC6Smq39PHHUEZnX09/j/
2w9NPGR5dJ/mQHW6lf7DJwxSnRrQEvsuNtZr4tQ8T+RHoJNoJh6M9Yn7uWALsVSJXJge7BI6gaxu
QQszJrDwpGQMTavPMpnxuWqsmdBGSv/THFw1fPvhih0qndqlIMje25n6lyvyaHP0zyjRFDBnMYLq
dFQt+QBhqSK9NKx8aVYUKZ03YLikUPi5l+DFRc4MhA0ldSY3Uu6aSh3MAULnsLeW8XJbcJbMuill
LU8Rm9rop+7dCJwdum5e92KBW4JA+VyOLqRz6dIEW7wWi95issIvgXeU/GiVPs7KRdBuJZ1jBMSD
4Id9iLLzDThVXeJOJ7W4dyG5wp20xv5QYsSDXE0fjVbS298YDg26uZyYgYE//lcHr7FW0q0hYzX1
lDD1kUX/8va1M6o9ax7XGtg1rpyii2PulDeSbGSr4+PY9tKfZf8dikM+BAU6QXjkmDDawpSkaviR
zNL16utxXC1ajdQG7T+CF+FB/CB+jNwcvBgDgaF2+2n8wScdC+qZSFz1p/tVkpT69mnXN1YKFHkd
/8C0LlMCmIRh4tpYvHPtQu5tw60pM2xYDJ5AOZmsSCtC+R1g7VhMRlAUEnWbl8KquFbmK82hH01S
s3ujDeCrAKZoHGdXoj6Z7bBMLU2cHrDGOSSPYGpl6Pk8nlzqio+q2Oj91zaK/x47XjAGVrcUNYbE
+Qpg9PQcREnvlofjkmJYtotKZvUsNlPlEYGbcvShhpeXU653NGm1+qutXhpLYwGVslPDAc3pbYLM
AsvwptfD5vhBipxk9FMIthCHGlNhiCbJmzVMYXRcoTl1LnnDOaytk3MbS373nVzPuzxmkS+DGlGz
Ozd/O0LZ4Jwy2IPTLfzJs2fja/YifiY8OyZ66VzcPykMlZhClBhvnCVLbRMh/jnm4o9hRFMIlc3o
BOjVwaS0DhJOOj6DuFjfBK8OtdUiwbMqZvdBD9EWhEZdrdSU3VLGBkh5Mxso4XiuxOQXalQSgGE3
5Ng0mTctE1YZ+d0Luzi5SajgUIea1m92Ulaz79MvGeV6nICiahC4JpNNYTexd2s4NzInXeVz/5kt
8N6fmHRo4aD93WjN9W8hipkIo4cr44G6ueoP/iYxrJbgobMxvh9QvSsdYawKqnilLR8xQqZvUUDe
OLq27yFSVobDrbTl5ZUY6WoE0YCMhYqtUkarAeE70epwdxyN+eZEfWGiYWdsZ1claJaB0azTo5I1
t1D/kSlkKBg3uonQi/t+8ZB5M6YwvUtyv1pkJK4EW2YhwmdkPrBdZcYaVb+b+Pavm88KimK3yMAe
cy2ndROez6WgqUoTNpZuto4wbbvMQ6t1eRrpozBYYgGp5+DrjArKGPVPGUh7ZlMl3rLTrPZl/tVB
AI2RNy8awXxUq01/9Gajy1/anvYZSSAcyLgyBXOpKusQGrwLADBGfc1TWppyRyL0EXJR6MRpc23A
9uAWeA3p6T8xCL//kXGHgm1Z8/83pJ19lV62jNThqa+iGZ/GHc9qJPASjkrRxOqszV1oHA3YguJm
HQb978RyVWfPazCFKv0tWPlIVy9VCb25Ip7Zi9OrYZZbaT2IUCg7xAozavxVzDsSuymGOHXtoFrG
EyInUj+kKIrJWrGuK6foYOy3yhm+y6iaAXLc+Y6bf1gHfNQhllxX2z/igNQT5swJtnJf2U4ReaR3
AV25GATGgbg4GcXwLMb7VZV6JHwmKeFRAUQDlOQCIRDsUNHo/tzdT5EiZ8DxY7yU2VYXOEvgB3Xk
dc/3Sub6M+4Adg9zoouLrkBX8GwU2aRZtI+G3HjSJO6WlOLxeLoItITVwDLIZRPZagEUqTz2cEad
NTFFX+zsm0g9Pmzk0nLPS3O97Lq096ALS7rgubJzecrZRY7WuE7sTYBaFHZzBCzcNCcsjIFOky+g
opfySlJlNw4HE8+NF14K+cKmPXDQVJZEfrx1cLtNxjtisEJQrOMlozJ5BBwT+aq76k+7qKwfCAuH
PRnrErvzaS+liqyapunW9FPV3j2gFwy4vb4l+Mst5BTEp3uYVD8d6VJbA29mvYVxNG8BV7tqTavZ
PrPhCg3MkCqXt2FoRhs+EhR+v5j3or7l8kQCrt59c/eDYYFRTk+T7Q0LX9hfhwQTJCFoMGQXUlWo
imPS8fBj1CVhUK3YgcEGzthtRIxLG89PXbW3fdF0VgLIFzyXHsgtwnrhfTfu+sH3KAJYTcEb/UWy
JJsWRn/hRzTiSMFwLp6/WN2zKGuRXKTNGjrMPGy1TFuWuN2xA+xwkNS9cAeqMNeL7n6cyVPA8FaY
f5zMr+Nw7yCqPrQpX2Xz2KSifIAScG7zSOkLeJcMmdGN0KVv7wxF5xk2SX0zfZjqI5l3ydclIPaF
Cone0RHwAXRCvPWlKFn/SKhJK3VOzoUUKI1jxSu/apT1DeHMWcCflJoWeyGBbS2MpFYbXA/fQEYd
qX01MRD8qO3KQHUbpFs//m1xezNuKLAebLtVSceeNFvZ3QV9936r/0YunS/zwl+NgVQtt2uHJ5KM
+8SI2KfRNDfZTIALAES7etwY7nuHoDQkXo/hP1Cb+jZG+fg6/XAkgMWIxkAUfd29DnV6bSeGoQl5
y9G/lzWKkqgzmze4CnpT+rImvdb0k5+7fTojIJvz1cKelAEJI21OeTnk2FT2ZUIuX+bhjIJ4qxi3
Ehc6P1aUMYv1DdJ1B3zAhlqXgMfvMrmIWaK0NExNCzSsKO3/Bi9B+6Lt1wM7Ni05B1k4G17/DK10
jYn5Cge4sXM/viz+XHI0ZNJEhiDIIkKEVke/G4R+uC4Xrsm8xOx1wg+mOzzxanVOUJ/Adho4xQq4
8DmLYjC8FGG4dUC3t6Dheo13+h19IUGNHfK9AMkHidW92kUzRWwZpEGlwYtDJHMRNd9KvfDQpw6d
gZSM5FyCP0mWrV6WLSrpR3pFR9mMFz3SvEvdRLXA7DkXX92doDac7VTaEpN0DfHXkBa/4prjsS1o
tCfYCPW8P0kGfWn2VDlgGeqLNc8V5s2AbNJegoFJQCWsrGiJ2cxd+GBLXC28ERPL7HjDajYy/0Qi
j+aI1Hb0g9fLjSEJVHlVlf5VrDlRkP2KPGSxdGMYHoRDYntqMUqE61NSj60I6b/mksE5mxJXpizw
ZRIORz05SwlI/erl5gof5ItWBzwWyZOYIps5c8DAa5yqnKJ/cW4qaclVYg3dyPEp/FtL2L6ZG011
ZofLopXh7BlLKiq2USY7PfujB+SJQLt6F7sZy3wmpQIPBxMa5pDA3x6q20jjKB/ekqCAnSxtsyPd
+I9BIxjjNPtTEM6hR/LTUYpgoYTMFOB6HuIT443ALXyk8PMYV7Rl5IWvuYreAfad8DMyV4c3aDLd
yhV9wWV6yHiaMbSVglKM8UNQRHjsFWdxa2lDX3WoH/M6yf/aGRoQMyizuWH5iyO09k8M5fQco5Ox
sgZQdVCzqGWevHgRVgRXhWgnTAs9Ldret62m6nxVPCC08s8oe7/8hfnt1mbGW9Y7VaNZjPz1OIaD
33dHoiej8BaS/VPWwZJyI8ZF5VUoSw1b+TnKmkDhHOSs36kGF31Y63w2Cvm6oM9QUyp6sNfhIeBm
1x2FbY9RqEiWY55Bj2MJ3tY2DMuZfssWxtIroiXvSvcrGJhN9Nr3sYy0+IpxEqjxcBOmFgi1oQrN
p3cfyj1zny1ZI793Du4TJ6jVpWitUzpzweufXpUwvXlKnf8zWd5QeFQMI3tKO0HOBwtsUFwatnQ8
Ti3RyhHACJ3j/8y4tiKSgRKrbzUJl8QGY68CH0ePo5YLpuQIKFjnbvviL1AKd5yJT2sDSl6YJl2Z
Ys34/69grpHfZbuo5Fqj7+c4IWR3EKxB7Jc9du99OTi5HgY8oUQkHmckitfxyZXzgJwOQ8BVZ1Yz
qokoAJzI+CSRb+SNwfAFb5kDW7RycBeFMUWirK4OktP79XYIv6Hd44b8+gZsQzL5DVLLy5YmXa0q
O5aZcNS5hLmS/MO62mDLJC8Zezw4+opoCzYx5D+1xc7fvT0NcUdO0V/BsJZ9wnvJri/jJil5Rif/
+9BMOLP4Sy6+zdd7dahpBQ328jbBOHq2fIKyhcag0MOvnUdWkCtB5Ke+6cVQ0U1CyRTFRkhS5r8+
QNP3mDFMVOeO4Q4UUkUYzJRQm6cHt0b2Qhmnp5Xuezpmu5p511PWWLZgUCB7LJTx3n/PWfbSeOjI
8AGpu3kFSU3bYvmUgvmwBtQxCoPCrxFKzCKeLdEIEwN9p5Ix5NFbqgxZ44XaO0Hyq0foxoKUwQdt
chsADIZLrRBGNFig81rsrHaevWy3XuumaLiuKHn4hFY7UIjttoaLsZC7oLjXMNuHtDPfvzBjZUqV
2Go+kbqM6QtVwa4bAPVQ4uJL2ytrqCger9ZUDO+Xzx7HAwJ3qOKJ6oXvINPQI4T0kWTixyL7UGwq
FTvm0GUGZYpfG5wGRBa8RDCilvispsozGxpP0RmC2XqGw1/xTHF3Sg/2m7t3RgEhhFzOYcNjjUqP
VsQnYWtIdiDmDOCENGSA62UlbTcP/74X/0RqllBH6RAKISk60ftO3vkAkwP4hbh0gREyZKfg8a35
KO9QcR7aA791A2ogO+Cka2x+H0Idn0gWbmEV4xnKKSgD8hCOco7agyA4k/fZRyvelhMVscf5/3u0
sIdTe8UvJhz3p2mUUzsH9hAZEOhlFtfTWjUue8sFt4pDxC1uL/Jlzy49W9Q07X7uJxkFfwEsi2F2
9xXwYTyACweLV55t4MKfmgMlumb1g3kSYoHj4R3cY6wJ+mUlzU3+me5f/FDHB3zQGWB665u86Dw1
Qbu8drh68hvRb0FiJM4m2VOLurnhPPhyhuuhHF9wMuPYSEycIV47Fr/zgr9kXD1oP12HirVgWidM
K2VTxMwGcI/NcZaCYwggSRDmdIIr4IArgPIcbUo11+ByrJeDq6OP4kG0tMEOkAYT7gu6fNfjAuUC
wzXjXvKABld3GBEFdfaReOZNwJ3+ZpVdLu7wRqv6BSVbiew24CbPZqy7fXqbdpDQY9L693y5Xfau
UZDYYshGYyvXcm0OMWWjyE5zGnB77Ea+/kEJCnVY3OLDYAD1wtN+h2DVQfI3taixC0efQEQQC66I
1ffVjDOjG3xkiOaOoL4FniuzwiEyezXSuBP9nigBVfuzyBlkhH79QERP3X/5DzPtUKSjbHcPIWdG
bQfnSrXNCKBTl5PaRjGyQ8ma1wydLAdknpEF4DdhijqgxMLTos2ZexIornA9VDTUnd6YbS9bi8Wu
V+KNDcG/u8FegQqNi2mKruT8lwc1znZoQcY14POYu2clfbNrxYBKX7pm5DG92QULBzahbyqg9GSZ
ZoimPoqjOpBhr0G4Q5ZYpK2YO7HoFm75u0yVdWliW72zT6B6bCvWxLZckX90i0c8cxOUvf4f7Vcg
uEufBfmjgjFpCJGHwU2JvYWcvuTIUTJGxCPRu80swwL7nXCHLkJlk5kTubCa1Ffe5fkdSyHWMgSB
ybC/k/MBi7lMy/FxqYU3rsnpdVt6FI6EdU0vo30pQC7fT8f4ATIikLoOLtSijJRZUbRFyYu6gNB3
Y2Fq23L3NgMyB6s9G76rJEB4E57PhrNTZbf74hpG9kn/LzTuWZbMSfGBY1wDGzsobukXR5/l3qVS
QlOWg0Fg8GhQru9NB4aBCQFi/RU5utEY+LVmAQBTS5hqHc1VmqW/GlhwwLo5f13Q+KppdOgcYzTR
A187X424J4Se7sFuhUqW/OAy3g0FKfq89HQF6tp5XYkkzCmLo7J5L505Qrhoj6271/5J6tkafkKz
SOjVKMOEMcrBRA3WeQJyue87MqSpGYedUT5jEKMlSlrFUDvmW1/F2sAYbBvkhYJNj0quAWSrj95n
zbiMEYnWA0EQGnsMbWH0ytzH8AMW+EHppiCJSsGDXHwqhnC3wZz25CGNngPmYKX3akw1zW412r2l
7cnFE8agmiT0AxvfbKaQJE7f4akl5nqXPoFCPH/w2WdTcY5wrE/R2iInDzxKsqA58fd4qRRfNvdw
OHZC8BNsavKkki96VEULcMI47q8ex6+afo3MYCJcSg0wAl+5BTbWMTDshlUf30TTDDOes2jtp2w2
5DLK4ambiAwO7Nk6+laTMXYmNLg7Ie6BkFlF56RmQPpBbhuAe3PnhRbgxzQu84OhgK2KeyepiSg5
YsATTejdBMlQWzP6/BqY5ecqqrc3MKj03j7x6GfEtJn0stx4s7lsTeh3/HvexmzJhO57TeF1aBxR
GOkxmlPFJKZNgSJe2QbGc8Ihcw2tdtqlny/jQr3Qwg/wBvXeN8n1wK+vsIF+ZuuF0lbv1urE89hu
csJkt85yfvgFdUYGGpsCbYaP8RcLmv3Mx8NhvuvUYdrYnDCEYb1WtzanvTsA60GVE+TE6QALN4C+
3Sp4b+H869b1zjHCGQJHTNvB9QMAfJsEl0w5ePMC1nCs8P3qZ+T04leq2Jfb/AVOMFKNV4Y26Ynk
2cUXokOhU6KCEyKaQQ+vRwxNW42dwc74CvP4EIcZ2B16eGYOzsdCuJgZS81lrULMuJ6Xr89c2UZZ
ppqNxv5ocqQfvr6C3bVgfqXk5t08P/7ZX1SvfhKrXCVws59vlTfFAKlwJr3z0Le/Bd6Gjq0oNeH6
Jq5vVuHthcs7zPxQANdYSjMf9DpF4Lg3281BPZhyPiKDtXBmqAAR2RjzhHiSeDSVtMKeRjgnkYd7
YclTKxl/9TRk22DnDr78wn4g+8tGOuC0wiYOc/zYwBo7AB6U+32hHF3FoN8RsSTi8Wb4e9jQC/yY
ratyBbCh/LyXiqKKuoqOT5gHpT/byv1iTo2/gnIHUM7KqPJzxmbTBjqaYYJ6A5d5m/u54GUGEh7P
WmKTUG83F5iHe9CjsLRNtKjS0UvNAESCs/W42O0XwEwoyD7xblTsKkiSQrak/U1z+HIhCxgOsIiX
q5h39tcvZpXO95/GaAxFVYNNgLkennW1n7B1ZJvrt/7ErWARUbHxSoZ5fm8BZkExhV1fyvcz5awm
T5M1gNYqBK/urjmph62nGrpvGTi5JuhLIqwuFSj9OgQVoB4aLIDxa9CpCmTPK+DRa8mseCCcEteE
SJgOMwaD/AYkzokpPXERQ0lFS3bRxX6aOaOBhlbKtjyGjTG8j6BJWAEjymV2Jp3WQkY+4hbPcHWj
oNlBhmLPBNGpTXKFxb1Ym0ZnmYjPY6qJ/H8Pnp3vH5r0cguPAcfA4lAIY2JrCYZb6qNRNXdLPwgJ
q2fJc5Jq06sYmfhIXMUqxGING1ISAF8tcD9yK0l85prvwxBnnMj1pECxRoeO+BR//GeUen52zrOX
LFUQj87qqp+Qrx4PinKZp+OFVQuJWZdV7m94KFdrcjNyqAs5Di6WJ5UqrdzmPtALaXs9zyrGmLvG
KKfToGUvgdtYbUjzdnzvgv+CP4mbN/WuxbFuw1YmxHKAtP1SGgJXnIiCx9VFs1IUM/tFk0c0lQnb
SkXJp9OMh+I15wg8iwC88FuwEz1Qk+1C58GrF02iv/PjW894zh5HwSC4NVSFKuQjgh+cUW0C73aa
OAq8QG6ZEHfEwV5rOSR+TLTkPIUj1Q3+URanGLMO8fJPInL8XE7J+m5gz6MRkbJha66n8wyt+R7x
TdtDdSAjD//ON8TlohDZeSJlimxdii6szq83ttRCnsNuGZ86jqTMiXrbWffI9+tfNMgcB8Xm3q19
a/YaeVGLFFV+nWM5sGJC49F380tAodtGypWVcJecR9qyOTw1YsQMFdkgRxFOVpy+QQi1IPUuF2uj
RVRpA16Dn3UfA6Fs5FHAAN+5cJ9Lx68exxS2zqhTyCw3Jpw30TjAJ0Xk64PF2fPn3LACZX9ousEt
kmEJhAQGHkrtD9cdOdB4SmAM/s+85HCzqEcMehj4RPNzSEf2TE8T0LXMRPqFgPUpCcVhE1Nxw63M
pDt5uvxUJztCYM5Ci3s3SYrMgTfGJGfFNHU3VGEtwFDAx8oiHB7spZs4/6xySShkD3+/LhR0+WbO
xWjcyGr2zB8Mn20MyZ2SPRqF3sNQIeTfI5O/o8iru9a5tWr4ZkZX7RXV6csnXaVf8J74HSyREGio
2aT2JcFQXGF5dsuhkWxJgu7jU5bGI1pj2G5H+A/MArWBuLyiWet8RxJGesDs91UrMs5/TOiGZQ8A
dOBcLgGA2zcDoxe8z072okSgKMOMbR+qvc8Akf1vwLhpwHjmTOwQyZDEbIxsrNk8a8FjuiCmCiGJ
O+xVBpkIJgE/G7LIRlX/qsflaiEPgo1OUIL6QwxAKKrX5xya05em+Lc65F92eBO2Pt0df0ewuepq
mp9ptK+rY4juMiDUa6Bp2UyBEZ2lx3qF96EjcOSE99bEDGor9oGP9OYrHN59+K3NYkcqYEYlShV4
pCEWiycfSdb76bxKQR0JIpyHiNvdUYYvlcGXJWe5S1S+qm2BmS+/HrxERjLtpShyS33LQtWH6OjW
9RDQtZBPFuXXgZBfABx5SLl4Lm1k1sVXWGK0wwng4mmMBXYb/3Rk06OEpiMHikmW+AeHU4CDP2pC
2TWIseX9Y3n63bO/Rpf92QK/l+njZuMcqmQgaeAe1NssVPlZPUe5q3z0LJWMP2GH3m1u0GfX+gGp
aurMMCcE0T6YZkPKAgs8+NamOz3W/a/wv3EsJq9FpBPH5qtyrjt1jRarzsbCCkQZHgCC38Ad8s6H
aP17NMqWq1uosAOgTG63t5QXxI1/347n7hCJQJHZ/V7jepqyD/qiLIVOzsCw5yh8SayEIBTp7aNB
ECuf/mkoFlRiW7Q9Bp5fzoG434/1a6mXRc20IjEpVDigr6bLnv6y02EMFJuC/iqgoLMM77xf8Mz3
vagi+8C4QnosTcA1EKUkIJzmHY+MZ4JS0jc3iEUfOCbxk3VOWQ8ABbKF1DVGsDZvXAKjXhHTsFa6
fHCC78WzOx1jRTCOpnJvC2IqMIfeHxta07VmE9oJFgK/qYmgh4oJg37L6XNoi+kUWMexkRzObQEx
SxVGeB2e81itW27yCNtADJ70YRmUSViA/XUwBuI5ZBFXZ6yh+4gEep+b3X5BcyHk3wY0EfzZaO9z
Ju3fHalGQy4uy86kTif7a15bYJxVoGV8lyufJ73RagPZ3fexBCNFHM+7YT1EL4y0WNMikduRdPpe
5F5ZGoY0YslnHQnvi5mFYlSuSBSXZYi590wDAGHk/UWKdVVAVN8Xom7caR+M7f7Nt5Wl3i1jdb3A
cKLPXcbUdrpxpopwZYxhRrD2Oj+51qfMHoKULENtNku0IT7b3qy4m1Dc/K2nWWXvZlbeV+V3o/vS
N1C1I34ZttDZRhtpWJ8XlSptm2raGHRGoDYzpwTogCUA8z/0iF9il4XryI9Ci4rj6KOVxhDJ4XIN
2X/8YO/yYMjrhzFDdueqeyZnW63x3REcfOTQKcnYEnxXAGOzgl2OxDAhsCwMoWv6S62GMe255SHH
CRNAYk8AXC06atgHckriS/5kNnV+RiDQw26q+qLUIgxVBfPN/d0ROI+WzdocySj4jL9Xc7fno9CQ
EhIapuUrACAMLEmBKla1Eev/zRgBtkJqU46r+z020GGqjiyLoyMnr0olizXnzkHd/2mEM52z5YkC
awiR2nR8GI2lxllPJQsdGKjfMQqPRFi+YBVxghY5RympRMnA7bKxibOzx3INXbyG2tlU8vRay6Tz
u3uRJeHKhX6QVplE63FLIxydp+1fAH9Pv6W6nZp9nVYQDdC3WcRCwoBY1dUDtgRlxqxBtf9UotVD
m+sLWZDLRbzNMvU11DDOhL0tmSoRgrvBT5kVVTjuexHNehJNM6HQ8AxqHLIddbAR1UERjRy7P5yy
BaE2KBCbpDQGYFPRawk4Dg/9xZLMBqP5Tj9h2tWHECcv7OMvZU9TOl0WObJ7BPPGMrgiHUTRP34c
rw3IrlS4t2pmSHIN2sRfLEW8Y/3kt+sEqtS0Sl6kKMUXv7GPC1ZpQB+xyaVi2K+P50lvVJi82iDg
Om6IJNmGwnNGlYoI/CtC3Qejx8FT8yRvRKGV77AqlQGcnvOp/W8Hi2P9KfAefUi5eUIx+WePJ8cO
temSmfuHn3nyi3uI3kB1N6sM8TXfc27G8ZQLyKMG2IsUhTMln1JhZBViWkst+3edbKhEU+z9U0K+
GpB/nEVVcKdrgJppyW0BMBtL5fnIB1gHdFCwCX4bJowy7LKa/0wEleaU6zl43OK7BcR1pIB5Y23I
se6llQo3jESGkgVLmsLm8ebXgplhX2Uo98hrTdZ5F/YOknmioSGlS4tBIVbZ7kqw1du0FgHiyRzN
9xAf8R4yKWMESA6XlVKKbzL/SClv2pVvkQz54t0mXL8iYS47mSTd+xJLm5W6po17V1QekTW0a0Ot
lznlGdN0JRmPjmVubeEJwwO4aZX227QXHhKrRR8iatckLJfpYAt34L0Z8XLh1ei9nbPiOW/nLiXx
V3hmu0DD3LEjLF04fV7batN+CAiyBKz+SggnO3FaUeRkA+gnAImStk10MpaHMX0OltPeLEJKMyQ0
8xRVjpzmOBzqH8ape5Ot3ahBeaxfAvWAjuWwIEE5ibybOKKe4YZ8QyXgujYLVt4hUklh7mQsAC5r
f1Q2LL4iacHQMB3JMizGWsf9QUmHc4iBSuwAElrd2ViZdRxO8C1iseL5sNtQAEwsFZ4pHQ9Z8dbX
jw3gV7xGDlUiAoyrMEJEmOlLUGmoi0hpVCatkY4MZZzCKggSqhjP2Bbl3rY/Umt70d+mqvuogWQD
2sDyiXXO2z+uV+mIIJnycccakCjozPhu+uv9J1ZkfxBpkoxpKxKnUuB84BzqZjsRMpZCqIugGUHf
hRW/BzFvXtGVwlQDgReAXAfAwTNHnfK9JkHHAO81dESwJESKBeSygYnALAbH9QUfktbC+qs/zSAg
hLZ/QdBnZSnMbeD+RvETPnF+D3XxDU79fsRTacSvQDK+LC6u+WXB5U2IniZHZ0M8HtZCBimXa1Xi
G2A5l7RFnNE4lM1N33FRSvXGycgKkn+VZROPoTKA/LyEaULeWLp5P6QFrcjPqsKXD1sSsDVEcl8X
8UCLQ7qrNj/rEucqUdNLReQNYPAicnNiIg+5MGjKC9ZUKO5+prCHMgHs7PMNNBOTC2unmcbaNJHP
U72/fgz4yww8OL2/GZ88rFQcvBOUUmZ6p0TCsmwbmRPZDYB9xKb8YLclM7CHtTcBRs6MzcMIaLpe
TMUbAsptPWyvcJ255xysHcMsVae4TDynQvAiEwqHVxF/hgwyKsoDCjDt8uOXa3fVb0I+MjZqZGii
5fQAImIICLUZRpI5FuLLc5MGz3Gtd3q8BDUbITAdPqCi+gaTbDAVUz2iaPXNuOMpt8rurDS2K4pW
zwNLL/tPnX7u4yZ/40ARSwda04Z+jzO5gfYj8bsIUmnwqeSMycYYdSXdT6+Rl2Xbo8Ddrt1HdfcJ
io0mgsErvI2QdxxR0LlbuVgghw3dA75+nu7Mc1aBXVv6iW/ndk7YGQXDY7/MRW2Bd3QLyDCQRVdx
0gJxurQMD97plMPn+wy1NAZA15x3MoiTZPkj12QE/7dkgZEngrXJ7gC2RaYjqL5ehu2TxhWiYr8O
fsCIKidxVNYIMSwE0dinnrdaciNL3W0dwd43oAOLQGtGNZ/PSQ1wHD3nJJs7BmMzrt4By4bta1Kz
FuhqOfjRyy0voH1q6//TIOdV+zP9vuYqPgAZn5DcmIxf04I400pDHSZE7oaBx7Jl556KxJ3kcUla
UZH+Vz+3F2mHxkscW8AyS+8AyX5jLAZJmY+XdD8G3Yfzv/VaXls0ilomoPqmUWDS5I71XOa+9v8n
Zpw7XX8nr80NRcD5YCQWDM2h9GwMVh472Z4a7XGi7CUOTPYy344p77jNDOkc7tdvpfJklQFhhgit
WRUzf7ip32oMa+Mel+/pnfBE9gaET8vet+9vhYQXME7xmSe6k5e9mKaEmoJ5f34yv8s+/DcwLb8P
2ZG37I33Ub3yn42Nn6aQfALWdqcmE873K2MuS7y1OfSt1G5p3YlnD2oCqXZrmEDeRf0F7wTFgCJ3
FmVF6Z9I8FjrT4/L8Fd6hhMz9GcicfnVogfIZQwUHIqeSHMkYqVlXfBjeR9EnxL1boiHd5ZJSTwS
ixtxQL1T/hJ1qGNfbVtXIAI0xA8LzRxjsttM3A/Dw2m9PElClCb1bRZcIcy8gFEZ4bNHFrYWCuVL
dVO96sLkw72KRFMOL4BlETCVF6Aqj+Y5SKFzXY0GcuKksN+TsOrhhRujQS+H3nBk4Thfi/fQxVo2
7driD1jakDSTDskLrGhNJ4+e5xNwIsILhCwI8bIYc5PI0PJfr5FlbRjMI4U/px8LzvYnJcOjxOI5
qfqY57gWcvviN0k2E3DQHI3Xyco5AADSk3qhwnB42twqQdn0Mk1b/prDa+6DzystlFr4TZeYwANQ
UTrqVOYEsqD4mNlNqiC1FZsAbBcmF+IL5XgA+E564+3L6l2SzE8qOJM6UO8clDYxQpIJyTJqvo2I
FfqnCV2Y+n4sALYmn+UPgx1l4PcBHgV6tS9g9fGvaeTucKuuniF6VLI1KOPnzLcp09KiJTiJFvBd
YK2m3VgsBMEKOuGbNfgYvDKMy0V7loop+7baMp6KYuyweF/MlxGNFrIa/7q3/wQucE5JkFqPg/PT
i8bE5egpE4QF9BuzB9bTd6ihbn1S9wo2w9UAYi3unXD5/w0iA/NRi9qDAo9aR9XtaZzP87GMKbVr
dE83FBhmHQna2Hac7FhXyMKFvUKjjdQ0O+zpGChdLFRF0OB4KH8jevuSwX+3SdQaqD67uqADryev
3rCP9rRkcHJL0oOcbRnhHHXdyruOERsjP/WiCa1TuGilKUnT1GNmrpYmLisMPc8LVDDLd8uqjuPL
fUqq64hKWEF6hHlTx4ytSVjnsGogOPUeoU37JUvdhVlbCelL+AKqhmmjOtJJkpxUjpUH/UI1K29O
i+wOQTKn00GiJns/aEQAfcLgHhd6cDQx8EMC4bTSLL5V/Yov7G1eA2cNPm8i9S2zsarwZaTA7Iy6
0YYZeDynWO5qWqaqSSaDPZr1/TWYV8R7WfM4NE7rkeC9qwRGoihAGkY5eOu5SJM0+IaDuXvSTNTo
nffXaZnx6YeWAqksNREhd26RCpj97/MhKdJYlC7xotnncCd3Sy6cfK83kzOukO4aTsbcAXJnLuJH
OOcsGnj2kd2gdRrU0gDJCH4pq5mozQ9SgRD8jEKQUyrAq7+hMhdPCgMVN+7kikGt+13esYzyS883
8ENy9b0daMtkOECDkGQcWP9zChsvcsrUTJyooVrSir1qhDAK3ljN3HwYipjGBz16EWY7N9Y6QVyI
YICjRbwE7SycW2IvnPCREzR4wRbWb9NvD2Z85dZN/Hh7RxkCly3lnhta5wkFXGecmdeMZCAC+2td
PJVoe2FFN+7gNZSTQMK1EX5kThgCyV9Wwm6AAAWzaO763ZNcbK1neP9bUwjozCVuZySGbPP4Mp7U
te1KHUG90T0UaRVYd3k712cqu1Euf4/7uwPFwR7RJn3jHbMf2YuAVUFJHrRyBdQ/BevDLE0nJep8
fQmPhSZQO4AsEuANbEFG3g4xbaHu/57zD8qcPP+l+u7NnLFPXahtzSMyKxcTjGzYTfem3ln+LD8c
T6TmVQ+oNZyfwv9mIOE2wxNig6WPZvfcX90Bbn6i2KlFoYR/NP+IVWvIWk0ZVJjYNaHbfX6PhwpM
L85HBXpgR+sk33CykOxbSwPmvwFn1aqyc4EAn2xu3zVSP6RW23xEiHt5PXboNK5Sjj5UfkR8yeNa
SzVM9a1VZ79vlRoTKe89wd+qy2fcps6Y3Ryxa/aeFjrbBnRgt6pqJ1iNvXt94t30pEpOYuAcEKvH
eKMXXZtjszDXsyTlt8QIc92U3tW1Ez2wBm4lX6oKR6LAw656Ea5Tlip3Ij7fMR9WiH9voEqJmWfH
3u576Gk7jDlfOkodMVESWVHtcA3U9XxHii6xRi0D8ymL4skhGjwtZ4FNwWU18HAqATRZ3YepYVLJ
N1zZSd1fOIa3MseG6N789QMwa5keWU0hFhbR9BRYq/1quz7VyD75nlEVCO9BIkXxWdvt/tZxVqlp
VbN/UaLgh+4j+HYa8pZBw5v37wzvLxqUYOUFss9J/SJTWn/7Jc3dow84Vbi2y41ExvgobjlAHN5/
WUIIj8PWYBmTTBavH6VGFUl+tgUq2Dk6MXAtg1n7cBPiyzWR4KlnwLQaoOegpet7+FDzH9iwEUZu
ABOhlwRbp2nfib2mRmy+shKzq/r4WnseqCqyVc3NvDTP4S5waGiFJg9XhT9q9v9Gre3da27KOsIY
xaLV08//BOpKwgLq+COO04+QcZ+aA/crzTPmuz4ZMwtTGpc8XEYNudR0L+WbwZm61ha7qmbDIi3D
8Td61EAVPfirhijjj33vLUh5dh9V/EfWZIPKECbzHwKGykGDiGyXnpX/E7xW5KJjPrLcTY3gDkGM
ZKxcTbqGQXDWZyZhNkpBG8osOioLYRFRq7ynlDlE/FrBzESI7juZex7YlsJGvP8Fbd0lNN31bigX
1SCo+uy9D3C2IePQNU87mYvar1yQZDa2swTEmFDIFjBEnp6uGntUJf9/SOOmW5h6AkNqjnpcXohU
D5DoCm7V2k2DgJssxrvttU+3vHkLRT3XZgOjw98uUCGHQgstYI9GhEZsB+7nxvNgcnkG4thpi2EF
t2qsjZWYBf7+IzdxKaLBmxBLDr9kfwiLK4+x53SCbjtQXL0rvFnjXiXSbGYVQP3i2z+HyHDAQojZ
9sI9GquWp/6FAu96dkidSyj1tbVmc8ZlU5ndCbEu/+sJgmhMNGTgVpdt+1IGdNpZo3yxTeW+6QAf
xFMVc4Zm4Ai5pN8DHRbOLvHMZPSi4d8TY9ATCJIG4wDFxcR55iUR9LBMfP8tdFILHNy/80qEd8lq
nxmkiwnuZxP2YlaEXP2QUOeEIrAJHQ2PGOWBX9H3jDdeyzsY1ctlzHDwkQm2kSvs5WlYys1IUzpC
WCOsAKwBVCrWVU8jln/t+9NzIgI2g7gTg1JJEFtfB6esKcf6W13sD/c/oKfoGsBbzQnG6jjKv+R7
P0QvsK6xdjNoL1J6sfeBB+A8K5sGKSui/aOLFiOewC1lspJ7YSD8S8vV14tditQ2rf/AzaxC7B1N
bGUhDzhs0vM1mnDNgmHRxCXHZ/SP2WKclUnyTxf2/LeMCSpV4Ce17TOb/GAudCql7jGspBOezQc6
DsJPT/csET0VVMVqaXzsF3Psnk7ZFIVPkSpcMW9So7r+zoqtkjsZC+xtsxTVF9jPe5PlTEaHGYvs
dfliShJb0QnrjrhchlGo9C9jrHIL34J1i3n+HJrTyiaMSBveuonF09SjAHFAWoI4GAOkc9llbii/
Ofhd6FulkTP0uTvMqO5e6xqmQ24UFTjLQL8UdZQZvcTcTZgWtOunPzmECj6Osnl7tvnPgrpD7zyf
IDvrOEygY0yyW3oLnhNXvuGkzzroxYVA2WtkrQFdcRhjjzsfsbukJ0yPfKnOGpRx758DrjsFJPv1
KpNAmJpokolvNXwbacQZ3aU6vNxgwEtIIuDZUE4q7YWQHp53ItCnI7o2EmbdJIn6Rfc99YlMbxds
xqJVbUVI0DefIpb1XfrPY7F3LIbxOcIiNuqxcIfVoM1OANmFxnq5V7omf+qJKSpVWo4SMM3DSsUF
uaK9QKJn6C/wEJgvZ7KEgzPMHSr9oy0jvhnQ2zm6NNPiNJ0MaVNLavfKm2ZmEA6NcvWUyujjdJTt
foqOyFmgq9auR7uwHVaElmxOGxBsniqIJ3wqzOuZfnNovsdUhXA7JPAswl34P/BLumQXepoFKsma
/V73MhDiGzq7EE/VZhMQY65GIm+GSzp7oeDjjlZeYL0Oo4qlhRLwN5jFMiADW7VS9LM6xlz6cPqG
PnVU0zucNsc0stX9Bd7KKTQZeS30B8U6h6BtBbisDUGVpqzmHbQRuSVwvY6n3DF14EMA1QZggBfv
721QTTx07MUUW3+OQP6zlfFZIvWCjo5+c2r3ulV5D84lNKr9HAyADlGMFmG+gLpjuw8fenImDn/f
j8wFQozj/TFq/2uaYKzya0mfV8PNlkmbWdAoS/78nJ3S4BdQ5JHmzNpjjdRK5laaL6bpGGReOPt5
sBvMYqMTeyDipCFGJyKcUvrLTp//OERZIryueqSij3yiKamiJ3mDSQrkvKuVitVgKNWdkLBRIBf0
EL2cg6BpqGiSaiZUf269iNUXs1LWaiTUjksJDgzK1NfeY3ns4yDnvcifPVFGKQ+mfPwwdU90sPWA
KPTZX2AJrC/LJaPNFQg/73e4qrg4+kCE72gaSmjurrJjdYXG6Sc4cBWZrMZwWsAdZDLdILASq5mV
bl5oTzHhPfRXw4yHeed9rRW9sG0GIqGRhnogqVznI9A+jefBMmaKmN4SQ+p13i976/2sBc7iBeSC
REgQ+9/5fyCPCg7u+h8N8HDy2A8T7ND/H9TLvL1OckO4jz4hFvjExtHz56CSOyWEBtTg7c0xUMDN
E9Edoqt0mW1oqF80IXmS3yzNi0oPolmRFIUrTYzXqwFSa7wiTzj3VAKg9MH4108ilVNt9krKcbh3
g4tKHA+iIGxi8k2ksbQZA7RozKPMWRLKyJIvvYUku61zzF2KoBA7YnVgNWAWPTR8I4G+vL19xODA
9jS/zyS1rNo3z9J2SnOoaNtmm0CXSDTQjRjTd4OjtlspZfBs54JigEjE17GESgg6wlFicusdWBGm
4MbdxVqPONSQ9Yu5/mkvBcyGY2pG5LKrxX5FaOd/Y8AGqt4K03k3ZYuZD1i5e+Cbo68gDOt1mjC6
xogCnzEbXjugW6TZ0ZhfKc6WO7mtxlmTRHdjl8irkJMIwlNkN06UiMIDb4cOSOIc6REVyUNEmlVR
S2glQX3ETUjgGe4oNGDTc8sMkhws7CuE6JlYXJysbLVA26BQVMqVX4QNuoXt5Zm6LQ78XNE3aTVE
awVP0skG8+NyApH7vUVkV3i+vqH4Q2NN0hVzkV/WvDSmFzTUtYQUrOFXoJ0O0BolTEr6FiIlIlmR
tr2STN+2QSJEi1MEENE4AUlM5rj8h2HLLjeg+XcsNU/3PNlxcXrkDBR4bNUfeBeTgJT4W8dyUpFx
/+ioReIG8J0eZoIoVVNSyoMKCy9aNvF3JrAF6xPq8C2/GoreTdVwh6VubRa5uQD3wnp2ptpW5/Ci
1afEAMhD6fr3EAtJs+hhT5K6l61GuGaAOEx3S+V5vmpHPh2uYqpdArGRHtso+0u6+jnSdbCZ7mq6
vAU/WTIrRISxPXrrVwGQCNUDnEmRLnilhmVLNOumydANfS1+7/ryqsC+TfmA/VgHqqDQ10pgGMXH
AfibtiOWWBO+nbmhbNuX4/hWQIhuz+M13MQs8hpsMVBlvF//Tf4x0fYjfN4CF42wKZPCtU6iyh1x
/ZAfONNaJjWMbtLI7cghuEfhc+S08njmg3x0Iisvln1DHSBZZMjPsUSSYzIr7VOiPkX/0FgVQ8eg
n+OhLcUOrhcxEwCRnf1olGJLzI0lQ5U0Xp+iE1cqo0VlLE04ZCSBsggK1xPpttgCCgdg6NNVxC/M
So5gt2kwDw6DbCkmw8fsMtHzmHZiFExJkutdF/vk3Kus9i0AhFz0RNhAA+hkK8SAjVwO/kd31sio
GnPTkeb7OvfXeclhs33tPkNJH2CC4PKT4+Z73hGImdsiJxwBQirbsxejeCsM7kADvB/UlckDiFdW
Av+3w1wFP8YFPotQT7wzibQBeLaRH+fYQDo2DRYGuU780MRxI3K+Qk7rPsV9E6yUiPIkzeJFgkHo
hILdUKurbcNTb6IEZYgz4tdxkl93dSdB2XJdRdw3aMbczPF+iZkB5V5+SgJLWAxeAiMj7vLo3PMb
kFGhzohitUTFE30YgD/fC6taXVMLQe24L4a638667RF2EBpR4fXNRgMAsLUv0VkfBueULQ1vYxFf
bQg5PZn2c3q7l+zlmuTsyPnE9kU2SinhvfbGe2qdPxLHir40LehBSfr4td6MmPtcWuW4QRQdvstk
fkq0y/PcqXjOfOXIfEJVqb66ERX9a7H1HbcOe13JY4Tw7+oumr1+2OEJ9bE4nUYTP2CSOxxLAH0h
wDRhXcbmrlmVo9ehnLd+Q2xwNkNs8UYBgTUrhtXpjPniTYb92wHdUuJuvLeLvQGVFPP4WQCuo2y5
Feip2Sq1aB1xH/K4stv/viwOSHFVNzxIuKgvzt9lOsqU/rB9g2riFjwe53EGxsamuVi84fQhwfSZ
jebRmicsSZwdl6BuZ+Zjsc3Q5hALNGS5NkdRclYivHnRqIhl5mPpmuXkeKGsiuFiz4Whq0/zPdWH
o8FQ7f70/j2jIP8XwtksZUWWKpSgipn0wxa5jp4cHGjwV105lPGbP38ay8LJ76Gqocu/YgcmM1Wn
sm9UCy6fvs3h6abjEPaDHfm92Uq1lftBuRDQFMLcbhPFJMR0/WbN9TpzJHNzSi1e1vQxN17fwdJP
GnZXwLlJ69zsXqrygoLpN0B/wekdM8FMCHbsj9bWbOKcg6YMvftdwzOO2LBJbOd2K7sgThivA0yO
JzC+QJuyEho2bIyxrZ8L9AL5RZA0sA2BQFMI16PiLNnwf1hwVX8oXO9QB+YBgnjoZf9koZbeZIbQ
dqenceyViXLE5YszV2mKAEqnPqkA6eyY5UfvNUdj/kpbAIMdyLRhxlbKYHgIEpyPR9bN5lN1jfKe
wBkeBDneqpbI3SH6KIY60QYlPiweC/QOi8tpURTT3QiXrNL189qodvxxmT1E55PPRb363wnvaE7P
tV8QdN6UMOS+EO38mf7ANQgAMWUhugdqU5WSH2zPgqlX7a00d+rvc0/1sx5xGGyJ+bjevCwnXPft
wKsdcUnOd2fXROW2S5R93OBTOOe/4fIF8lE4HvkSb4jVfbfbwySyzTX3G9fLReQZXTxxe3f7SDOX
xIjOIAEoXP64/6BY65mbhub/vzjb3jEbES0RxxkWJTWfUNwbPGJlbKkW7glcg6pXav+s+sISYA0s
FkzWyPhZHcEOnDW9iClE/0M+2mlBuXizgOPpqMRWvenskIquJ8De9D+LBhwzLJ/umrHLr5ddgQ5y
nfeasklCnLjgHVUN6SiV7Cdv8nP4mvT37yzm6GFovUEHJ8jLAFWAdKsPhdlogxdygj7PtxdQZfpA
ZKGcEAGwQ6+f0Pwv++eUKxI6C67tzSMoJl7rozhxYZw7p/L8gDHDJDwCdndY7e+KVfh9agaYC1cU
HuGcvkzSYA7wawn7GC2HSXFKYhuFKc25RwMEKANl3b6vfkK4uwZx58Vb2gMGIUY3Ad6lWNxzp7Ze
Zw91D34zqDeSyN5dgz3BLdkO/ju062crbWkMQ+p/LwDyI6owOv2m6tDBGMM+/QnR7T8D4kybOFfx
UZHlAdPox61Ikb9FG65FkcjhtKDdJ/BiXcs6mni09xJRLQ/nXK51/63ofuYHxwsGYBL8di3LiouQ
hh1h2ciZJYVUzorGrzMNIafTe7VHmYKDU3i+sVw+ZtjB8yWyKI7mPsR0RDoP4OY4+8eu7ULWvxOt
Sr/vkbHVs4v/wixoDSRX1ksSEW/fEJPEKvvx247A9U9WwsNHKawcTeV+F+JStlsqPDO5L1FRoHaT
v++oG/0sGqNdnv87ETV+bjPT6uvDFUBZ5GWj+VIbE40pNyPVtRvlCtSErU2G0JP7A5au1X03y9Fk
J52uX8qJcFoqwr8nLYvNcGCGe35ETN4BwPb0Hqu8+f2X4MGqDtVSHZASvyAJ7xdrhamsW0Qxs1Xq
a2oATKY4yeRvYDMw0OH60Jqanhxq+InQRgZrmza6Zu1k5JY2wSeb0LYJ0pTbZagIQvOrXw14uDsl
15dda/A39wVCs3D9zVJxoxO5mERw/HGADAz+mOm5O5+szXi0v5J4/HK+xqVWZO/ZvSuVggNdKb0g
dOHzeWMFp5RQxz82ibhz0sc79zYG93Ih0Zu8ScmEWdp3QCIX9VjTtfEJljwHjfEYXq8rn/QCoQB1
c+fCLS1AFaJ5tnN0hBPXed7m647nP0PeqOKdr02PPpXC+GSBERSp58biMnqkPMiGP8CxIlmmhXUN
ZaveMFZmwTp+/wp9gMDft+7mAHwpm1MF2HQVS9rX1BHRrFe9e2e8/WIS8RzdKwYSL6OZlPm5CrTi
JZo3mD8Y5v6D+AMDqKRNL7Dqxg7stWbRJZtVgDOUYjPNCk3t/FlH0S5BulxbVJrQRtru2MTe5ZMv
HfyZfZZ5VbH/9Zz7e7XaqDXxM5hEVSSS/S7pxaEtOhjsCadd901SI68PTg4IKStK87KfOh8p9lne
NVQxztolDOB1cN+a8qvYBNykzskqucaGf1d+abUXyZUAtGHcTHLWhINIGnc+p0pjFhWJP4nyEawJ
P08mWBBAZPHmOx0Dpqq873ov1KbhnaY+Wa8IHl0HTWjq8yCJHLzCZNX40YBn7BnZV1iBauto584A
4WqjY9rqV1NT2ST7AW9ddN/VMf8IPzM3K6iUD11Wc71Rbj+PhBeMC+Ei0Dmj/qm0cZm0L4k6nu6o
zFvSxzchzdk5/VgrdZ1CxvWKHFvCc8H+93Ai1R3OK+9h3byNaxeQMWmU6hplEvRFo9sLuILf8mWx
8Vo9IZiMwAXvdYy0pr/Qp0mafPu7OYdN2YtBQruCqtyfa6psVTzJ3IWvFGomrAFhY5puupvGPOlt
tGFwYe5+yVgr97VCxQld25mtM8A+CtS4VcgvHJF1zlev/8TFIjDFoUd7d2z2SY1murGvXl2mzBSM
7FlQIeoBfPMoJTES9W8oAulpxMI07sc2esdwjIL7CNyREu3PG2SHclxcTddZ4CWpbt93gtWWkI/u
hAi29adfGCZYDkxcxYevN28wlMNRrNZ1IEq14lxy35m3BhLIk4/FhqE199+MpFI0P2qbYUk5wt8l
RXyckstXnJEgJSGiLD72fVa91Mlr3pbo0rPVfpS8ch4XVbQDiCTaJyGBsUNmHHfVqt5YFcP6gXWa
SvbQJiVCA37vUwwz3plfeB3+71fvcq1UKO2w+CS9zhBcYpk7cMmPPf3jwAaQRzTZR0tqysDbkSOd
c/b8+tPv5/or091tXi3XkVJhFKoTwF+c0w+Q+EKTIoDHiGoAORyMMVWT+d/Cd+zYUV1ro7faAMWh
xCDNNCX/FdmHbIqXP0SJ6WX2zigL0QG9lBUQTEZah9cMCz0xDpq8zAjA6P6Go26KtuX6sVXyuT2c
VQMoe0wIiIuRMvYeWM30oUr9tDfMYIxXpWqYg9LhUC11CPHYkZLyHNlLi2FNVr1Kw1QViopCW0Ea
wl4QbvBxCp5sc5yj2U2Kf/vG1pgSv1KrTCdezNUDwz9s8Qsr+GDLTX5x3VzMMRbgdCN9Wxarr/GE
1cyo2UvVc6ZU8TKaIoQ0OiJDXGN13X9UyvxKusN26OzzwVCCNliRX41ezi/aSZKq48yCYu635UMj
G4n+Y0HNsBAS0VEolva98k2px5M8b346g94PPjVqWgPYCKJzzZnlCtV+A60kYErf2JM6/1gBOysz
cgLhMNr+zhdHbLq4e5VColnEMguo6ZFxbVI1a0wq/0PG1U+8DqBRNeAFlI0Hh4mNppIVYp3CMVYK
8b1nGbeBgpELWbmZvsupEbpdurbLSiAyQtpiBPYoi8axBOz9/WJHEqwdRwTwFTexSwO8bVQuk0z6
b+Y9QgAqOqccgmc7pF1skMDwpNJxi28BTAq8IhaqErraPAU8izlKWVLzap4oqjmL0CRZRdEvoKB1
i2m71vVrSzBjXrS2opSlziYOGOCZshNEKJNRodtTTZAoVH7gvK3WeljsuIlReY87kv387WOp1oCb
MRcz5jGHxN+xp8Ypew5iHAI1CXkdrEouTyy0+nW43s6iyakKwry071nBoEmqIdhzjQpbdDlalQVw
wp1KD988pSq3LJNHT5UTALa7zflDFdFFmCOnjVj5P3VbEym6ov1CumuzzzWDV/z4toqsVW4vqO79
5b/0IUyFn5ExVk/EHDDR4y5Up21MEX2dSw5xj306XvGpCS0gzBzoNXB60HMGovUKP/CKAdU/6M4s
ixi3LO6u6vXAwrW3Ccf6f2mWALto10rDooos+o9rDtkikKe90y3dzvE3b58CDjyCKSEZ8XlbTJIR
n2vbjHmVKEzu4zTy3ZlwzLTvCopONFvomO5AII1YnPl6tj3gbCOeLl+FQb8wxZQT6pY9kCwBQJfF
DtCg6bQpft/KsaJXvFOzyGNsryy5Kt2htkb7Eh1HanrQLEzegmIjYS4haTim1oF7ONXS9dcr+NjK
fCMG5MOnUtnB9wuIZZ/nP701GCGx2MVXX/6u3lDeOg7R/ROcPzbntnQCumlDJRmPZDEJTAc15eFM
RO98iuRdyZpi0Jgu20VglosRmFlknlo5azO9BB4jyfOYJmXtEceGQuzZeG8v78hdq3d/ed5cAvfp
Xm0QsK/pz2UpbHWHOttTFYy4hMsDDCKxM5KDU1casN0e/a3OqchlnBMvaSnJx+8n4nWZvvJKWLnk
PzPCzCgzHYfPElx8LF7nHxzEoRtghfpGJ0Q2R3q7nHgKFzPLmF51bdLELRdG/DNqo74+lPRLAoiD
9tDyqad5sRFS5WvwHCKCm1deSqYeTKd3VKlwjYap1FUgXqkpgpVkqNnancpFV+PlfQoQDor835yJ
upRQSVWiuLQUELyg4KDglFlfRrrBnShR2qDZCr0R41pHRgyxrI73Sf3ynXYo7Rck3/ClOIo/gEYZ
jprS9XNxJ/5CBsAV9iGWpO+KnJ+2971EGaMIim0p4npOUpDyXVOHj8F7gZpyko69TH6M7/Ju5bIP
XTFYb+w1ZOFB6Z9J30jGuE+SGvjEEECO2IyyRqZzPOdOBvuHZNbB+asz5d9kmb8e9faLpn5PN1vV
oHrFgIx8E2KKojc4w85qFQ+pogk9UJtXj9kvJxhMAgMVtaNI0Hc9w6eNxqOpaDjdTYcTJ6uyQujI
a/F6mFlW5402zFdBZkArTNqF+Mc4bR65VAjSIBj8UKf9y/noxMK7j8M4M7d0UCFmd8w35l3bCz1w
8B5Q87YMlOaJjNxXcefeaMn8mcpfwsXqDH3INTUrPaOEofko+dKZzqXIET4u39OGdK0P1qge5yjc
MpL+OAHxKuMU28w6E9P0la3bliPDHVL7UoB8atziZ/rM4XU0VUBluiCOnUEQa1JHzGmgRsX6/bm+
50kCfQlMUykRubVg6UXZ/08hpK2QLX3cARHKk2nvibC5DjAkbWo05iFXRc3vdT0NFQ/KBNnvK+nr
jJdVMQ3w/GiKAdzhSAiZ0Bri8vuRK0UVOqBJHi/Ol4w+P/LjwwRsXIu8aZ5o30Jhd4FaUmRZH3Ht
chMX0vWrsoSX08OBa0EzKZb1HGeKt+mrKEdsWVyUmylDDrCOPFhlNEFt/V/SJauHEGC6Cu+Kx2vv
nJLlT2HhwjPIXVqONTeha9gDfNgunBbZmi5C3Rdh5I4hH3E5Abfrca7plSuYI3Bbj/mrHl9mLVJ7
MpmfiTiY6x7WXKbIi1cV/KozTyTXplf9qLTp5ts06iyoX8mU5ViPu+9eljY2PklBtNHR9cfH0P9E
P3FiMgvbaebXOtZTR07PyF6B+hBpH/UcyaIfFxbjzWvlAUPq0OCc+OD9CzjEduMn+33bRRnEZKHA
KxZcI6kvD9bXH+UXcunGCq1x6xpBMdd47NYFoudZsvAT7BAfQZyjiDge3246ME9JI5sOT4xKJBWr
H4gpB1fgMeMHLdp+Qbt+3ZRXRqjbH19qqcLDwXrVTI2+2CqzXrJYk9vryR5l97fY3v2z8ZxeTAc8
TC0Zos/1xBUT7kANN25lwoCCAW4AIL7K7d95VCPG3TrkiduVAj8TBy/PruEkbO9lv0EyFtkwxzrv
OxDam2Zshk+qBK2gE/nT726GlWXpvD2VFioQg6PrD3UBDXvAeifj/bhG4oEPs8YkJi0G2lyJpuLA
aLzVTxegZLz03xk7rGD83+0cXL4m0Q8Og1iFt8zwB1FcCmzL8GhVPZlda7NhMNX3j7BtfBOZuhlB
2Gdoc8sN037s5OPkZFzCg3XEGOdOSsUHkPuE0E9o/T7jYOOfDjRwpgkTC9OwMnwscxNjqNz2DBXW
VdvU01iDcBaUvivqxobeBxBLpqa4hLJ5Txqm6Ctr9/AY54FkP/5OTqeme8K9fimrQlXRzcin8WTK
9rsQjkRAQkpXQhXU5OeJeN+vfLSYhJjoWWShGQU9FCyRiQlwu+1dJ7JscTyI3TSSIxQ9eyz2wrKr
Ttip57fCiiQBkMdRpXuaulz6SiMUqL3llbh8i2BTlTR3LGGiiDgenAuz6Yjx6IOM6T9ZpuQhbicP
lUVlQQnyaXbopjWcRVlAl6Wwpsz7B4g3W8RDqk4EtCd4n0cgXxXZ6eiYPAZerGwnyLKethdbFbVq
y1eu4FrTDL1L9jg4GspVyr2Rm9YfL9Wj3jX6cdzZ0In26agVwIKMUlT+idpeZvMtWEFP3JXij9Hq
b/viOYJGgdZm6gRlG75L2p6LQpXmPgRIh93rahUm1f1LrecuDQFXU1F9+Y6kj7VY7GtE2ztY21V5
eYY+joN1vH8xFkiLdaM1c2d40bmxVMcoMbbVvRD7xOUiMTzKYfHgXhnY+o8+GGO8ClkCHaNjVeTX
pXQOaupId35YEGTOfkvV8MMb+yoyw+og8V1nwcGn5Ng+Gw68eJ5L2ZDDtQ8NZ8QOgK554wt581cG
iET/VkWu9SlNLjz3E15fHQ5f81ou3lmlRRlOnMNWo9Ll3qwfIG/WTEoNKXVwullaEaQnVI6GXroD
TlU1qwm7fpo25Zt4q781AV0O4FglVAXvuLbdb6XZXuTZijoP7OsLrZEcs/Rn9lLVhIse1sZLSblH
umM22dSJvbMfIVKIzDMvcxgFPLgaTe1CHrGbp6ha435T61cS+3BEXElw+IGmg51bF9eSWZk1WNGG
v6B8VLfhRu2Pr0C6lKcO6IMEuiYhGll/iwxuz4pP5xmXFujnTty0xrjCVunXidJWG0uMUC4gJ5Xp
szaU6k/+SpTgFcT/tSPNyuhnX4zbzm9CaXc7QmGI72Zqo5sbq6dDRC9dnqH43Ewbk9Xgc09VesHT
KdJlC/H88WrZwQpjahunCDPA9NE5lI0lknOX3yVBPjMumCYze6Sp+x/S+7FTcuHSQj0Eo6DCjV0i
aD0oED9NnM79PXZZKuk/Vrb8ia5nyuURIZarJdGnAlfjlZ12ylNGuJ1Uv9W6SA7CWdaefut4mDGW
OyJYaTzSZT2r/MZBfyJ1eCCbbpQ90SQeECR1KdttohPUHZzQIEVHfJmxrFNOo1UNM209mxm9NYml
fm9+4Oa+7b455WAzdaCsZ9QVUEDBoicm8d4r5l6GX6jwpvWO9S8JmLLdsVRzMbD5FEWwDTWgJ/Sr
3wLho9QDmv+1xbtbC82Ldz0uPvSTwf9Mwb41yWuQOlrsiJpzg9mKfy1z4iimSPVZmJ1J9RXZ/PTm
w4mzRdk8BVtXXTAEauxQYECtLEFlpNLngwTWoVaWIbi+Eid72736V+MADAzMAYi0ph9+UHilkVSX
upi+Zeeikky/mL/earN74K9PbW41AA1lpbN6SNRGxjc02MP+WLayFUfW9X9lmc+StkNHiMG3uioe
/Bi/A7YwGFf/KnFSL2AA6fV2NVFtY+allVs6Ed6mp7k3igdX1QZvBxrvEL3HgSDIhJ2XehVPxg1p
6XwskuK2HKedM5SSLQfGjM8w7YW1GtoU6enW8vNAYgdSgoVvicS+FSqyAqJOB6JoLBhyq994Ftda
8WXOpe/gIGhn5E0E1s53uW9J+/pHcHy/qFe44jOMgqe+3+WfyG+YS1nLFCUeyBXtbh54c+8xMscu
/gQtusg9qaawGnKlBFEZcqUpFvVKHlkdyX5AUYtJGmp9v2oIcqR+PpKVoV6yeH97IB28OvSSd1RA
N6LuyLLG22SUEmjf3K3JKGmEqLzc5mxcnL5SS6DLCaWxlFU4toZg+R1iBDxuKvLGixiB/xqIrDKs
JxiYemGvobsxKFEGOhSQHLUEeHSsbzD+wY23xQHi3Uuo72gsH9dEQ2bPtsf2kTc73MpZ47BfhBje
V//Jb0tBs3qgNwPLvWsTqv7duWZvymog7pbFOCUGh+J6BQKoE8L5rj7Y0FQk94/1sHl+kxTgQdkH
/BwTlMGz1ldZn1WqU3/AKWudomfVfDXnpyveiFyQQRvem7usly7/jNelljLyd/85CUiCu5ifwoGX
aGXZgdlR79VPYmxedQSzMhe+BL3OrHSwwm67084Th4vo6SkuA2p6B4lTiTJh7BROSZQfKO3NSM1x
EmCZTgL/A9rPkoIXiYe/N0BP/fRmDAIQ8+m3w7H06ZF/8mzcBH6jwOUZ2JgGgoNZD/zFJvZB6y71
0FpVsEr+gDsnQE+RyzbVAJoyk6Leynv0oGcso7dNgeDwlzKSzeK88aW+uwYgK+Xno/NSszacrpUO
e6a9Nc17K+xlFcJE00lIju6wLRamZdZ65p/P28cO+x8Ofg3TbpOfCjud1YSM1468ruklCLjTM5Kc
1Zgsk3Cr9hKTHEJwHbX6sniuf/5DVJDz8hPTA2MYaDQK6w0hj9uf/6shDx4exF/e8Az7lS9ZQCzp
YnhsRDwpHOhpNe+3cj5AHTZS350JPUYoT/BKxhBDq6szWt8f5Qo+/iBv9sGuArt4kjZxmNpTfWSr
EpsnhVND0ZM4TelmfSdqQzsFZORikwL5Rd1KZho3ljGxRWNyl8+bpCFxDmCTu01wRRkoZsE57hpk
ZE5WFF6n0+pfDx2kPdVfqESh8NVQk5YnnEMIbvxg1qKYWqWk55MHW/D0glFjagj84eqXoWhiAw+q
2iuIbiuIDwVCJ+zx05Ra9oDF9mR9ucXcgyinf1k+rSCuwpWQzZ5MmPjbZpPkU6eEKKa8H/Ddt1dS
sPQH5CkzsrzXT4TwawSZ658O3VJUFNFPhYW20DjIXahsir5z9go6f/iN2OZ81rpNDnSwYsNjyFLJ
vJBIgotjtAl9ntzscnqnoM1B+bUNYrYbJrN6/Zt6+FzZNgHWZyoW2jYRGkGOwABAyi4FpFtshPb9
EuJkAPiSbi8KhUz6rcvsO99E7Qde2ntntz4ae2ed1YwElfj9OjU5wceWjxIuokZGtWbpLTzhmzLf
psdQwmZUzNwYCpv3IfjioD21yNST2U3a4E7i9vHxc7URxThUIpER8mdQDEdPmaoiJ8xHVtf3dJcz
peZyY4D4zg9AmlmoH5ZdEspI1nkjxNCSsp/eH2fHlm6lyNp+ALi8gYKBQTP2MV8cQPDjOSCGDDye
lquuakLgG0Y8izdepAMAs9AAWMfzFdDO3jaZGVP0UKl+UvAIRUaIy3nP3K+K23kD0QwphYnIxT9k
IarL9Kn3xhJbLOXgHLvuv1Ok5ePg9KhVIBV+oDjyrM9BvKmx3oxBk4gCVGlcpPiwiRVDl7DN73sw
shHjkaYTcax+/u4IEjlhw6ctJvp5CfdwYHgLJMtICEMDNzKY1mhAqyEa4ec3WKXYesisLjiFlLvF
gkbBjcxUd/0CR3TuLKVK7MdjlO9xq2ohtEiqT90OY7eIl5nHroPqD0LCkqc3oo+PMWiajdESSc09
3DBzEUmLyCiX0CthtGsxIqG/rD6IxypCCDIw3eo0ieCYsYhZaxrNLNHFwDDw0NdgFGMnz2IyrMrm
cF5SFHH9iBy4svTpDK7mhSOplshfYBrrFlEgWTkEAmgtu260yWREH7j4kv4knxUbSrPYmXjma0ns
I49tLKDoKB9scQOgcdWWLA7t8+soDrLnM98wvJEzQ9PR3S4C/QFddOOPyoxezZ8FaNQd71LOl9Fq
SXPRYWOCl4IlQnBVS0b+W9CCx4pEKusOT/9p3FGww1NLON1nfIFIaDdnZc//TwMbsecCaAznQlte
V44m++vJ1ioRZIv2rMvxZzgIiTORAUrG1MS64KShLyUR42OywburffB4+xepxeCXAZX6lgk0tNcb
8OHzqH+Kx8DwnBS9YuAVwheV2qeHCJb4BD1GfkuFECiXKMucTexbjopecLeDGP/Nv27ueaYGBRP+
otRMKmrHz0P5FY7w1IHlb0IH5tqWQRs4q/8Vh4E8MdnaBl5zUgh/iN2Kgig1Nv0LDx6HE0z4Qij7
u5HFlAa9SOf9Lu5qva+CwrRbXqNuZ/JY491Z1m9oZNdG03JvqMhtdvvtukZZ+FlfuC9O72BjYmIz
L11Z6HDzWFOqjX1Tazxnukjgy+9oBNkD6E3hoe1NIC/w9ZVmU5uYin9eYJxb2LcQNTU5sLHdCKjf
EeJEajNxtgFL3XJxr5zmwtqe23gtzbbquZR5/tAx3wb4l5r41KSwGlzq1WoQ3vzzPkg0xPtpShK7
W6oM1j2SR94d02pedEtmjHIyAWCcgm9nJSJ9zfrzCFxum4d/BMFynCuoXLK7GZNlkTS+XRLw50mQ
clehX0DTdWNoT+92XgTxCxqU+7E6hOKiWylg6JrMtTLYnc8TDoQB7W9tj4UOQ/+pSDwrG3kMbqnA
8W5z4K9wSHAk16//3kNfxpXzBG90X4LdTnv/qNiOws80k1JREyK4oX/P3QXAg3oojLOJ0dBRJTm+
CFMTuK1fbNyz4s62q8t0tmFOqCgzP5Sf/N63Q1I3FAWzPURQyyHUBFZFAaHo0nz1bc0ANwZm0Mpl
08NLmA6DUq0US5B3hu8MXEIa9irtI3gDe6s8wKeLn23CjrCMfMoqo40Ji08dIpS+EEoq8jZIteS1
/W+F5oVsMFR93F++MkaDLjgYz1AD6T/+kOFsthy9FVgC2+iLyt4SBR5LepU8ER5H+Ts5Pc+yyoDD
U4tf3VTm1qHCVvwEy5e/ebm2LNp2nQ21/79rQ8bftYzBh3GHAUCBm9FAtAw8gjV9QjWZAU/alg48
shJVm6T3z/5cn4QSRWPODdh1MV89+FdHz+WPgGXMGx7f5w9U2lDs/BZWua84F707AgKwV9qL9Gkg
+1DkETad1AhsHeClhQtaZwR0RFcXaRYUWhpbAjMiRjFG01veg/0WDZ8ubYe+3wHSoOpXCK0j2CoS
B0Y/HNgikyLnXOaYUnKVTxoDx2Lh60wRiRowaPvjfgeZEcpOD441Tx9GvLztFe+VK/eICCLKntma
UnVHctHCw1VRFGTKexfON2F6C7THSfAKLBriRke4/vhivpgmSoNtJ0mMeJUi61n0c2fJOSAP8FaM
E4UPhyePmZ+27bFO8PjGxjPPA/6zzrdkp9RgXGxe9lxt6cbHLJPAvRfdG/XSrxrZuFqQ6mfpCwwR
kzrnmxYEnH24Q7SfTNNcpcElMocLLSTP5SjBShdxA2Dc8VcOIPWgDTInIghRnzqUyH31IffahgdN
hkIYv8GzC0kIPx5Aoqz9zTy6YihtW2RUKxr8YQG4iq3r1lFO6iQA+ad+kU8Jy3qX4ghLtiUk9K5b
y3JLMBLeFwwre4g1XzIxaUsz0jGG0k9eX0MaT1O3rInkkrT5dWhNMFzhdURXWM5I74gZO2YZpuKc
1A3mYrdJfa/tGUjnu/h2McDcrwRWevXNE8oLsARej59k6neUlEH7l5gHWu2Ww2bKKQdKr8GJjw7U
v525b1xN6WLJBRf7lT1aIsh6XR+HF31juEQW5TZvzPmXzSW7rfjgZ7f0g8kyrz1rbBbXxv1J4j4L
9vo27G+rnetkqM8IdSMMLUzq6qymEF7xgVV7vn8tOPxj66y+mmC2Nx1UY1Z82iM81FknckOVcsNW
kdMT0ilB9n+Qu2PSuF+nyESuTGtbX5eAIh3n1u39w6K80fdRDqB7IVy+Y7MFXtYoxUggxCCcU+Px
rd7jD9hb25X52MVodUV6/XDJz3q0cFFLAM5VkuY7x9xbNWo+kdnMIrGzzS3Efh1K2kKMMi7ZZsbo
ou4iGVy88oObgUjVJjqDhZjeUNWFZdXdhXH/uCIlRhbi96Ka2Zm1NFdpoydKWaf/5mCg1VHNAoL2
jtpVVf3p/sQpNz+njz4POPoqLNIR94qf4HgeKTp24r5tDWjQR/JWHJ1AecPQBw1O4wywOB9KL18s
zoFwUSq5p7JlUNWkOVTz6hRbV3qtKPxGMsJQ06nRLE40fKeitnEKqRA0WUakCM9zxUUG/wjo/8J0
9hdXHP61PKFJO2i0uNT90xppMzRW9PsSJ2MUIqMrZVT38CQ9H+wTK/AMk1nsDHcIY8t0SUTbeEf0
qVQHAkVSuHXmgSfQj/3bCoMPJwnyxDofjsOivKjZLKzcmYVDisHdfbJwwvc2Jj95OG/iJFdy5y5J
dKuQZt9OdVGlUEGOot6jxfUVuifW0vjbv35g/ifII4BtIhpOleneTL5tRN9O7EdWLbSDEF0C/1iy
4feQdCVqa0c43dcV28Me7hAkUvkTLo374JIFrvPpUO358Kv/G/KHJ2SzoTOT8mu7OKtO95GFoxNY
Mlwu7ppOTTjsQCZSIabTp0PAEcAQ0501FEu2xtGQQFADILvkcqn2roRaHdKVReeU7Tv3ee6TY5Ix
P4pkHowDZZPQspu3bUvEgSt3vOEif5f2YZb8ts/YFbrO6gyXCsHNFUuWBj3/B82UUZcEP4DMH0Ag
3Jemfipa7SzkB67Vq5dFQ8Fz/wCL7mdiH/DKxOuDpwuHIBGJZeVVE46naUo/ZopCggNgmlLkEYDH
R+lQVa4mqqE1qlLmxZVuV1aHmsN08/R5f0/cgZDSwzFkvHRPb/xyFNx+mnXBMPgbT1miz2iDzZ3C
M7IW57APFjS6eV7O5bI6wrYldlWy52C6h1A3JoIuwQZSNWGUAlmGGNBrdkcqabj6OQsIguyV30ze
maAneFmXKht1O4wXE7TaF2OT42PjrlrV6CJQ5XPTRpFQ3bJ3/5PRnaNk+5JTa4hyraHzHZoaJdxG
/U9VkWkC3sO+7xPzAMWBS2CgcCRB0QaBFNvAW8oAzvopEdh2dSKr6vbeAB5+SgDC3lFnwzuJYyX0
Xc30yufGHTdsXFB9pWLcEaY2t63bmv/+AWemE97xiqHxzZDclyDMu6y3oSkfDCseE+DQ7pr18ag9
QGHpSSMoEDp0q1fJ1gO9Mza09XeNnkItW96tJZp/771gmEFCubeP9wZqlWSAAbQTGr/Bt3KfbQgp
tFBycEh5MxqpFt2lvVIgEoDeAldc9A4Gl4n+bJA9lOqRMKhXlf80ezFpB0FzRCnEOzaR+N6wnBXT
6ci3+ANOJqiMlqtxt6rZ+FBQAJLieQ2gLzrFzvY8IUURc4bo051um2CNSWhMVAHFvDAHqpVjf5Pg
d/fTrpKQnSRDZ5jkTQTorDpHqDBbF/W6rHDotQ5iVVX0X2Di9FA/cfHBk6A1hOnFrUtArdRbvW0Q
PUQIxkvXC1PoNQGK/ZdvlbIO1o41H52f5QXcwK2VNGi4kein0sTgwuhmL6CkVnkPuZQcllrBoyD4
FiqXO0Pl1oc/Fdpe84GA6+H5joapPD2MkDoh51iDD3O5pV/4fGLOJOlQFh/yg3yYnLTAjyhBuPlQ
xtINMtXA/AkckRWD/NcvNdctwTfnRT5yMY5DrBFDp3uvuggBZT6UEhy59uA5D1woWCXojo0inwnm
m1fH0jgWQcQXcOGuwX4rESQzACgDn/vVf5jV2bwksUfJTrzwS6sKPDbESJtPrmlvcO/+UPn66Q6L
KHDVRree5xp2GCiTXjq8OsT/5nOmj3wO3huDjBbnl/MaOKZAZ5A4n6jZwvVLmaxuDFve2lUTQoSt
zgp/4BJ/IewnAug4GiTNVQJD3FgLNOLh87KsA9zgKZLEWh3FNSUIir6M715FCWdqctcF9gvEz/dy
QAcUjbqRW4Dvr7Y/BQO0cpSxzUs4gfXIA9N4uuWcceTkVvlEVF8TQZvUP3izdy4cux63f5GPqEIF
8Giu1CfpgHrGyyaTfQQEgJKcOUbv9hClS2Koj/GCeLisBcmmz9JdOf9TMrX3f1otPvVvwX1FUVjo
UJuLQFFa4SYbdLnbG5ZlFHgu8Dk3L+8LFEFVESt9yjgA2MP+aiACXUmcS0Qitz6yaOeJJ09XTCr4
QWxIvZJysRs/eMDDr7bCU5wxX9EuCnGR/by+7W/wGhZtlCauqgTrfOnFKx9yBkg93E4im0qV+MQ9
xMVEtOEg5gdxyYimNINreFe9OFfpIrMqIsxMPWGwHjdWGdjlwSEk09/JAv9GilOK0jZrCd/qbYm6
0VePUjgFdXi7UjBMDocPOOnwrQuNRGr2UNK8xkaP2QZefrXvNJ0ZFBPaIs2Qi3kw7D08rAyBuAck
ko6LZSxZ2N9p2raYndR2GSUUEUR3uLgEmNXEEoNE/DmXxZYE89jiDFaqk+itmQwte0y46VRD0e7W
ge7448+U0siAb72/VYgtXfjltdkYN4RieIsf+N8vyjbs9vifb0A86cWPPfuQP/ft6GNMQXXGHSzR
66YF6/+Zk1rhy3lb5R6QUXIfHXwKXCcHOWuoNPf2X9k2ub7bXJZ6w7gAf3kzIqpqTaZ+7Re+A8t+
IOlSDD5rMgIvW2+kVBjUuYr0Y15FZ2XPHLK50JD62txVOLHHtW+ocLpvK9Pvgai2hU7QuBwfv7UJ
0V2UON7/FyfLf6GQ2upPY9+Ck1R2aAYS1YOByiNv+9EpHpxCTRBaFVoL3hz3sP2PC3eChyrGL/NO
5+dLHqDQnkskA2IM34t9Gz3O9wvBLdobu5u1O06MWj9GEA7NzuW46laL4NYmI0Ao39Ywl6j5+1/u
9/EgprKinHERKAl7i8oGh8nLrp/ww95ASjvtnUYT/5PK9kMH8objMx9NA9SK4vAGzHm63lfZh9gN
Ywr3eERRpkEDpLfl3czCM4GiysOjEHfxqjc2zAhLDfZ821gJbeNvFDwa6bGfR+8NMYiUyZo4ViZj
RXG0V70rBm2EUBTo4/cEhDDyOpdQs4NUNH49Ly0NGcPHxG2/P6X5o3bvMrbrRUuRyphGhjN68WUT
GVsaJ4iaj/jRkxbU9G9mD1Ry3d9aKtwu0J7NJE9fGIMyGQPsVvOnakoGR2qBoCNOQATtTveKtT8q
7akaFbgAQnZv8uVI1n+CDBgXZKuDIHADQRRQ9PVQ9lJ6zXpDfQteFdO3mttsiN14VhJcGjIdjAty
oShfBjNGJ2JAJZNhhDP2nO01ZstDdfxu0dke1bZjwN1+rD4Cl9Ig/YTg+uHyhWKY2uKPv23E/fPi
7wWXb8Qgp5jBU15h+fCutElPs++tNEoCH4R1hgMMyn2Tu50CG4CPAJiU0GbPZ6NQZ8xk/31E6TBq
stItgWKghpS9moiP4IPaKmrTJXn0GmvD47ATXVgybfytkSl+rWxu9/LqWfoVWK4whg5TWZ1YUxNl
ZP5Qk+N2vYdzOajuy3/rB4lOS8R6AK1yGeAHySesA5faWyuMTcm9ow5aRHSPKj1gRyxtjmjzMKs0
++dtbFGy0RSVEUov6I2tluieMTXilhMOabTmn2WuL7lDrLUY4uXRMS9tqpanJNmcuyq2x/REXzj+
Nkls7Svi8lRXg/VKkAAwzGsA+6Fy1ZYn+uOWeDsJG8Jbzs525uKW9dZ7usDPMYL9yngXicvIFUJn
jlA0nsY6tGrsKftXeCBfiSns6ymOUW5NeLTdGL4n41GuOxBRKjbmbfeOjYp7A5RHr7gMLlYV7Bev
mGvf6erUgHcGHr0EL3yR0CwHYly0Bh66BZw60ZTczKyKCO/KqWFHVx3VF3OQfKNiDa4mOwwosHe/
umwDjQ3JXskwWvFGxqCHE/D95pO8Q1YlhGK3pWGlJzlsuo7OmsiEPL09oy4+RQ82CtKDW1rC0fBL
nZYdZXFKNBJvng6x+bPwgcvB+9Sy8qwenJQObeZrDqkLDiEERUeT2TAlLiWRmbSHiMbL+gLfa30e
ju0eBtCxkxvUsk4P3dwX4vEw8aFl5CCAc4gbBnQCTNtmQwmeop0hOSlo3sL3+ejD+ptpqeaCbM+5
J+reO1Cr/7vz770t0rNjL0tWl8IRn4wCxZpgqM01EWCX5yW8b7auEJkv/UrhjZ0VejZc+M0I0Zq7
sTTha+5f7tCPFOquQBUzxW/CouEpkoC9/UVjZ6l2x6R7HKgSOLkl7ScgrByu71gmuFi4r5YhwdD9
dUbOkjB3LoKJVLZkRu+ishVmKip8ewWIJlDPRQjBgfXM9KxTJmOkYgsjeuH1fCgKST2NunVa1hmy
2kwC4ofX47wDyx47R8LmQzWjnZrPd2Yk8TpMyuZzaxSJq9OTE6KYb1GcrQN/Y1wI+D2cTZpuFNp8
PKE8q6kDRfNXigbE/9R4UlGvyOIZFniLZiAlzR0CH8ut/INRC/YHU64WISfESSgOSxwzRBS8WTDi
EZL0iOUWBHa1KYCJQrFjNBxI6M0ZmfQaxZwLeoTILrf4WUJn5PwLPUcyBAWTiKIyJUkhJruVU/Wf
OTui2dpA5CH5LaW3NdYy6+rA2qfyVk25uaQGWKaCgOd3asgDwqT3cOcmhMbsgts0SvywIkzRwneL
EjexlhJiTErGq1e2wF2lF47LIiQNAYBPJ2eIY2jrQrtRDoE2eCN3LH+AYNO9rnpzXPa6UmldOUeM
nXsbXI9453EVBQSMY6KO436APGFAzXryXWP01aO1o8DYBx2Gf8Avlc9YQQLXAEPvEO8pYd26Pucd
v/yQdfb22omzstbF+55s+NqRtFwiZUEXT6kDdS902Z1sRX2ewOsHJFvhraKaxDUkvu7+tW3EJ7Na
0KZZmgYetYIFHQipm7u/AKKXrml0T9YWuWYqrMFZ6Pt4gpF04Ri0KbRSHFmzPYW5+13MF08JU9H1
0WvVFTeJTnCr0RPg825wvH3rTMjiYDltI0inxXjF7G6dybTj61WHHNzmMP9S2yhLg9gXqtsZvOGx
tjSTZyjDpoCOkFCTLP/hhNVRYJWOOpt/Fq2Rrd9V8Kod67olWL2ft0hHOBSaIUdd34yMVvN7xbU2
PuagsuAMoiLTSWJJXJ0pLep+JgaNcCzdfqHBKLmcYR6BILFEauZBc4h0fyDbtYIr3in4DFdXf/HQ
Jq06OZb+7R9f9dJnJJo/HKKR502pHI9tY12cUIU2Zur0nVUSFnuvl0QDbsR6nkVX451P59/t9rjL
ICTJtP8UONaFGrQM3D1vStJ2iE4Q7Z843gzsiSWByFKDnW4Us/60AxwESoktEy1JmZCVg/AQ3Iae
5Nw9I+lmciZtH37THgZhaJK3FlLjTELTQyXSXO9llF7cQZL20rBanEIAl+izawYJmG9MTEnL8t+r
mYhxYYhrhKpNG1lVpS0n8rtfjLpRNk4NPDB5OUk6CdynlQG/d+LLLI1KlGggql2wnyaeNNF75dKl
l1NJ3lH8YSZNc7g2kcSkbP8rbK+PhuYAMftTfy9l3nNdlEOzB9FBg5oUmyqKHso7YDGHAn2bnOCA
RI9LspWKpZmM5Re8OM0viXb26AdJfcmbHGiK+byXKG+V9ZN7+11YuyICf9wsr7yhsGW8aJq2fR58
izAh8IboBm3IuKSeLJWPVMyASMWOHMxYvVlxTHfDhq5WztiQ5MrPpWtQ6OCuU1pK/0cByZmStLu0
EDVTFLMRW3yPy8pc9dW9sqvghtggw/ywBt2nqwdk3qRFnah0YXd5cUxOEN8a86luqPxd4loGvV9d
bRla8M0bBsW/4wxnihxJRObHQTvvI7xmqCbqggo9fgBs6WVYGHlfNJtCfq/2AW/Fp57GEnjXh+V2
HWAOtln7AV0bW9wjljKzUhp65vPLvF51Fq05jbv+1jJKHm6zMRYnAuH6MaaD/7KnlNYSpWPfN3mb
1gRzBJbMLpJo7DYpp+ga6xpvZNvXXi6kqw4uhPRKPnyui2TikPyZq4wfrFkCajOmd2WniUwCfg47
asLfF46G2ZYGerYP55vwp2VJFZboPFxsSnEAVdKyXLedq98lZzr7MVFgNNY2lgTgIwAWUHE9aKCI
A8LkACaTK4FFFFJq4DYmBkemdCpeErMELZoKzEijx/N11ABRHwk3VagxYy0eo379JpGqWnBPY5Ba
1qwR5DhLt47lUlTq1cGUj9Es+kfVaaJN57M6ljk11VT4jSizcbwKbpWbE2H0oxGlPN0fRXANHw9S
1JGFysDNRyDtQqEoFotcnkR1aYiihg1K03dNJmSzo/YEP26/Yn5K5+Lu8+DcB80QYmdcQOkRiaZV
cMTom2x8fUgAzakSXH/5aorLdgKjiC1yWTYPz0RGfaH9bqekN0PJwmhi+pKwkJt0hJsidY9wLOnh
J7UQfJBGE03dwJdD98Sr6ucmYmeSTQp8wBS+ddTIo3M+ieEUGTbqAk7dX8/D81lE1vlZ05HaUhMe
0iJgAn/Tlkx0hn/DF1KrKYkyRljcWbDqpu1drg+p9HhowDAmA5pNjAJVpZx5D+oQcbcyE/aAmRGe
JICR5rbXKAeCBFwhQRwJhKBAkK+uK14hVSnFWmXgXwgDGkMrux+PYYHtUHXbgC8FynLZw3LN7JUx
DljRe+ISh4/F2QrdjBmJEivi9PE867eJJkRpNRIqPY9IkoqvmWNgenN/UrVHTvJE7bs1PBOVMhb9
/NbovXWMzxhp91Giz0hNO3bd3MG6f65/WUrP7/QbloDDZeP0RAwI2+elGct+EJBZlW1zFCf900ly
XZcyI306eOG1yl1lPVa8kZWnIBbalKqkf2/LQNvN43oZnofzIT/jF+22djGQCY+80aSXFMuLT8+A
FXRNrHNVoGBf6j6i91kQRQfMyZrcUBmb5auB2sHI1EHnS1vL1d0jRx17YtMe5UjVdkRAthjdQ1gw
LBTG/W05noi+rfx9aAfaGZpeOs1/OpZSfa9+HaBO+aR7S8C+RcFGjd4TdbIaiMZftPkRnB6uf0hu
EWR3s1DRxdk8k2rxlOuyzNRVIc7zJ14fKGkepYuPVP0GODcOYUfPHU2ES8rglo7JuQv3GxusKRWH
D0nCf8T0mcekPQ6SPRBKQARMi1Jaa/1Fbw9DlpAscFpSalAfo+vJBNwa0Y2JTag66wnWHmEq6kkl
mCHaHdIRNzQB5tfFxyLWh20nXybnxNmVZsTXB6doJAdU5Pj4L7hXCFWKhtp8UqfIqPmd4ZA0icw/
nQy+0t9PzSBNrHbiGRuChwWci9Lr7/xZ+o9IvMp/ftj9HlE6/x/2ACKQEMhCB00+CbcCkpZRdUR2
rypiY9mf8c7Vl1d2SbvRg8TmD5Q68DVbdXkVALr1BDyrhxBuwdivSABpUxD2ZtvxY3k3TTQbQDMv
ply+8xGUuqb7Hw1kjMUpxP3F7fttNwN83w3ACezPX1kU9b3Y/AL8pB7fyJKz/ybeNihr4/A91DSz
ZSrIyMyiRuZvOsrw5UMLoQ3opvv9rnFBa3TtAqOHL2//M3Sb8vu7CYQcI2VapYna21f7ULqxj/uu
nnl0pqbpBhP9zNqKFybe/kdkNAJYx5mnOY0TXi/1YrT4iHF/A9QT5bLugsQ6lh6kQAZFU7s3K2el
46KkdGu45puZXvlpnVHY57EP+8+gkxp0yrO/n0pGzTloeSexSbOQO3iO1KvF9UgiU7y2KWrO7hrb
6y6PG99fiZevTVzR/VoAYVV0MrT+F5msIjFDQIJ+yQUsCDyFWY4Y8T2suFyCMZqefiK2Obxxxbjq
nSeaNJDGmNnTy9b4TzMJqHFtwZmgpUGS5Ex2Vx9n1+eDMFxN28wJjOowHn0BKF1DhXVx2ROFdc06
M96Io2QE2oqmDPhpNp/GTALMAqjm35s37uk6hoY/kPvqBAD92TY5MjKaiZadntvvc9GButHSVcL0
fkwb5D8TYW5lvwf6lNaTALeDtA/oH1RJKO8rgKJjT2iaZuKjGTCkVwpc+WjgZ79k+b52I+M7eyJC
TTZ6FWx95Itx5IkVLYS/PBioT4igTxFUN5Kssf8vjHW+/A2vi2cgDSq/lb5H8aYlQ0RIuVTq4yy8
IPeJs+tEGS+JvGjfEJu+7T16VE0uuhoAYgDTQfC0ikd6fDEVDpiBPZNy2UXMzAR3aFFGG3Vl8lKJ
7eSEcAqgrdtpusi/ONhn8jBoqtM3ZLZvtz7eDs6ekPBoa49wl7AoeaTfa3UagqIPMBidGu4Fc71A
MIdQMQPtFbkGQHEmNQxxJBrwMY/ENUNNsACGDLlP5vcfw215RAVQF4tgMApM4lvEKR6+cnsDx0Hn
FTeYrr9FmLFgJfNbVAXLzYzI0Utl4AjHloD/amdGMi9GAfQ3m1Q4wLdyknbZHmlDJQolHmyGBe13
g0rwEi3uKUQd583x7TMtSjo89UOBxgJ5geWzzH4yMBdk61sk7ClDiSaxCoqfQ1qf+z6YaulLzRAO
FfJM3ftI0fdHCQ9Dyfxgm/XtlU7tP+79+X5rTOxVP3fNIZamCko5tPM2fpf+uzMOLHHNHeBcRWM8
COjZKU8UprSDjyzs8bF9jf12VCHIbT3vJlMPkQG65OiQpqNNaVayDzYVL/M6hOVfRzk8CG/Mcb3s
yZdCVCDckiL2iO4aIDAjM5Oet8zYQwsTbLN/zbTk8ryuyke4NejAVUFxMqxmyW+FROj24mX6AWnv
Sy3hto71pn4ixuCxZ9l+LJx8eEYBDxzrfpE/oXIWqZ+C/mExcpKkRYMSlha9ocneNu9RKQwDnPJM
/4PFMz43wT6Da/EqwpTNWzbtyqlUJcGlhku5n7DIo3hdxtga5LpBGhfoKw105b+NOs8NWm803+Le
cyHsZ+Hhdfcme/472u4z2SVHzvH5b0eaRFxSYpDPzRyPAmh9qXMr2OXYbJpl4WVG/zH+ThvPPKY6
ze0s1swTILmgo8AkbXQjI4s9HLirJJdkjh32sMpmXdMKQ/Vyh3KISYJbxaIHj7lXlqipssSbHkvr
pPcAEY5CXKl/UA1ZgBP4X3/054kHZoek1YSKuS5vRCO+jc1z23O1NJASaawXZRudvYTKIUecCCSO
JZzzmur9Rzs+cGqZISqQ7LYB0YIBOHl7jbs6YI6dLwyJFoZl/QhdLOK+GVV1CR243wx3rw0IrarG
mtKvOa4VR99ZWzJwbDETfyQe4ijb22tca2pDYUycD4Rr6pFs7gfYZYc9g+GSUDg127PQ6h3sD2yo
AMM/e9QYFMuNQOayVEZdE9beQjL4Uw9vh8VFAPxnjbMkZ4urY6gMeT02t762Nx9w7QyparqjDFDt
CYQcZa10BbPdW30U9jGI172VBMf0VZyhPUBuY6vUMQpRtU3tz0y5ENSJwHwp0hy6OxZRGszU/QB6
5RcY8jyY+4jVUw7QGJgOfN9l4AdxANM5p3DUEYY2XX97A+ZLeGtPiX0UDHGGQq/i1F/tns7kAk7m
MLvelMm8v55FVrNs+xDdOwvQj1wzIZ3LAXvueMolquKuATRQz/X76iWUo5Q1H2T1X4Bcr1LxcBxx
f6DAXy6w8PjDlWGqhoUhNh0w0t4nA2hz8Jj47Si/OHnh976Ok0/BKACyhug9jpy+ixyGyPNyqszk
htNv3hJtF+RaPq4GI+3ZjLsnSpsgLj+00+kNB/Uu4me+rVV8n/UfjP9FrqKMdKfRxhlWbDADn0yf
k+Es1u2bJ/IECfWf2x7463dFymWKO/R7cQc1SoDoda642VEtRwpTPJ/QWHuG8LopNKpFhpOVXQNJ
hAYNYtF5W5bK8/9YnIIP0qfDSp047jED/K2fzgzQcz1AhcOy/1XvnbXh2dg6q8EdgSULbNzgGrnz
03Y0o5osySTVrqjpzHPFentPzpdhtgozGTnNZkSDisTF4h0rRfiGOaLY3pJo01fR6ZoUvAX69Gt7
i9VyCKLo757AO389cg9Sur7iEr35KpHb2fDv0E/EgWxxVoj+3yQvIfaEfo1ookc6uTRbUt2DTdnX
wAAtDqL0WQUzus2TJGDIqA7T9iNmlTgmvEmrxkYVTJlIB9xUQGmc9qfB3s7tSysG6218bIt+WArn
lgOk43Uc6Fgl766Nvx6yt3BmLdjC3KMtxV3wFI0+33FV4IpG+NMyliBrRuGDs0L5x8PCEJd2+8BV
ocaC8mp5Me1YDAT+qvrqEiwLKvzYE/kqalmYJOD+byer9HtvZhnvbNhcXt1A8gc59c9/NLHWeJTG
DQAbUn1aJC2gByZFsMHrzn1BCOOkNAJPcWxtcgoiJO0f9ugC5dfryY5efyTZZouRqBeT7IE7mCfZ
JOMf10W9mql2GQEpDJ/c4MWa5AEvPT8PI7mG5awgpiMXx9I+jOebYOmB8MF7CjD6LegklTzPsmss
GfsRpVB9LT3ulzZRnMTltwKWaj3xsdl3t2bHz2a9uNfW5UuQCOl/wyUGHRS89qUFzTuOc887LFQ/
lU5Q1cpQVvPhwQPMZ/5OswLUvg7AO0WZdZG/LRYK98j0FovUbdK/yfJ4csTvYOlXbXSCE8/SlRUO
RNfHL4kUVf37kkox49+6JhPp8AuMqtT3TO2X5yjYA0iLD8wwyn3s+ymKi9Uy1HaAic3I+yuPCWD6
qwmgDab9dg3YB4PUzPAIFy2eaNdcRynJld03RKHXttpTch46ySzC0NCoM8rMOIYKk+W+b82AXRbn
PsstBTCK+u++h8CNuBtINiufAu2BnOPAfY7KSHKrlR+1OJismnjXZcZU2EdGhZbOU1A4JEL17sWw
Ngd7d3oQXcHnBU/fnuky2ieYhpk6X8CjVdW1IDmyaS5pf27eM4t5O8LxmITtxXzppxxuP1IghyZN
Plvu/oSiGmXQNvlgCBMUt9SU41GqLQu8vGx52ab7fV4nTRPOYr+WGtSrlPsTvVdiyXYTJwkkA2tk
LefuOC78z4WH1F6sisSjV9aek7ebKEx8t/6Z71y7o7L+ShyjriUXJPK2Rxdn7jYLW3e/85XL9ADs
XjMFN3XG13L3JAFHQ4h7ziYwsGhK++QsqpLXgeqf/H004c6IyhHMfi7dli/YqF1pA4eoJm42lTUc
M97VJTqNJ/piMc/TyoQAPzyJ8m/zQXge9tiEOF1OQauMlG/eEMYyHeengf6NcE+CoPFJMSNR12XW
jmaQX37JnDHB2dbezu2nf4JwroAi6vCecf9s0ujn9B7QrtTpnP/I9LKqnny6JVQCYlOac9Y9h+xD
2DBmFnSlIn4A4n5Ln7fWeAIad08+z8rLeIDzdjhDWehjqQMC5asMxE9Aqp2kmmNqQwxymqliPorU
Tzw9n52gTMZxFxsODHwWLsomXjrf3O89EOd39V3wep5YFBJNU1T4ESmV5w3USWpgqpf1pL2vp6oH
ZxBPky+im9t9mNSgkwDb3VZIYwoQLyB2mv1NYoXV247hBR12+sYZR8t1WQLL1XGzsEDPJT3H1YIz
DFnlyvLj9CNjNFnswYruEyL2H5Ca1KljDSUQMZPHUu3LgAS8bDbUTl0rj+0NGdCckzwt1k9tJ2Zr
vLkJCgdyPKPP1EDy7MnapIkrXPSjZaELTVQzvMY7tjxqHXkPyZYy8G5xLWR0rFYJ0/UAv12BoQY3
ctgeKsNI9CLGhTfY/hZ5Opy0O4OGOZbNI/sJy9GA1MyAcZIXK8ydoPeMLwRTtPPezd7fNCyU6oaZ
ecjm3cIW0syAf1qehCByiMEJgBGfk6HR6TsWrCpCQB8aXewriB/B44ziB6SZjAB3i/H4BbWJ6ALi
Mh3tnb8i5zseoEQ9yF1IDKAl3UPxWwLIdxj8Fej2sDTjOulgcfHanWDGyKDrL/v1UtIe7Oc53kH8
E3ELAIOjHlDsOvMc8PGtDWlLQEtVtmFeFqfk6eZbQE+6UjWN+CxRJMjt9dsp0xFZ0wye40ibBFSy
BooAjYZ9PmjZ5062CPF5tK0gSS3fKmz8XaduTzpbPYXHKer1pxVQboBGEhk+ZHorg6QwII9BrGTQ
yy0TY+O8bTqky4nt/CovsMFT9XfCcaiL5BNUjhnVareQBfUFnCGtcHTwD9aGVAIM1kbSkwPuGHzC
tEDlI5HMKLBNfY8m5S4O8bCAJ6Z1+KAYOpHge90qhEyh1TYeC/5pG1fqHy0oZCZFCOY8geXttxzR
19tBaOvUOGfHk6t1qOniqN5G2bP9BOClAuqu8j4VvVTVYMv9z3Rayya5I4pF0mIb6FuMI9DXWj31
1xB+AvUMm24kZXIMsJAUXZ6cE1SQosn2wmCx46VbpMgDNBAztj+i/Woq7ry0d00PNbLFqQiWy2/Q
p/mEjaAfhqn3hhBdTeLmIeSucwGqIrXOLcWGTHsF4Lzy2ew9tTqsOcMtRuXeAfO1EBsv08N6TzgW
2g10XKg0kN+4jNl6QahB0el+odcktRVe3YbwJmThSqtBSjU+v02mfY9b7S54KZZdYas6ippkAnec
+reS+EIdMuKg9PzjCYVVIXyqFnfAboBddFetUmMCW9toQBPpwX9lg+oeKErFhiJZa3xWMm3r+RCr
SXvNGGydJTnwGhTch93UKOFyfH7/L7Wrr07F0NTEh5XjpJXCyb0d2+VWnqiYzjrfXfY3UrxeZdro
pE5Wip5xH//vJWMij4OJLgD45X4tIMYMe925ShUOQy72L62POMzEGc2oa+YsOtjYsP+59j1IyTBV
gi85iew807eAUMWA7elLA4sKYy/DCFJO6sbBg65embsfVlRI+tpGB+3jqKgjf/gvNm8xYVcnBHZK
B5Bx2waDvWmL3/yVN51p2LQ1IqaRZYwpGLeJgy9sgVXUrDSZbsNVHqFTjM8JKs+pfRnlmfsSse5K
4pyU9X/t3v/XgoId2H/z3/gSKlGoRSnEUeFPUAQp6cCdXHbHZzuigsBPSI6AVQ0lELzrUy6WOeZf
YQ68bmXrJPNCKQcCi1DL7X5llNXEznktT0Vqu1Ji7TGIgGY3PlhJozOMBh/u0RQ+0/6Z71zKyjfn
l6j6C7y+NN7Ufg4H33l6q2rRv+g7JoKdTGdRfZOdqL4doapEz2DPGaQfj5xPiOzrbFpMqRekGLLo
H7bGA+OZ5dlCJVB88Po00gm1omdFeynWfarLRwsxZgFWVtB8P2t6+Gsd6pwGaE1DcvZGnJXZWyXA
N0mKj1xeJ6AVS4HGBmsBXQxL9VVAjBFW/IGOZQ+1fs2RPbo5ggTOEe5uXs3U53AMDLpBxandifUf
Z+aIKWlgp2OXNR7ni/IWnCpAOhzmvs7uEJPX9e/v4rKWpxaYLDFxjCOnUv2XHhonEazQM8o6fgvR
tH7ql8SqBqXoaOkrowZBAp1fme3oRqMCr6u9JJZHESdIPiBSCWdI1P9q0hjRkPY/8bL+d8XazkLJ
mi1A8Mryq/NHu/9hli2wRCWGrmf4Q6qwaEIy4G3hkZpa8ihcRhxEa+5U6oxsZL/GMmKhVjvIhT+x
8ZfXc43iQ+uEhwkhC37xDKlNhaCINSoTbK4qwub8BG6/OgrsKnb2w9LYsIVNlJlFxNvJl3qkqVl7
EGjXutUkyBnrx8J8QES34GHtcYjQtkGQ4YjQZ98WogTayWBbq+3P6zsw5ibjR8LH9AQPpr0ZfeiV
G9dfovpXek9x+hCQ3TKQiQNufm7IXm8rmCjzVFQd5Os8KffQiurnb1CE6V1GLnCxbToN+6vUKERV
8fGLxSyLENQi4dZpj1CwRcyIPtuHw7SnX/z/HNhc0dsTJqY4b65Yluk0JcJMSMJkWJwxTllh4IA1
JcmqWViJL3BZynbUUfmcO0F0gjjkRTC0xclpQ4z8Wv2rQpUXkAKUuka/7eL8ffUDJtp7Zaa8oL0b
KFt4Qe0cmRgD7ktb1QCMAT2bSoiOOXBwLspLEHDpip/llJw1YtOEeVTpzrov7btVLxEdwQr55TbL
5U06HcDqDVJvEvLPV5UQZ1P5ZDMy9a5Mb+fCdLSa5ZQrGuoReGFAsmUPOVtQF2T05yLJru26Rsul
ApjKvdaGPt5leXHnkaxmQKGy9TyHG8rw/+qxpDQTxdyZ4vLnnRQkgAod7BlKTbf8arpcWJ/Oqn3j
r/ccdp9JTZBGJfyZqmdIzsoNyHOSsk0T5tLm8Sd0Pcb5IzuxOBkszMXF3qEgV3aRRgA1prS5G+WG
4fPtnpI7OLuXqFpLAV/ipXi9prAkSjB202Qb0QcvFc392rg6PCqAitc2rugWTH+7zUbGwE5aB4NB
9c65Tx43X6AYfwcMmwqo+M6nswlR290++EweHKk+qXgimJvsVdsO+g56GzA9JgBb7MXqT/4zQXrR
jeTjXGz8SLlx4hBDdsHWpvKBTJ6FoTWmKJw6jZsbLBofqgKjYnitk6owoIdJY4ddQE/K29DqBHz1
FGAQCX7vJ5kbCrHJ8NzJE0cYOcTsl4Dd3T26bEafO9stslQoJd48kOUpf0gfIIatxuinb+abqXlT
o4kGQcQdTeM12bYI/GGPT+9f3UboSmaOd+MHiONjd8vwvTGwCsHdPIV96/lcOd5H2caI/9H6CAnY
CAEe/nEw3AvrcADhtjJEjQWsC8R7P25NF32JnDPL5n9s5GRDas34NWjy7fffqZnfpvL8EggSq/4b
pZ/QHizPBasitz8YR+WysIAqL9VYY5okbaKwSSNWhxYcLzSfPa7zFsUl9c8o446mhbSTe21s70bX
EqeKyTdsT9A4ExjvgmoBbJn+8aDOhYvf6GysWryLmksubfd2Z5np13MIiPfhEQXAdCBDvYAZT15n
ExkFnmvUwLcrrifLzKPPOgiyw/W4KKCyuHKJi2p+v1ysC3hhqwS+yIIiMyAarBO32qeqqPkjfIZV
OLulU9EGXdIVpPEdyec0QkYpzG7c3E9KthaTq8SE0dkvmWlgMuzkXAxLpnl3rVNalGo0HhMSgdWo
a6pXGU7cljsLnF50DsIVO5DjeShf6A5A7S4cQTM7A/dv2jHtIy9hQRRRIWa7NK/0ELEWvGtX04Oi
YXF5UzZTrSXyEkC3zF8vSvXSabND7wx++wLCaQB1kJf27cwRBBIX0d3dzcmnKlDvCSdtzvlGWFnS
WsNHIpFJItQZnxVnDMHKLLVIIrn28OeIOWV3fuuE3WJXMxAdc+rPX0q6ZMG1oNIupVrddFn2xIXn
dmZYBbcxx5wh3pbVHqeKN9NSKpxO3OG2Rbs+TEeEhroECgtYMGmVIsTq2tLMMdU1Ve+Z5t5at8TU
YWlYfu8S8jsWFM28jmNTgj4N4CQapuc3k/AtBGpQvCVQLCmOB+LwhAi2InzxA3frAPwcCF8yZLdn
HeS6weWncezFeNC1GjP1ciIHQqtdGGGAvzx+M75DlJ1hu37ot9oT5q8xPfCinisS7uNVK1KfmyBo
S0smzlCW4/LFqlUP/VomiIDXUIuzjpiBZZgs5QxDL7zow3sCPEN2mB0OsxbcM/TouJsdg9ywieAk
wSuB//7fAxXQUJEuNFCv1ID54Vbf4hcOuAzLJd97TLspXomQgM36oVp7YlOmgPTZefgzPKtGpMwB
KLo8K9ng0tReRVtPOQKolaLAFyMQyleQFhuwMIAw+YavH/fTsx/QuGIIkB93Y+KKwKwzxE1nsMsi
ZZcsY/bCGpNmqQp9T5V1cSoEYmdSg6eJr8MTj7kLstOiZep0jvoiEhPrBuLjCEue6Tx46AQ1ZfL3
oes37UYhZme0LLPM5pYmNi7mSrsNtB57cg+Q2FtSLc9wj4KgeazD4naAs2Zm60NmLMqnqn1gQwT9
z7OCHcuUTI2yHiuLAJFRv9TU5Ltn2IBX8Ws+BAtioFE8IkPY4wgnwyFpZ2jgcHLscNH4av/5/ChD
VpJaWWGmp/Te9p0Fvy5cNZsX5AxRIFEsqYZE0xB70PuXuPrtmkMqo0dZbRK9XdTuMVijJyk0jTrX
SaLBG7HUn41aG4FHxMyvlntIEWlHPSnBlYHLe44noPJY7P684j/j6I6wKDyp1rvqi4CWhPJPzaZg
RyYkQMSJZRXNGjbsVT6zf8UwQBa82i/b57nJYyD0UYvL2w+CUs9G/mNaBLr1fiJhvFMDUr0NyFfs
JpadlTZofjcW7dN8MGK5qbA0+D6+NXhpEfchMy00pgpCzbx5iuk/DnSjl8sNTO51cLj2PP7IO9px
pdmfkvGP8FtL9CLghCRAEvgvTitSvfkR0xIDvS8aBAPe1lP83paCBxiMmM+PvO67obflpUaQLtD5
qGYdTaeE0d5DmQIDa4ocSpMqT+zeE3FZzJ9SQbjxWuIBYV2gKgTbbF0RSIS3gg3EZT7Y9nXLBu2Y
rhPkFF/kAs7idTsMuWBBNdiP/yWKzTNzfxaXcrnXIyqtvIwwLJFZ1jXy2+HN2FOdGHRzS6Y5TzSd
HYXh51OYvwMQME0ZQ4a+QVcNFxOdnt4AH2i4X1OVc9rgW+Oq5j/+w0oueGr2UGVWVYKo3NIMs7Yw
frH4KGzZSzssjgrY6X+hiFLSzIVdECs76hmqS0tUL5WZUuJ31uMjuVnVb9nawPJLsrV0uwgnChvS
MaWx4y/zMjNX14UgBJLEtZjQXGUlkaj7zy349ALbX3ATj3aEsGUtxtzAMIEDkmGCUZGpd4YP7Otp
mIJ1V6j5/uR23zNSny5oowXGVog3GxlkPs951UxBQPYNnUQoxObXFzG8GOhT6tO767sPxOwHcwKl
r6NazkyQVTr8tVq5LNI4/k3porSdAlSBYFk8BNWCxGI303lEkBMquyWpAfYVV/HWmDGCKc8YW9ZR
+ZvPatY0pSlVU/+6uZBgM15FtE+F2RV2EuEQgPfYG9kub6iijFhBGbVfqo3EP8A1ejmeTW6Yy7Qs
ionMr/UGHv11NnnijYOMEfw8XgOFsgIVeAX3ntLMW1xYma3zNb3fFoeApoFE7150m2Q3vMwg7sI+
Tqq/iEGw28T0RPHxnr1zrx5oyyhDGRhYuhw8Fv1i/U/T4zCzMadC2mHsu1Ep91ZiYoy0Rv0huq7Y
Af+xK43OpA6KrhrMXWl817Cj9/F57h8P7EoD7Dxyhg/OvXHjWko8x5UFailYJ8Z6WWmfo5PXVaga
zUbFhYuhmD+qtqk4rDq5Ugyeer30PwG+L7qE+BP0HqZ5eC1JMC7Q01IwjJcM9wafa+mTWCxoGsgK
KAX6bSMmvT89lXD4UMpYtJZmK/07opraxBMmTnq+3feTB6LGSCBWdr1N0JXN8HXfMrtUyJaCI4Mz
+7Hezyw4M/FS+L7dfsCNxLGwf/kCd1E8j9+xaxGAD/HYNvgaVKGb3MRS0jLUmGEI7OJ1uDSro4af
VLIbUHt6WkVS9vL89IgHLXWlYo8DSYLWe/lhCS7rKdk5WOa8iU6Cv5CLVcM3SBXFwypMNmoPlCX9
BH76xExnuaO0GRGakZgQgIci0NNeOY8aL3c92QOA8KDjJHXmIY0/HALCwqior32sYbSkxIeZzP/m
XjUjQzBvfdVqOzkCR0HYid6ghLiIdTbsr4+sTkqdlQUiKn0yL4klFV9dDTcRHy0bL4WGHeb13SHd
Cc41MlgldBJ29TQoRAXiPR2fvw5HlscVNBu5TwnTUC4J4Ak+tjOg8vwPQBYFDmGfPfriF16mAECs
h0rPsT2GTsng2wHg+MRJlQpHD6L2JCDszft8mNgWrRbQyFGG9/AP7fOVIANGi9DF0sZBOvXVH7TT
/NSwvkpBFgvXdZYg6nvKg9gM3u+E/sjozKae5Zns6aoX5Yt9VW6O+Mx0G2DuOMltE+pyc2o44dsV
ENe5TBg3xZecp9FalmO0OPYZQBJ5pZzkYvic7Ahp8mdKIO8WT/vR6Vaq6IgkOVJcP32gsP2HvrQi
FegdN3gQ93wicYlch5bP5tbJPqHK9TYKuV7wxXGI0An4DkgYiWXhnRW0VnalSI/4JdsV82ZRkBjv
IqqrUtvbVvV7TcT0qAem/3SKGbT39wUwXeVvIZL9FRb3JnnEr2+YmL0NEwjamv9MuVAMGBJekbwp
cPZkW+Vv+8pdubSmCfowhNv1SM9ZwRafarPthEKo4xuIk3OCPEofoJgMjNxU9j5C2m7+SAwu9whQ
wxG33/IOwEOl9QMFj1HlVFsN/5YLMTXGkONc+su3i+QnHr0eZ0nGGPtL1HBVDAMefLHtm+/j3Gfi
1+iCHBoWdjF1WUhChV8Ua2xZ6l4tMqqXIQahzpWmCSlAT0L9A5Nu1xDG/3Uq+mJo3qhGad7BAzgH
arb3aJA0ypoTfePmtw8VqZZj82ok6POXkzn0QD8mNP8ys05qwZNdGnFWzbqDQNiMuADd84zG1iLt
e5ZZ86naSSiMI/17EXwshpivbe/CBgaQdy8RWBeS99WMxrdUit+4928qmo6A8LPNRu/M9WD/uexZ
EG2Hoe6JaNNS+ZuiOmfe1gh4CpbYuszv0zUiwFawcywvwx2UNXFbxRn6Kr/fbGTKse+/wjgLayJk
GPA1ofqF4iaLNDQbi+Jqbx7Py3PoG5EsgUFq2cN2X2jtYTHj9qSz2IMT3/7u30scma//UY/b4q/Z
yEjMnCgutaFLpcNAWGhsgOITerqPYwgSqN6kB0L2ajowbXZIssS51RIMYjY6hzYd7ZveL4x2VUt+
eFn41dgCzmdhXsm/h1pNi2U/VgUhkkTDTxJMmUUhqShKTN3jp6yQV0xf0zujXisuiIpEsMibyhvS
pZEa3kbemCXhW3DvZoEP0gvHeJ5ZB/9QhWHsJBN2Ikat5PeVrxvtZVUieQTMvHOUXkSVoqKHmR+l
mVZBPAIZZ1ofKlrlWtlDTR+Jkfj0t4HzmcrDWu972CFKF5rcjnzKxa8k9drRr/n+5sRxPCl+4EsW
cIIIxyKFMg6fSI445qHj5Ga2NoLK5FUm2Ufn/3jHDY78Q/2Zsim4iRr+1uItYyFTPfthrIjencGy
cE8C7+gPaL0EPMxrepmPevk0sR+Krzt4+XxoLhMFK6krqvYWBFqjRafw8e65Qq6Kiien1s/N3igi
oGmjqyK3v1oGebfWQPhqcOYrXkOwefJt2s/9dU3sDztNlznyK93daiZGFwtNTSVCZheEIGozOoUW
isWjAl9T7XW72F4z5G48diR4JWTYeicLOEn4Wn8y3eLzMkL0nnlFZ4J7y4Pp1gd3fSCqvg0dMi5l
6uC+nEOQmrFdqN7J/qAQ6ncIR9+JRtocthKYY9ix9ncOd1cQXdZsyKyIVvRZaVPwJ4Pqq7mQegSt
hXP3ilnhgy42bMloHMcQ673fDdJVAOG/P+HSOmouM4e9J7LCiayDaQgKH08A8wPlhXGlsYsEiUVM
lchi5iulZ2gkl6bI1YNXAmu9Pwrh17M89WKETa/joCBkck3sSeXBaa74OGnOICbMpgHkuGP9PLxG
GWKvv2V+B1TqpwUfQX07ht38NxpUDtyYyEhlhWMekKTiHIZMm2n2cdX4ySv1IpRxvhbPBXNZBxkh
ST9/ZOiie5cXJWVks0wiEsbLx40UW2KVhEh8Y0ScSoM3X8AezkqNt1e7QT6zBn2/p7abaoCcf6do
mhXftOG+/AoUGKj8+5noSfdK9H6PCDtTaFmSaVI41+VJz4eS594N2WLqGE9+8LiT+XJILB4bvxEW
wKIe0uz8Y5TE1MAbvBNTt3js8Goo2OcViHJQuMP/gAhgR6LCU2EKix1F+xPBI+U41DUsuUZ4LzBL
fHyJTEapXP9wDUL8DIh2KiTZM/0wTWzoBnVf6VjHZrEYT66nn4htizMwLgZdb9SFLAwnrsBrYqaG
v1KOvUTf6PzntTeu8pF6OiTaHr1sXOh1q3F2GN+CDEHFN1SVGvLnN2hjVH29dbCYoXQrla7l55ik
3OQNtLiM9xEqAcOdAOoGvLRTkqKnWu+1Ky3nX2RKGa7RxFLhKNX8NiZDMmAzSVxIAQktboRmhUjr
1njujYx0n3kAdsh6HRqU+3mCwYU7yPNtrfVoX5W0T31+DS25RVkzjdupWgKESkMp2gJCWtgIFRD4
sdcB69X2xF/KkhoX+snzog9UPSTpWs3br2ne4wVPMP6Koq01Twf+KTSwhfGh4NjcUHkfDjXsShlW
sBhp19rfYgcKhnrOprNVIKpSG4VvPFHWxyAzwlqqGKbbhmBQgEkL5CqTuQiODx/vx4zUiPACdhx1
jfZtxZriVUuDzn1NOhAuo13CxVC/cAfEAe4DLGbLY4iPoHfevxImElSQ9CGcdd9KxJFykGuU2SFF
TsB9jUMeGFP3b40owZK20GgC/duEl+/mXgwjG2IrVjQ80zM2dqcsZfK1do0i6iWPMHIDah1dlVMV
0EwYKOAvdl/zB9ndJKMGd1Pm5ye0cV3sjtHCzMKcS1feEo1T6SDomCHfDLtmJtshpPIbc3ru0nqK
7dqqJ/FDnSKQwJ7HJ34Wki+l+NiPNmQdN9Y21ejEK2CCtqqN/tc0OYWSJOKwnYeS9M8agvr1g6Lk
PEAUnXEP8ki3ATupp2fGvfbXrKO2QrsBmA0jhZxDyBorfI93okEmhVfpCxOTLYP3eRKUzc9a3dmP
4QtRznZVnXUIyocWGRPqjwFwIrEkKaTjWSK858ufvljCE4iTLuS04nwv3JcnRlPbmh3Ct1bxGTjd
eW/t9z0oLrxxc77MhuYd9YvOLvi0MMdh5Njq9KG1E487dzbmGv6Y+fs6PDvUbpFe04jpbOADFT9p
Z9R+8gl3s0TKOa0fbtp4BwfpPSu0+WNg6LjtBpp5HsltjjOoE0inYWqLkiziyCp5moIJzRrm0kF/
vG6CVTUN5l5YNQ2tLBM4gHXLfI0SZcIWHP+0ty3WwmQfUwn0PzsQJ6Ct37Yd0ECO/b764OHMHDsB
CcvVLFeP1b5mtUZpLEWYDOqnYptqxbX6thlpYGBSdtoX1hldA1mJP9M0KbbiWCjgg3fFNIC5X/SN
ASYwLRQ5UxdRjZiQ+NBlWPkMF8qke7AoKqozxyrTV52rM1kVY9OxgimEYmKc0FXn8tQeXhQoOvfa
YrdQfIg+4t7XOaI1FVK8xnwM1KWrqMdLLjEVHiNJ9fcrcXeyMALIwasabz5lzPJtwuuo/JVeMxeR
5o1req3vCCGehhVz5QGL3UnXnR/va4/fSz/UFaNUHU1MORV+LN1BiqD0QqZv/8Ghpd/p6uQiM9gt
8l4VsY8YSFZHAA8zP12JTg2/HiktgrR/OdrIOLe2UR8L2IhR/W0JAxV2MY26HBlgA5GRC/8kvd3a
E21iWpn0laIUJjvo8iTG+Ms4WlvZomHykjP7sEZJiqmqg/qv6NEvGZcjGlgqeuZXBdnl3S1YIPUi
5ZsIeRJjkTXAeIxKUeghKWc50OiQ6cU80crpEys9QxkKHHNpfSFbH3esY0uNEewP50+GEYpTbod3
DuttY14Hzh1XaufLrATM1Cfo4yta0pbo+n8msDa22Xk6jLkh71ek7oeJApA+qRuI7ljEJaS/r0yE
oXffi+x+3Nz+/u/f4VqWUYi0ipBD3arbxg/s9cwXx1YVHlW/Y18Ufet6xogCxtDbytPFwpr7YH5A
euhcV4y+ozRuY4rn/nr6Jf/urQZewoIFPF7rbxRv8OUm3cOYmam/rkCSz1sDYAcwJBPM5J6Y3eGn
gOw/22ZfX3kT+3f5RWslYxn7+q9g6QxvL0j8gvVaSxDFCxLIQm6txvbDyGItBP072FYq3LUA8zgK
z1W5ZAjf5bV1NufeVHLEZxtNcqHm97JT0A5GwR/bNY6R7fSHdkfaM1uAWCmULZkJ3Q/iWNCZ4fQy
mVPUhWkeQT9Pv7FsGjpj8dneWvuhsC5ULycr5UAT0FEG7TY3MUxf4j3jRI3L04TGMCin+ueoHZez
Pfe3YJckqzgcbBE+WB23lBdyGf+P5rG9RCoboAthqpizRsoHL3h1I2vhnxEa/9U+dNQ5mzUFU9lI
CL/aL2u3OC90sQgLNs/BwpSUHaYPUvc2zR35h7CfCbyOfvO76viA3BLYOmWwnGKXYuCEj2HrGPsE
7wZUVk1Lhv5hzcfMv8WGV4KDdKIngnpwygy7cxRWBYVKIVdoXoyhoxuLfzVFKim95KXYFCxBrYu2
JYsnOxEichgg4OeaXlZ5Wkr0uJgcK8jHoDdeX45ADvsnpK7dGQK7oTj+GR1q16aWLSD/8HUpylAS
nN/4cKg2o20cMcx0jTA03B7eg3SU4QPII3+uvm9mfCSS2iZ934PJWVEb51/Podbp/Nvd88wg5hac
GMXseS9MUXk+gIE/QqzY6VTvbwaFIicFIOkIe7+sMkwhiE4Mv/ZMzAkNd1CW1k3JJHs03pOCoOrc
Ln0aNHCbZJoKSDCG9HBhH7gFVE89udlOuMsIMqIdYtnDjZGBvLCuRYyzdqTlsVE/kerwn7AizKWV
i3mESA04ddgvegCF1bpLJvMTpLXnhNn81C0WAtWhnLpicNMNaGGZf1rzYyapjn2/k/1yv9XiWc/8
CiU2KWNKAxWx+ctezgceklFZSJi4T1GeCoks08SIlvgnp06sDEeF6soNr6fKMm9IcRkLKpcGoYlP
72r/FLlcy17Xk9aiY5Srx8idDe2etSDO7tZY1h9yLSAnkSDdNcqQ0nZBnVylECXK5YTWAkOwKkzF
xCNjybR0S/kWND3Q7dX1MOHf6xQS5cH+lc2/N2hVdlqI7c3JlJecoxOrMfS1WG3oG6ZP/ZGbTk3K
fy28fzX2Qyl7WZ1T9xuOehFp4d3iS15+Lod5S66AuvR7pbQJyM1Su3mmIJbeE+b1pYJz0GfTvBAh
8e1EfmjDB2N/xd6V8egHastpWsPJfp1WtQXy2Zcepiblfj+KPJMiR1T/mwRJsS19+N9P2CnHqPzz
DHTFlNsVTnxuhl7LWuuGr7WI5Zot5IYUQkP2HshYDR+8qVuGyBkqxwFA93cdcKfka17BH0ZKUWlo
aUYp+QJPChe/QsF/Or/2siNHPq1YGyE8ORZJ7S5eHxvF+38cDRMMb6KxcXImRFZBmr1jl45NUoJM
AxYaJTfkRJZK4wz0pmbJAU8FgRMFz8RI2F3f2QHrtSfKriowisbZ7WUE9eOFDLUYji1LXlYe9ag5
zJaRGTKm7ccEpXqTkNxDoaSZI0izR0Ad38WP8B2hZFdiJwDHYZOZUr8fgXheTVxpFe7uXy31qSd1
wAa3Qdj/176n5C1lKukCtfF9yB7UNBiA0n9QpwuEZ8Xcoe2SUE4IblciVezR2ogRlh6NrrvC83fH
kpmds7P5rGVSyt03Z+3/0+Vs+KU/q2wu0SEwKdd4kNJhxBT4ptAF93MA0TDSIH+5jBK1wfmzpSKF
5UOy5cLPjhJH+3vFrIazYmtiUh6pfTAwF24tMatqn5gaEZxH1C/oxodrBvWOQv6WsEMAQxFh+L6q
C2abFWBw/gzRaBCgVfkqELixHhD/+mLIveHY9H80eXJQiVgm1S1NfLrgLS4vG6TFeqw5li4Bsa5I
vLTUFKitDzXxmTGgLNv+dmd2AWCIOjmKKjHIowmfXExzW7lP+qfYm6tl1rCKTx9b/BTdD6mndnM1
zmdIWlEXwKAqzj9Q+jZDk+fexQY/gFEIPlqMNmfyZusmRI0iMTSw6qQ8GG91kdRMupeYoM48qyDJ
pmL8skwRIJiO5KidAFeZAEkPpQoa8oLaL99oroDsQ1xoXNqAnr/ibAxUkwCpJVeyvDNJl3pCtYuI
HxtEzNg2UTIe/iHpDjH3Nle1Gkmk1oET1oFHQDrdLrth1T/Hya95Qh3FwHFjvq5H6OZRdXiOcimz
rpeUYRvLsWhLgkSVhislUvTPrxbfp6zTw/d5J8oJdzLkts74PU/Dsw8ikjgEx0ZTHQCYYCHEfRte
liDbfz/ajKCDnwg1oXdZA3AsBUY5fe+3+o2/6pmunRW46x5gWn1lS2zb2nZ0CCjzIKg/Qf3fi3sM
MzQZdEwHukMT969eKsgsQsB+XV4MkJQdFfxHxNgjgOriYUp8u3X+KD6hLtxArfCvkF16RODZ6Elk
ITfJbpTTNMHfGstDwVPd3tWy6i9/sCFhKHB7HPOCiw2BiUvnTbO8XJj7hWJHKma2rpm8t93MU1sz
bqBkpDeX8a/2ZafZ7LCnkvTKMLBMcBWaU9FgFCZrEgBtvYMfmZ/avTPFxJys/D7t6OcdbsXN2xcv
tCEKjkIQjjg7LHkRout84GgYzcS2dHsatVDXksUhYDOnvOtJqvg+ObkJ1/RgQAD+iucO9qmLtawD
7mzeG2CXl7N6bDacuslhVq3ARKcBIL+B1QKwTKXEY9EwUZYNYaMH8fmd/IcGWk0vKAOdtKkKDrr2
MK3aoIgnKVaJ69xhcK5iT8qWOxcl/oT+GbHAw6Nkow6cSIsMDCvU/mCXILXzcLPtrf9Xuc40un6H
V7GiX/JhGGLA5iH4MVT6FWm+sZZgznX60RHpSDh0Hvp0GW464qhEHZ9dpEjBS/jw4zTv/0/ZXML2
gxYljt5e636XcCT4ZwBydP+cMfEPrpI6TMgP0UXBpVygi8sEJ5SZmOBQuzMAPC4XOl6BSkSsbI2K
bRU812XdARvct0IUrYee+F9kDQunhAjYxH7955C5ZPLwhhjAV6ZsTZ1db9p27BPsd0joBDWPWr47
4n23BPEQghhnDo1NJdVlOgxdpQpiKSjdF05L7AH+1d1FZdnWWNjgMf/DCFh8+G4B0mLvKF34yb98
Y8xTb96aSnU7N/g8mASJJFG0I0UoJ/p54qaSDmjVbK9ohNJTSRNue/v428tKAiAHiWBNhhISWfEP
X20FEFgayegssHvktDnMYGCMiJ2WbU5SFyVRpLtDOOshfNOByMXUrFZnzZv6KMMaAPNkeiOcLTF+
Kp2YTembee4uoj5quWWocJPpQ5eeimT1BHEOLu7b6rNfNdzIsOiTmQQeHETy7LZogjrtGQ0q1Ijd
BFmePfc9JtAYMg9VYfhmTEeSS7tjDGW9lxKIfbNZ4xReokUpHnmyfq1NY+33LCVtcFHPx5+Q3ZtU
l/lpbKL2L/9511jd2fqt5uIhHwS8nG2WXRvSCy25xQuyH24BPqynIUn85bapiBwEKcWlgmdPJJo1
es5wwFWiwAR8/o+DWzM8V5xyJUL+cIs/N/IlmDS4+qyNzGFlYs8RN3a22H1oFScC3ij5GNATKlXX
UHeOd8Ja5AYR0fOb/PcO6DaPLZh5mZD711ZiqqFk++QO+e0fJ2NHLR3jBTKEEcn9RVLYc/6NTPBR
6F8NCoKOND2lEE+X+nCr00pFW5fQjrfDb9guq5hZccXVJVwLVhFyNRBqzZsK6DhGcR5qRJnHNBUg
g5CN16dL4h1WxAECHOZLMrTZVFm9Mmn/czkPW/jcAHE2GMMKTcwWuhbOOIDAZa5OUJRP6oqWr2rE
z04H2g2T51Jg2Zy/mVQUB+C6JSVPwEXjwMDMA7uSk2DLB5bCTqmG1n9LIO99KP7OMpJeyUC/WElE
DxAIt5EhZT7/k6oT5zxKLVwnmvkx9b/ha44QH9U2tX4DzkzUmauP7mKf9y+wlFohdbQ/nQuonF3K
TiQiHoaJeRCwsIcNV2cg94CtAKG52FTFHEnsPGLmSbzMvtwfqsvPZLscPapOKALtZWVAnifKzVBc
Aol0i8PxKJgO78PGMp6H1unl+B7PLPOm6iAVPxrtGHoD5p736Mn8A3z6xk/UO94FgNFSi5pQZSSG
lbWvT4xX6sJwTEdrcZhACQBOhNV0JFzm6DAdQ51KudEJp34Kwrd05HEP6QMR1xL12zxw00deR62O
dEqUTKvLEdLUmT81NgmAGRmkL2orcZbWuExRU2E/6bDlvV2xOYVVLwxBAFtIJMhjHs7YbFsS0+4Z
ALGOo8sp/OapBpsHVB+rWg+ZN7hMw6nCK+FJB+0ecWO6Z0nsyUwoBuC0fFpPpVULjvj36uMuqEvw
gV1d3UC+ply2CWvWe+Dn6rYJf1l2DtGZgosJwuP7TRL01ER9X9RjO5Su5LlZxIUMncwfwXvVTWbc
njcSyqRsgjdQvf/P9R9mLAmVU+LiQzBNqEUyL5YhOWX0qYCVrcUBbRXXxIkQTQYlfeEYYugR7rGc
FlDzBhVq442YFHnKm+lbV+NkxlJPfNr/xWj2PC+NnAzh3CL6Kta2WXGHqJx7EOZz96fq12A+8SbX
EEB6WMD7e3uNMWtHjNJrbWRslhRLz2jaty9eJSFISZP5FwqiURjwutb0QSKJsO4KuZdvrIFUms7p
LrjR+XnWI4JFtzcuc5uEZrWHUMSSfHkAzDyFbeewqWGd+Z996bKRUm3QwMr/EDNoMJBxF5qJOXQy
3tLjBfpWZhB23Cu6WkvomxvXHdyx8YBLS28sTMYtsbKOIJOAMcrL2WcR2bR8j/OuS4nIqwEdNRBe
8GEVTfa1O9SE3+m6jPP1rY/WIbe3/y2AF/wxGFB61LQykm9ae291+SZjvQ2bsKca035whn/VfiVb
k4zoS0tWJVEQs4kCx1VNHAUVe2NVZuIuwhimLNxaN7xeRNw4SmD4QxIFtA9i1/7mQ5tDm2SbQaq7
LLB8TMA5ZGIqWNhf1TXK6fX9QoFskv1soNvLRCC4swe+plwnw2efqgp/3VAlof1j8rmugmKv2FTG
if2mDR2ddqYXYO96upyeDGWSyP9bW9rukUysnKm15BgUlopz/Mr0YE5AURSkRrEaO7i2gWH0n64L
IobhWTgnkoPNd/eyRM/99onFYhkWV15/g7918QbeLUht9GkxkSr/ihcPqA+11ChUnwYSJaC3d5gm
vR2ppH7uMLMVpNzeagslsL4O/xQjRXALPmUemGrQsuvEgkLgDrO7BEbDFdUSZZcLx6am2C6jhiP6
sl7fJ2X8Hi2NkZnYpqW9IHQVtIkFJ/7Fb3Z0BOmr2XkhEKWfylZsmug3jIAyhvjPpwmu2iDBdAg4
r8/lAiHPXYYFtGG8SGeIGd65auC6vXYSMox22dP6Ki7LXivEUsljg1ib1cwArebn5uLkeJCt3eOh
EGnFS4AcPRI7Fz7UzoMTRRp9LYutTWd0HFf9VnajdVdiHWuAP4vLZQgH4EUSGFB+P33q0ZgNgUP1
iOYfp6UJytIETCDpwcLG5FL6Y1Xxj5urqzfdiha49vBGFDqIMYxcz2HArU0FiMH4nmu5BK+KjQX/
LsUI9PMDeGlUVHFN5k5QDI6FcLNX+YX5N6Lm0i7SWhmfc6umIgJumdh84i8IJH9+HIAyHhneDuJx
cb6nKgNtkWUHaDl3FvlNc5jzGdob98oRu2Hj+eUONnllksxAdPBijpfjY8z/EuQPjZTaFZkHV2rC
sezMS/0bdRzUVzLuydGngnKcEkaBZjMs8ocUVYH6p8pOSfWAq5Zavek3SsTw92eAPh+hxFfen015
LLXv76k5+jy8VjHc3rK1iqnLqyA41ILtp1/yoaBLtHPdUtcBzoE6TMI7uCgQ56w5M2EdnAOxak0+
OCLAjrT9TqHM1Ctk7oO2n2AIIJL3CcUm+KvycYoXTmdUemBaisvHHVBae7bP7/+h2vS+OS3qK1Xl
/yTZmYS+oYnapacOyL/h+9NpG3Wl5T4m/u1RvUtgDK3lfOTEcPqyc5AIcTRTGmyhaKUV5buT10lt
b5p466NcJqvN0EOitL+zJJF5R5QbRSCFHKzSulJunvjM6XHw0wj6+hGYXRrmpse0TR7WH44ZN+vJ
34PMfDzPxZSp6efLhEZvJCmKW2FlecxcLegQ5+uXboIjsXi7G1bNSmOP/gyn+bMdkF+i+p3YD1wq
JstDO8dz7qDjsgaEJrnIHVCqW9BUJQLTMwCIQENL1sPLbsRmYVdwlO6TsLBBRGFS/GEsPjuXF+vG
jBO8U2Uqqdax2lQ6/E2qCZ4mzjSHqRcI5MIFlABJ4udQhPi+KpvH670tCg/1NQwpUxyaxmt0jyXd
kZFQyfOMhJWnE9IOZ4cU9/PrA+YKIW+EkldgXTQthbS+ssX6arQ63HjOKm7sKNcCkWEeimMHsvyN
+Jz7Q8a9E9Yj8cgj1uerpJ/9kTyyI3JeAxbAB9i7DUFuu6N3leNZNE+yenHdIIzSYsQPXaWXI+Uy
qG13VpgVY2zWJ8nQm5T9z1HkVNeOPv7g7kSqbYMCL5DzpMSwWzMp5yPL7HsxMYnj2W12eHSkhmD0
8QWvE0l9r+Pi6PJ3mpnt59/SCME/YUtMeDjkUEjGhXEl39fRK7UWKruMpFsh0G7wfaRvDO/okftc
pEhUNoqZ7MQ1GnQcRXonIthbRdjnpAtXegpPstrvy9fb8w+Bqs17Uf3pAcv+BgmNc7h2tiG92xDp
9LGSL9uLmlLxCBsRtj42887DyHORXM1NxpKPAY5p2du1JhxnlLq8BUZkKJnVZPdKZNEPbo5Uf1Lz
gMrGkSyOM5MhssC3jHUg6Bvad1koxnUR4Kb0lJgWFl0s2l+dw/rLJZLsTLXBGiKOYiE2doL+0EHs
i10K1njxEz2AFua8GAGAprOZcY8xsIepcX0qt/6xpkbDrs3xKCwppjrUwPrBCKT8VMoxsmputQqV
gUDqa7N8d+xmjt1ggK/ibBHWyNReSyNUuU3ZowdObMblRszal92+nQtzJ7bh12aZoHH2/MNL+uAn
E9yITpArAgj5GF2dLBq18rm4s2A6suwpgkpUx3pp1MaVRnDOn1M3ErwxCYTD6P0LGURs0ekChR5u
N4HwV61az5+U8f3PtLyjyLE3oiekjFfmAZiY5B56z+pCyj9rhWwglfrdi2HtnV6+a4oWRrIAjD5Z
MCClANyKeKk5730HP2zf4k6N8zH7OIPiAgR8ikbtKxdXCARW3GJ8Z87N+g3ygfgAahvX+s+qXySH
Yk+osG6ZnoMr8ijz2q+Xw7x0/dLHOb9THllQu1FsxB6HqWgPtuzbJhGzvCtjDHTGkFIsrqK0wqbT
qCN/izLabWXpCYTV3wizxE8IbsC2cUz21YdZYl/ZjGljCYTKrA/8tsNsrFCt+lzs4/Ud1lpSrmGW
x7ZyoqFBkxuGUVOBvcrRygirDiQM+BIgT9nsP8izkGIObVLtLvcFddUcJl+kRGSQsrK+HOnTifHy
3iMVV06BY+foTSCdFJnOIUjdsEJxgc0huWOtzHTCTmLN1XDPLV6hkag8csM+pEvKGMWx/gx5Badd
itN3JFdlx9tzvEeTrcP6fh94FD8ywVUR3BVgAO6hjoO2rSYZl51rtgPyB7rWsuohjyvE8Eja6/yZ
v4ls3Zzd++W2dZe1ziJUIAZnul2YpysOXegN9pWtEWrFaAaaKtzDvRDLNDqHknfbUpEd9IQPRStJ
oznX9arSNMLKmOCiA9MpdSgReW16853A0t8ywURZnnCzfjwq35GXjHd+6W2S3mY1VbTGep/c6JDZ
+W4eQI5/hYYeTGgVI9CNtatDen2Avw5mOn1ywnV2eChm1lXgxDkyio3VSjDxmj9rAB2+hYOsQ0YB
gAhwaxH9TbveIbLhF15M0Wrng+TFcbD7CNZI4pVe+j/+hQlDcINxLkvF6T2gZZr2q6K3RKUdokzn
9pVQavmV+kPob5uAmt3gm3E9V9/cZA/aVipsP/MPpOfnSNkzhTr1tUGBfDZrUfjT++25dnNcj6jS
k1auXbEOTaM1eND7AhaMhgV5dAOAdqHhgRGCyUqsqL6FmOkGaDtw0B+2I9+eoHJjPXwFl3diJGLN
hjUNK+FZogjL0Q3V4fyIuY0wnGtPilXDbStw3I5MFuL8F5BQILumohlCPlpMhGHLGIF3JtJi/0Eo
QJ/8P+cdI9cOGgcZoDcLAAjpRH9SQSq7fWzGh9IZJPvgbeB/zacPDqqFTF8HzecazON7Ysxdh3y2
2ty3Vjih4F+aRMXnjbIbmkXjM9L6a2uW5hwrzKoMtg/FsfawJ854Xrv5BCqWDy2qepJ2bO9WlvQ/
1Zwps2kvl5AUfs362sS/pRGPNDJWLDw3kUKJFppyL0QzeIFaO+f+5eQqGll4htTyRAXNZ4vKUPkM
+Mmr73sR537y7WFPw2RollazvzdKp4FmcYIWf4cUZ8j6ebUuOgLj5gCt8VkLjRLszJBvp9Ro8gtK
e7DQ9l4JvabGlpCPMkONuRpdb10pbcVRdmXo4l5svs+uhwpi7dAS0E44lY8KhcJf4WrZhhjdDQXD
H2oG5gJfmc/NRwV6XVFe9M4Pbdy3Zj76c2Oza4jXhzgH7Lpo/oeEXYimmnVsBdl25WWLzqJzP2NT
tXEFNV7W+5EkveOAeLlfUfrFhL3i7PX242wt8cg+tpj/5JJ+Vho87YkNSWhuenbtkUXOGAN6tkXA
BA1GgKtvvUCIasvWtGupGGe6izPPk7E8IPN/9hOuGYoLINm2k+xj3rqFxa7+4c7tiS6S+JnFC4hS
SPTkjjVx0fXWXah5hRPmRAJJ8ZhClFIMbSwnpWv1yoTs0A2Zbkf3ZLtyvsdLjgryUKGGDjm0i+DT
c/0eCKui4+9PmOhtWoCFgfjOMZuv9sH+KZaBffuOaBuDg28lkM9NPFKMtJ2dpLwyYPdk+4LXy6zO
9wGnaGAH/pfVJZau41kGj3mdGxeZ9MJ2BVKl3qgSxx0NBSGMH+U71rodqD6j0NYBGRW42eQX4oP1
ZBCvP9jxPPXx7imaiXfYZRNTwRAOie4HIGSDklc+hn6NNhF7sSNaPBrdvubRppiYy6FLryxccEzU
q0DlP8kHsWFnFM2zxiWNdMjMYKEe2EW3pnOOJscDyPBcJwVFh9a8GqxDIWTKysh6+uW8WSRqnhic
e1ZXYG8VkFjBdVs0MzUq61lKWHDR4zryZjnpvmZ2pA7ZVo6WlNLNzUWV34yHNK/8EetNy4q40iw/
6s/bxxwJ/aOa1AGK+KyvQYtjRPUk4dlOVg5hzHKGqspLt/8DoN4/5hYqXv0vdCH+rOJx4C3PXySx
KDm8WZj52U8vPGHrpzvldAcyY4uRmNcBvAm4Sd3VFCtGzS/9HihActYOsBX5chGMVbXaCXm4lhwI
szM9ZGmbtkE610zEThXhlMiLnW8d8mSlimeQ98tZbG22Tt0fwwLORPdj4CtYV8KgPzzOPYi8AhAY
v0HfUarOxK9G2awpvpBTtKrzy0E+blGwnvGDw5D1TmzGiEfOPRUFEG3Qz8LzlB8XirAWJRxhmZf6
ZUkE443TJrVYLQ/PibugPxhScVR4W2z0J2F2tEpUi+4LL5qwxruRls/8KOabq9ULE3EJ2P66LP6t
oSagRVKyRmL0iPxOYcKa75RdG3Qs/1OwUYgBfINNt60wmOFx9KH9qV6TUmLyIJ0If+hpKDHYC+wv
xy2M8KTlqbMrTCaXojXrwH8FbMwVz5OPHdeV7NDHpa+PecWup59fo5BaiOHewDeEGad6UydoWQTp
y7g0/4q/13O0jyziiMEIj6AQ4xRqMVt4nAstGITXqhSv2QhEXW43AG7W+7r9YQ4JSb/sZFc8P0EV
/8LlpcMC30ERcNOm8j0J5UCHaSb4jveVix4HXi+vA5ZCqdJJxhBiuXyS5H4hdK7ZXOIG0z6J/XFf
ZUD2gk/8O0wwzCYRtioMX81u4uFqhW/Cb5kSscA6Vq6rOONkvA0juUKslpFc+d6XEqmtnwWKScfH
JYbXGEf9BCxTbs6TU0DA7hImYqtk77O3PHWHPYWUUFcX9tN3LI2jpAwmYFx9XYme+Tk4b0PomGxl
dH5wsxEVX69QqFpt5mQGrHWvDC6C34a+OT97wE0kji4/Kw0yM0NgxSySOq7C6dLYRevvxhKmt2ya
t1AjLQWO/5chiAWULQEld32MUE8JRlzJ/TRBs2w4uy/w6baMVIXCS1OaA79SROVaYQMHv+Lqafns
7pDmds0H3/2JJZ+fk3f31SKaavu562wD3G8340OlYA7MdfcadZK4NLnC+zGrLhiZqltvpsP4yZHW
kvFUgx3YqXgmi0rCfodE/9toib7QDrlzd6vFQCeU63txQGUTGlYp2iCsVM5Q9ArWnCa+0GrHy3hR
DB7Zo1H6mkaB6YvzfKHEI/DeylWv7XmnAMEWHOSWRjs7cgQclNL/2GvcJYCfE4fN5rf0JaYZ2VZY
JW4S6fUPHhgZ6Vd8BAKZTN81mVmkaF+eWAzn0CyX+ZNYK9chjFniV3RGOy/FUKrDYDEx4ibTYb/Y
X/mMzld9Cimp5+2O0OZv3LOZ2qztrdrdMSu8Gcnii2Ckxyolpu3mB21du4Xb7eC/Mc24OzeUxfuw
aN1T1xtV5Niiy+f4OO4cvc7G+l9M266BgrkN+uWdzr0M2F+lPOXKHPH4NAtvtVfdKQ/pijxn+/ii
TIYF2/GH/9cOx90ryJaXLNhEmhRiEY3sYf+C1Xs1p8tXMrT5Rmloc1C4W/fqtEmezF8OjgpiZiUM
/tQ/m9VoSZccrj/q8rSiL1tkD0LB0Rsdu6wcGKKcYWtwe7S4PerKlvvT1hFmdF6jPH6z4+Y915yr
8PqnaIC5LF4L43zsTn9mj+H2WO3vVHFcV+Lu8sZKUDl3yA6KD5uOkZawkGQSuwhRmWyH2plaQK2w
prKNR0FN/kD5iCO9oyYjpC52XX/6nSA0zU2P1XiI+rqFpbfd0FDb4IStivo7B5F9ue9e1G5eyGWU
OsYAQ/DAjBf26rC7lyqdqvBnccBwpzKH7uDTOBfP6BQiEnZp5tJYXR+86b0d2n9004/sasX02q5d
M9Ry8ecBf+KACdKk7KIpP4FXa7HCeqgDHzncwl4H6b2TdDLB1hqcfdOOg5avDt61kGfY4q3wFZf7
ws8Ub1kbRJ0FcXqN/XFA2bKXI1R7YljDjwg57seXvVRIrMCX7NjkHBazVe/VgPa7LakiplBVt8dP
/CFbLxliTsQel2NzVIlL/Z6JmZz4+4hz+ZlcwozyFMG6k7tgiO4ib6CtDpZ3o5D8k17fOcwFCCBr
MWnFzeMSpB9m2y6Fog1D2amldOD+hECUPrW7Foc5htLTjFjRhYrg/knE9DgoqKLqvnNaw4JukxLv
SaoXXry5CoHMI2d49BeDcswVdq+HYXyKaXJkA27lpd3Le9GhlcKfbBqQbqykxu0f5UKG2326Q+mo
7YsAlghHA9LUjtJzOroSoBuiAU/8IUWckmwAJoFOzyt0+6DlspCOoO93G7/Bj1pHJ0EumnOqdUf6
kmeVOvV+YokOJK4flbStWqMwed/BZY81ymeMk3Wvifz4j+Miqnq5kTUD+0WIKTFlfPH7kgwBfqOj
XM3Ch6ZH62HPdH7yeR2zMVETYubK46gJReUq368MvMhxITa4o3HYCCyBZhFPTVjjWpL2iIMSuWZj
SkMS4I2RVJxRINgQnlTKx4IRZ5tZrPsizNO7jvCOjyMinu/+fAsvAOP5XXuJcLDeT5qaWx/8yZbv
76oKaGhldvRtsg9xb/97GcsGfg2uLnkHVwJ9sy0hRWH3lY2NVD1R1iY/R+onI8Oq7XH0bXcV5R/1
EGjy4X3jSe0C53ZR3AzX3jTu4+z/a6GWUZo+bCM7tXfeSyFu3dlLpI94cwFGKxHi+2WKX1qZ1Nos
oZoK/JRS+iQfYdV4BsVqq1llynZC5SrEV+Nsr0N1d9z5iNhenYR9zk/18k4g5gUkYXhjBw/UPp8d
IvccqV1roQ/FQELUR30QBoTr/CWpISK1Yt8j0OOIVjnTNJ8HEA09zH53ayR2lFo7amT88vkBA/da
T+CWhsAESBqEMqaKQseFsohKvunW5A6qedAjqVihRysX/iznRlcq2FqMXtls8G7xUOj7hE/EIyfR
Xq1k/1Qw6oiPH0kEf/VELdhRKUIQ8T8TcXRNotaaGtKAUZvlh/4PPHM75o7kz/8AAZeJTtbQ1wXZ
vCywZh48MO7aw5VTz4WtDv8Y37kbV/bhCISQxyB62MJKgKpsDQ7x6rqsi9YOEySDdi8kC9Ikhcii
uSGJ9QhGCGnHf7Qo8UWL3GtYBNP1rpjYmsOEdE5gjLNhmiDbnOxckNyhEyMTpasCRGejoGpW5/Yi
TGQ+wwSn+JfmHZ5e/HLGYJd+ZTx9iblrkgZWJs6OJCQiR13sZSAm141uRSdZ0TGzv3gA/Bh33Wwf
aiYuQSBE7pz5SVKFrqtF7+rwGxTC9ryBdK6yyrH6nEPaSq6Ngk2HgHpxzEkIOKq5HesiorXL04Js
ZeUqt+rmJDGw1dxGB8wB527DDFyv3aSBzJxTdlJgGo7bvW3gUrAyb4nPfa7YQjmab2yNAITnLyna
RUlO8mvH/RDF3iIcHjmG/e1Wy5zIQour2/SDQQ8kdNyqOnrp8iDJ5jApJFq0AqerEQFZI1KHL8Xb
KFk1HwUjXNsUmmK4vtToaNnceg8dpyyFKflzmmfJpV+wVMZytN5rlVmshwB5Jm+V1vYCGcCX1ICT
PJTmio2ZD06S/e/RBNcZM2u8AUx8MRVrYvj6Z2ljrpoIOpAQwKaqNBLhtZ77JW5nOuu1EZHj3sQP
6Slsvp2L/9pQjvLdxRchGmj1S3M+hcfHO1A45gR9mZtttXSYl19eNSxU771TM7z5WShFBBRASLTP
n/ks5hizY1CkyRMeo4Ib9JQZqN6F79JNNinl+d5Rbd/CrTik/BVpkuU7J1DbYbDXDoXeJJ4U5psF
pq+UknIHwPzt/M5WEiXqSR3iY3v2vBdWNTPHGW9FzZ0SZoENN7B/3tFu8HwTF44dl7HAOXrk2MDd
oBnMJ7adge74Kmy9eQhRpI4RUbmT8Ki0ZOzc4SNHu/L0ITufGQWemC4Xce7qf5kl81njloNZAbHK
NZNVK+NWNxYnM9XmphEMxIObcfJicAwJSGGEbSWqPfKh87NdkeXlIzofZPmow5fs8DcfxXSazHLP
bz8sbj2OPp5dg2GJQQTSsINstQJElNgRDyK7wmnlHEAY9hehW4clqA+CeRLUzYx2IaHu9J2YuX/V
Js9doe0mZDrAre4nw438Sh1fZ6K0uY0hokfwg7AoURVhVgK8I5Nt59ve8Q1FFhm0AVA4bg1iZJOo
440XU+8xoPiDWve5frAUqk9Rtwrzz5SGoRdEgulSITC6uMbMBFhIPLwVUEHfZnTvvSo6THJbOfAy
VOFNaRN5oqaR9aduAY6WowwWupB8F2jhb+ltsYBgU1h7/1ghjBUtyvS7iPtOEOIXtNcGoTNjghPq
gZZetwFma3PGvKob+5pSD8qLWhB9+1U6KiJydhSsoGaVr3m1cDNGhYsSSSV61Bz3bktXPLdp8ANN
9Vs3WILwd1NrYVG5dqZ/5T0tLi6e2QvZo/gw6QAU97LwXKHgXRqANySRc2R5UvOM7ckufgW4O6Dh
vv36R5Gnoup77mjgZB9Z+crJSu7Tz57W3scepSnFxF/9oSanvwvNrIPbik93pO7VhO1J+Jaw4S2Q
6lmaPThnsu6L9PaLmq5CY9tlhnVUJVw8hXBSSauLqp0l/ET7ZgLiJLpyfxXi5LYeadUD2lZH5wgF
saDXxjBrVHt3R6WFtYhRqxQLFN/6wV7OqkA+7Jc30ZyVGBgPVbsS5IfeJ0YXJIDmD+j+/GC2c0Gd
iv1JcD80dq6GGjkMKBlS7rpyMoQ4VkHr9fMb57/Geg6FbnZhfFykIPA6XfYrevBZv3A5qCjd5LrH
HAgos3F9qU4vhTFqEqgV3E5dOAEvjDM3Xk4AjV0LxSfAQVUpVqHkttxSpxuL32p/6JBHwjHL9vj6
wBqdwhanmqXfuxu4I0TP2QtHOUf+fnAjwQSBH8NL0bIqW6JliZbf9ACcwkuIFOg4CVg5ABZbUt59
cjWsCHrE6uKXwn4XMfL6IGC4V5agr4FmICKPXt5MKch49T/nMAO8nNe7kvpl3h9EjGuGm+nMOwBm
R3z8PXPlw/nLDZP+5rjP/rTGYuLKHtH6PiKICaozr1aWpBoU+hAW4ogRM5/OYefUUAWA8gw/OV7O
uALFliGqeYSFFwWTCa6WsAATVYLIDWkuWyTq4fm3awXiBoEM+MxOI2uom/vBfpZMoUt7QK1vKW1a
3uZJkgiBZjiIZ4NNhZE6X5+G5kI5pFYrxCAdzgQAkGoyHwQQmCs2QdDH87Wf6QP8DN1Rx+YDFg1R
MCumpOpE6Teu9kf/JA8ff7gxRXqwlRsUCQ1dvBzwlsNBosGlfms631nLDk29RbjWoVVFxlhD8Rgd
tw0d8wxg+aeyxKEmcFY3vNGZA6o0exXhYV7PxJmk4wXtDnI/HnCP1q3NUP4IRe5lmw8Ws53UwUeq
6gC3x+DG07mybCeQo8za745zwo7mMQtw7WJuFJWZYEZ7dq7MHD+FZxMBGnAnhjMTdgqL+5l/ilXQ
NdIvARUkkorkIA0bzseYPK2nF0En9c9MCIBFTHNFG6hW/uvIx4OMt52duAEwKt9JRR1IdLVhjqd5
/6CguF3FymmY7AIMdUCGS5GHLCnPG91yI61ZcwtA3ENCOUAcKk5aQ5Y1m8mSu6BuV7ErFcp1PAB3
kbD9Ep8mmSSmL1mJ4XtklsDbgs3mwelKRtPd+6dM1kL4BCe4ULzF3Sbh+axQZdVt2v9SPFDTl5no
/6fILQniYTa69LZn8ikjWn94IMC8ODHTk1iSeLWEptK1h5/KGYVAd6T2qZoGw2MntHJIAhm7woeq
Xhm3hm2WkG5utmpuOvLvOBlyFyaT5hRgULtIH8FNTCmkBHNbEF1vTXcgwBKGCxLP+yy4TgLuOm2w
cqRWEon+EeB/yZTVa+o+Ib0Gd/C4XHZymCL5RsgKlkd9YqZHEu6jLCfesDxx0is3JQYet4tdr/w5
eG6Pmx572ah9QjPSSndIr0uQmzWKe8BjoHvn1TOAbNC54h3m1RUwx2ty+3iXL9ghSk5oH8VLkzRC
tLpg0lMpBTOaP+prlwlUdQLHPoVWa++lZu5lHWNC05j0UkNVn9XBRv3N3lvv7OMrYUYBY6iDL3PL
91W2knFr4gd9/buDJsc5a/04G4htUz3ddDLPOtJXmDTXl+hJGVWobGIco8DOI+3hZ10Ocpe0G5uk
G4grdLZM85EhiIbEnICZNiGO+f4gnSR6akC+1kDyectBjqNOZVIz8PzUCl9E3SADh8Jf6/M9xWPV
uXsPKLylMsV4gvQVyPQ8/YEpGOzeXzxX46DnjVT8f5SGm8HTX0DQqz66F+UEjS8wdAn/oKUuVeR0
6H9G9k5nmEMLEIP3QELd/0wRtOZtaaDU4y25Qm3X4cScBHdmyMuasW/8BS3i1Vo9+S9uK7u9U89c
HTIgNXL10kKvq4KkqyCGbq2QhfoBhZwKJP9SzpHZbDiyZg0H7kXfQ9BJxHUs2X86gbMhhLowzA6m
4SPN2o0HUjzez8CZnyTJHUTgjo2cWMcRPBnkGskRdsbcwt9lY3T5ZKA4QDAcWBUqb9nv+0IIg84/
aMx4Wdwy181qNweZAOPUq7jooo/cIkblBobuN/S2jH5SwGQoTkgC8e/Dfgi5I/pZiS656Apdc0/j
ERG33XGQVd/v+P0sxkmxxhoDnxTlEj8bNIJ6o5OdUYPl+8As2npz7H/iBpBQqS92kFKAMm4gQBR6
VFcZ+10YdNKeHxPoXa0rKMz4Y/q8Nn046A93YFr9RCI+6Oq+BJWhupbdjXadW5ZvtGRoCfGy+Btp
Z4sqYnW/XV9B+lpFYbMpDc/uuFtQ25TUbDF1yqEW0OQxDp/jDqxwc4duElk2ZWq+L0VzH6SQV809
frBH/VAfBRmpmDaP3U52zQzp2uMoGKBmx9iNkeSxfJnYDBe8y8yyEfaqA7pE84tERHFlUWI4cmiy
J5b2kkNK9pUkjxsvvUoNsBcr9nVF+r9XYBRJ0x0SLt0AT+v4ReIQkc/QExjpiW+KsBwBpbtBLOmt
ncplEsDXtD9xlpWvuBS0dIwJkWY7A7jk0p+Sa2RmNyjGC+X8gNnPKqVllGc1k10DHIZ3furhsAs8
6YAtWuthkUNhIa0X0DHguWijJgeBQIx2XI7nMroT3qGxiMLfWXQZXeqeHLtB692qqVK0ZWJS7jJB
lkf/440Nnup8/afUNXdM7ef4RgIIwIi3QBNuH6ZBkiEMwBEySzHnT/MWpfwT4m9TrDLNaI6RD17y
rfZe4D7I9+/actPYTxReOSVLioA3YRym5bKgXiLCErCUiKY673fxPaJcvsufP4O/YnVOmbI36un9
PL26Tpxzk/W8Kqvw/1ABlKwA6Shsms12k1dCCWJhXqF9xE2Hcy6zTAoHfJdnCvE9+t+0EwKMOl5X
W/xWMqj92LMs4kXFdp8pf8we7vZYzF3cN80HgvKmetYt18frEz+JsCzY2esL2tQtiDppztqTdFaR
nvJnEpzW6pzexjXddOgWnqjmwCKHPBWNw0NT0SZ5FWeu5Ca536OTHM4e8f7TfDvVBKiaX5Dvcjo5
XdxBUkBU6OJcXZ9Et19tYErycIrEm9rZOSWWh9LE1Cf5YBB/z1Adv4+LU1k7BjPF6/5TFrYhJqdo
ITIuqXLmvrmPVFRzS8lOahCGFoJr3CbM1yHuvn+UiNXb++H2vwpIzUxm0iaTNy1MdjaehOOJr6l7
wxW123ofsDEXAYtxC6CXn8L6ADTwLKBTdcUDzs9HhVa3YOirhAFNZGBMsxa2NQ/RFq9d28cZfBgH
hLmXtwx1HoD4cNb/IuvE2vLpdpUR/arrtUYfFGpvRgSdnaUn+R4NbAp3LMxqqzcQhb/IURlswNmd
9b0Hx4fjXY4hb+krC6M/VAA2d0++fGOJmmuS8I0R3ANIg6JN5kRhxYvErQ/J9FQTW+eflhpt+lbx
8evEUSDf9HfFbZ6TiiAgZGERuIDlcoEeqcRVFxhnrTGnMOz1s4rivRwtxrpna8+px29estkwwbx/
Q6aDY9PfbLoAcCsbhG7JrtXL0335t6QElqmDGwkaFHSzyI5WQgUH5njHdzaMFRkWdpUaSQYqhe0z
ASCEa8n7VvNdfg+7kXfBzIsDq4zxcaingucq4I6Mli6yFGE9SFCQxSdIKKH2hhhG+l9v2jF6fR8r
kP7LjV7D9jFXLVN8HjgsWfgQhrc9zWHsh5QgtoJuTLQcrs1YDp0eQ3oB/B6Kt+szLpf/K7m+gtMM
jqsSkRToer9HXId2wCBDzI+Jn612ZtI586Jq3oPpIpKTjwmMFqs460/0RWURc6urMs7YR3T6eehS
J5z/CIttyplo8xgIk+we0mLKgbsml1lWQhJWMcqvxqYvq/5wVAXDqDLu++p1WMDUYR+WGhpqvRCi
tUOjFxl+uTBTm3TCQBl3zWvP9XZABId6rVLkFRHbDKYG7xLZvSi3Ny5wMCaVyse9XGTbSubfSCZH
qVE49Wi+xaRItCMbU6m74+nWFm+vJ3a+qtDFohHjlzTsgwbhYBWt8CXCb9hH/1HE/v+2wFTednj9
ieS+3PjLCWuQyF2caXSzD8z2wR9PTaV3V6L4xYH/srZ1TCUZN6ka4M5qHwK499P4xdiG5y8TBOmQ
1ogYIKnpQ7n36jFiho7vp3hgWuj6S9agJbefmuIgD5542RFlutn+kLBIaqCmc+wJ+1qmIGo9XdnP
5UnOfvN9R/1aQxcfk7i8bO7FswqyowK3Kw8Zi9uwNb6nkmUCJ0p2zStOizK8uUotHY566zNFNNhn
WLm8azF8j6p6q2y3meRhb3SGNjLLvUw7OBWx8wE2RdWA1XHKh9i93YKcuy/DHOhEe/8vJSx/1Uyx
0GhOvfozAgGSyEFqnWJCKJEfQIvYYIzZCrSDmaeGQwC6NrbKTwm70Ynu2BOVfRcSM9orxiB9FA6j
5v54j7wBTfuxpdtUY3H7/DZYufz0R6DgDgTH67IXXqvFE1ZkhGKPvxKFVaeFRyh9XHQvhSxzc18D
/j0AJw81L9mdXOXKfHUfTriLz2JM+sR2vZ3R0NSEzArqEYI1a2QKNT5JWsbkF/PLhRPaoPgWAHoV
UehTIejnnWvhsqIBdXnwF0PNJ88WLDUK3l4ZfP7/l7Evj38PX76Ov8Y7Sy6qSsO6neS5pLARVgVg
AJgALJdC36F5UpZ+ncCjykb++mhNUriDr3MRlqAmC8umJD6joVq1+g9nusqK0mjtHABRm2wmS+73
H4wLmOq5LXaw5GeAlXnKqY2ql93dcINGsrG7JyBiETFzoU4NVeYUJFUTGzWMy3S43wKRFwsNjcPt
8IsXFljVB/HB77oe8oxDDrTvmbVyK3UwZStusJui20/lSbk4epJZ9xNBCTbck3JOJUeZr8OxI5SR
/3/3TXiTHYJgh54vM2kgBhTeeSl6r4SKGCbrlgShhzO09SzMEBlNAX8Nos9BEjRrmQXTBSH7wNDR
cwMRYqKGPtVvuEKp5hb0gt9X74PCRGHPTcLdnrEcZwWl5d4Pu03ucBhbaPPhj6CXf3TfG/BXJ0jh
/lKRo1Ch/w9RG34cRnx73wyFNC7UZDhmxCNnqmzG4c8wcDsKkieqq+Ot2sieCj/R5MFbLgZcqZhq
SQ61Q2pXw44G+eQ9AEG+Hz8BWtnNdSLnAxtw7mCa6mErUSKSZUHTB7DVrQ19CduUQ2G0vOUe58kE
eb/HmT7q0XgfTqHnK8FHg5isL9ebTpxDeKoFrFJjIQQ0STSelb4TsAcme/inSJSkZweHtwMEeaDe
mxTqpzVdcr0FAzzlxcE7OEeQAkc6JiYobCnx17L9sV2yOXUkhMJvV4WL6fHEc6hhQZAAcQSqLitD
ozRjuN3/RPVGtoxob5c8Ox14DyFeaWY0MDuFf9yanlIN7dRtFfs/j/KgDcxIjJ3kk8VqAbOHCTjO
xqhsPBnoQZJzu48y0/+zwvlwJNQbS+RBQty9S5r1Zedu48cijdTZHdUGfkasVH4ydzOHF7ZhTX5D
R6ZLYr1AZf9faa31jM9buoWoL2XQJfIQwD6nVfwvG4hlB5JgqOOcd+a95CB6V3dsET8YE7b+yA7d
pyeit8twMBZg0wujCF936d+xRayvxw9NH8RdhRmkSz8OFH36bhu8njOHPArOP6WRx+Do927ZQjAJ
d/y4U0T6SqQXZ2olYraDG4zf35fAgFRbMaYpnBfCfzKcgZEkLUv9Ne0+8jb3HYvYVPBTXOE0TCU+
+xElyUilnjgewT8MwmSJDNPaZphvJnU9dq/HwS4h/G/GMnz+eoD8md1Kp5ipOmja/rZ5YEYif/bv
77B2k4d8UCAslemE9ikujH8wqIrIMIfCEa/LUtPiqSBExvEg1bal6nbCrVnPZl9inYB2m6uyLA5T
tMmfEPOimgYfnUIMCmKFNTZhh89uMQjVwv/ia6bbnQR2iKcXK4wVNBAr4aBOSN5FC5Bz1/aI3RFG
xhIjWA0KFTRmzslJQotg/oV0t8wDIHHzWs8Glvbj7+vXV4P2Q+IKp5Jy5qEeYcx94tZAW7NPDlBy
Z1Vs3IzekUK0qOiDTfu6xHtwpnou9VoFC1u/CH5Gzv8sLuoSooNIo2Zo/qmKv9qVoRVuov4KeUay
uw51Cnzs5FFHeIXPfWf9RBZwPI9W+xYISFW7AtHhhz/mWzmHUeNClWhe3s8b36aS89ARNeIoQPJy
Ubvgj31syXS3BWsGhogJ5dDdrM7qJkkCEorZvVM0hv+f+ARgz/I1NnnkbvjEQrEo1+axYU1iRxew
dmTxEDcnwhSKKkwELIczSYPldnMXEAl5SNjSn0Gs5Aj6TPH3BQROE8Xb3TCLZM7WiiFymfJuS+kB
7N+4sYcRbAS5GS4QVL3GGUMtjaph/hYEmU6y/41syhfpzFU2y/0riDRVispKCKGoX5hO0dBml7q5
0Qj1UYzONXDuUZeZv2xhsP0vs4opHQdswIsaxTtn2VCmW0gc10MWdPfG8qzrdttgTHfgQsGJA7iS
0937savjXvrvNKDhjbNK4/Oha+/FQGQTyMyBKOBe95fn+SBBTIUUiRMOqWeEgEDBaPM5dWQaNLkm
8NHaY+FJzccltXC+jFVPg8hxoeBj4O/Xbl/smcZCs8YMXo/1ntFsdPS9UWd/H6TX3JLoDjeIld6y
RnpDv0AwW1O54T4vk+iNDDEjAxGYgIgs+Ojy8s1KqCSLWy3AqMslv4Ts6WMryeoTeHFhoZ/BTTFC
pojLnrPbG1HG2Thv9Oowg5Z1SlWjnwRbE8gTgoYsLeOGhJU95S0cY1nxOcjl0noeji1/GZpBTO4C
XZHNxLebFpi6GcPwiiNgYzaLxOJyb41nJGCgY5QvdK6G/GJrm8FiwnzT4ElKPVVw+pa9fu9DoPPe
2/TwDL4rNh1zlTPqZKdg6XP9j+Bx1SU2cXrw/w2PqV5fsv4JDJ1Gqm/kXQ+sUAmzEaG5cO4b2Vda
1q+6XciiguDc3b/wkxB8sIn89iwVCUYRTHbiipBIL3f6ns6UzTMOVGe/beN741/BgPBkjngaHFX9
qrEq1EXvAqY64zwz3oBFXwJtcYu11HXlWZlIjM1acAV3K+xtkgCN5AfFBELrU4jbb2gd5+4aBMlo
5uzW1FFyKHC7JYHf+F10pleKoNreDw7tYbbWcMwBzbC/X8iJ2W6Uls6e1aJaRPUvExs5AiITi2SP
JumjadW5PYpLwwwceMfUXfhSBJ1Kzmhnk8kuSsayjFFrSQCpZEJsv+c/iZWuuy3tCGb85c2inXDe
7prZb9rpdg2aKXnpWk8HtOcRn6zJOUekVCxnDpHIYL702IqsMQW/Tol9d2SeduTwLx3oJP7As3f+
IkB09kI2rKZ0IgXQeI3eQFEzGeletbd2fdk5QnBt7vupQtdUGMa74gEQx6mCnQF7KjJ5on7opjii
Dy+yIQtcyMKqKlgZzdINQ+EkfPrJIkOvlV3A2WAp3p0DazUy2bUcxv/jzlARjb0Psh0GW761+dMv
K2qwCt9It6vPCmZUUmxnTHy02sRaE31FTUwiSJyOCAxelSkyW4tYvdGkJb0uYGmt0AjX3twH2b/s
UOyUleuNF7csozfpC6srcIBFR8nnWxVSrR2xd8OaRJGx90BD+4yFUL5SkMbS8u6c38IV23WMb+C5
zGNDlbY4WU1s0ps6MJ/tdDfqAbHZaUspgMzcvhcARZyZUJBXMRHdNDwll6YGmfQyNzwc8AQnByb+
eMjny19vebO6sVBJM0e2Q61e68OILvWjwzikt0cxPgNsd4Vj2zpWG5r6osjfZ73SCDmF3bHeB+8J
l+RTxtunArnBqEFbVnZ5n4USjN1getW+GvZFaKYO2wnjVs6BFNUxL3ghdQ44B8ARdxHAf30yXRhL
nTfgnoIZpI2mZuWt/PUxNXddLm9/GOTGkhl1aNg+cwiW06wV2NGsEkgYnl/vGlHGreVyFYFLZDvX
VFTpJSckiHQNnlmS5Pjrw93QliuprHg9IN1zhxOJH2E4D2QgVeK4gGFCG2jJIhi4U1YYNnXdhYSa
6xRGHV/eLKY32rHBWUQG4I1X2YNL6F4Etj+VhFTwaktbhsJkEJ2TEITtwB80BPvonm1KxOrfx2Df
RjjBe54pimZtYeCrNBeuqn6QqZ8Fl2/APDA0hkMysF6jX0tlRA3kHO4f//K96HPwYG4gcpfyItSo
C6UeqDR51GA8VPbbD4HJTxkXKov3FGXROu86AAGxBQlXk8UrfgaT/vlvCuxeXJ6VUq9+ko6kitTg
YiV1ZhPPZC3sZGiJOvR7K/aMdzP1S+RGvMzo6f6kJzs2fS7IZV7QPK7qRF9g1BeMBBjBAwroMZ2p
gHaIv/6Wf2HInb7akScHD/4rstxA1V5WLJ5gID3mtjy8V8kCv+K1OY3yFAzvuS0Pm3C6+/8uIuEj
msIM04AIDObfKDUaAhZJV8cxK7qRSAfq+0d5u+vDXHTPc9lknQAags+dvnVmjt3+yDWPMosMls9J
6ko9VGV1TOsjjcMvzvtZb2mGr+uli0Su4ilrcQBlSyprUslqBMW1yQoqvByKs+9HHXpmDRDaHlay
OvUoEwecxQoe7BlroyUNzucwhhzsQ6rg6ePHEu6c3UPyNE7pzq0qmcryK9Z6QD8SFkFUExwZVqkr
O+EjpSdcQMR6o5xcgHB1YIeaIIb63hiXhoq2h9qWMtzR9lcLiEJt2ueQsbQDx2jIYeOgWZBKspKh
oZ4hVydCUGWdsMWMAhSkvM79ddAtMGit/1ZlkCpqChs6w7QEgE6dE1mbsT4hP939owOIpPygauZe
ftUVwGoOeIvogvUxvjfPLxxB8U0fj+La/xI5F4LgbGw/7fLF2D5WZbG8JdIqEzlKo8C0YjdkoW7h
sdvZina5ZKJPyQoid7MoCUecb8b4lPBL7r2OKLITqjb8SsnHUCT/TuVPnGSl0aJyJf6sUVxFQbQq
k42tzip1Z/XeGpfdIrst3cK+NxSzCj1pxIobiGxizJAr9vtpKAAhH/cUu3Pjq0Bmu/4uX3X4wfR6
vqljaSuGW3lebnUQv/IZNrJGgveNDsRMMq5zA/9BYcWY9vqbXuK6JfAG89Bc/hcEjWpe8sLVEMCW
ewvIejPt9xigVJZrbtrJlDLWLp7+ICSjLQRc9FecGMbbNyYhvmjOnXD3nww1P40BQ75L9ld7Jrey
gg+W4/IkAGRbqV91VCv3LE0YqUIP3ZrkX42DkSsYypKW7R1+WAhxqr03o81304aOsjVAoBO/Wo9w
0dAqxWCiXNBLeAbATBfEz/tnUjleYSMB/i5HmKkPP/eaLsOE+G+PsbB9WUc4Y5YVOOTRcZSMqjbp
mIWM1NQhGy3GWpCS6iMi8fSZ1hGUwXkgQBUpUan1rQqt0AOOdg0eRYnYgA7T8SRGAh90uZDUFWRW
7W8W6CUj0tJlz9FXJMI41l6qN8NRz9gu7l2Njo0YbbfKUulGnGkYLBXUBYiL6BypP6Q15d08siJA
onVYkDwxPZACY6/nXTGJIX8cYv9OColbi8++GsuktVkJxYYv7DUIaQCwKkWqe+FE+ZVIq/3g0iYJ
tTwRsv2M/8kWc/ZiE+xyxha+WMEUqYNYpFMG7e2m6JcJjsUYN8IE8y+aMOuOQAQVUaG413exdjpH
8UljOZJ4DfiStLC0jNkjJ9K/pzxASY24/ZcYc/fdHBjEp2MEutBuoHLwHL3lgJLUT0vrsIz9aFVl
VCJglniz0dwFTcdaQ6rvh2o5mi5XUHzjH6pmcN0dQUXxCCr/yWWjROp1fb71KXPTLWtmMZyXQAfM
CXB73fWsDV+zgZdvh3GY2cZvjfygvMr4jV8hDs93o5u6DgSnjEshRlG3O/LGvoTQIcEuwVM4mEpU
3fT9o/c3j7qLZhxQe80wHRxZZpEry5yXDXlCoBG2GQrCHNpuJ5N+Osz6hlFQkAbDH9NqoX2b1yKI
JOSYv/IgyO8bv5iAc1ZJaB2aJSH3qbel8BnWi7yNVzazM+w0GIU8TJihfOrBjNsSObDY45hAP95P
CIw7Gpp0MUPRDVulMmEP0UktlTofeao6Q5LbOaiaXiF4xu3gbx3hD134wtw2lGWJ3VWVXmzz2+Io
HrNaUHE9rlIlrHKFFPT49V/EzjJlZ2gWkHzertVedqDYhM1OJEe6K9Y7UgSrHIySTRe+9qmrKjJv
E55m30Uo61ldewcmJZHHBrQuz45buM+MhVW5+jo6eaUjxmdhdKX6kKd8aPSHwl3Y3+7sKUCW+5Hl
CTRTwvr6FyDyUvvtk5LuM89/kL50yR6EWBKUABr+qmWseoVDJ81+3mYMVRA+Ug9JsDfOHy8qUZkx
QhP7npUPaYpX1n0SXXuxXHMdey2qWsNL0DcEMcnoVGfBctpmZppYIWcwQg7t3Q+rBoyVdtPOBX0C
VPun7K58OTPEbpw8GVmRtJYE6DLVAjmvrlyJ594Xm1UiDaABwb9gXcWne6GfU41SgmqbnFW5ywH/
X3qgXC6oq5d/Eb79kTNMV5sdUPZPM4qY4Vpdenk6PIOS8gHX/EIAvXr2zVy5ODYN4kmJA+YLDIEB
30zARZpkj3nA91RrPG8kBYJ+X5nNnJOaS265xRC++6tWkv+6YoBNUTZnk8NwmSSQkH3Duc0/pYw2
VnRnxSh9qrVTD4xmhRtR1GKhUA5EnP3tXHuDhOr4+PvpaKZHeGFtKTLXRpP2HIJB+lmtBeuUNRps
vzAF9iRgpzQ/IxgpfueueL45IfGExAmKDjPG089oIRn2omcXXTrqhLLLskts6ne0nhBOCwbfyKmd
uX7cYNvv/G916ouPSVZGnYxiBn2nnQC4gaPukS9Pn+b+I9lM8UXa9ie/wxPohLO9EcvLQKKyn+Tb
8xzYNDdZ4Sdx+yKg0k4lpqeLCJITjQHfrUDGbFt/qWPOqRnZtBm/sAXgtIZxFuJK6WGlgi7prfPc
EE3dKF9JaXpgyp6Y64Xd6J49ATq/6hSe5TvyeZCv+aFJmyNR58ux1IcEkmRt3xTcvrvtlEvTG19V
wIoW+vv8x9SecGctktqdSQeqs5xDEuLCnYEzaPr28Wc8oqPuf7iJiOlNohFVA3b/QOMMFm4eJhFO
ZqI8+HNO9GxHa9M0gt+jcj9fLGTxxbIKNDwJeblpkZKBF+jny12MhGtr6hEZrcyuERnMjMrtWw5A
Qcy9oEoNE2nmtt7vj5P3NY4/NEDGorqisAEcWi2LITmq5Gusof2/BxSoeiPCUYuh5n5KEBla11t0
IJ1Ok5RW6uUD3avtp+Dd93+ju84C+rOBKtQabplfV27rBHRoXlQecyDTdMINgLFsLXhtTQO76gTz
/QsKtMkKWq2R6Ir9EKH2vh7x5DyphA55EGPxcf+JgnL/wNDrW7A5SwQEzkG12EsdmavHPgMp6oGu
N0/sciOeIZ6acnm3i0XeI1an9MXJpflXYnECifdVuVAkUN8fugSfe2+H+/73fsSl/6GUWkndF4XT
+3Jb6m9Y79H956xYISAZSmv03PesFzTZKekAicZE4ZSBljiFUc/PX25c7EZ/YL++9yrX9Z8wMMCF
Us5+345aHTCpvocbCNgltukJHa4YXz9lpPjMnxONNe4tnwLhRKJOfClV4HrSRStwHr/PGKYbcuAb
0qgk2r4HRwqM0VdsnaBfuwRIWhGzOj89eb/HlrxebDm3ZtTWMLgG/hyg5UKHb4ww0ROxBVd5Tn9f
5m6ri+Y3zSkGACy0fCJHvpPKkKjVxKbuE3FJ22oQBUB6ABQaTBy1y/Q2azCdj71bvIrwKmdTlFtB
qBgumwn+SV7nWme+M50SseENe/0rsdjObeMJcsnXe0L9Aw/PFUVbPoTCJId5Baf4IZVPn+5DcbpX
R/UUpx9g00mc4IUXjyuFXInDplJPDfW/NZcO9xumHbkBIIa/q1rUe3eiW0arX71DrQ1t/79MePPA
3CPLLp83eNDzTAKETTMW+XKFGmke43I0y8gzhGeQUJugOWPSimztD6rGYAjbYG8x5CqCqyb2CyzS
JWLqyfpDvYiniJ/z2PNzo50njdZSZvFhoW/ZGR/ubRwFfcYxXO86b+FP+2FY8UFYMxXjNJOMsy/4
/Hl7X6/NFPELhbyXNWpfu/PzD/YXJ/WopjoM7fGQrOmBSRQiH9TPSVjCHgJYOWEZhD0ZfsXExjpk
sZ3BSmOmobFZoAFOJuN6sxuCeH/NQueE5n5luJo/eRTAGibRxfqLwy96becWb1rcc6nvmlqRGFV/
XV8QmBrN8TQs51NKPZ9orSbY/qpXvbHBmyFtbsM5FTr84CnGeNdaqKD551fiUfLJgEiI/ajm6sLF
QrsmpwkwTd07aTT2rLT/5u9XvFUy6EctphknDrbQHwPBdkf68sPVIMXkGory1bQWDJS9leS8wLkC
44fXX1jn0sXI2+I0Blu7T0pO7YhuHhzrojx7iB8OD8LE2uPGPSAW+f4UtmULKdiywSLZ+pnmr9Rg
5Dd+vvjSPk1msDBTTdV8097yyS/PlF5G1uIPk/RecZ6uZcG4OaflqtrFOfcpNawjBzPenQw2g7sI
xcvDx/zg9Mycy4lRQ5IHskne9CUTlrd3doQ67esNiolIyb4dUw4AYP2+IPah/Qww0YqNgVmMZD0H
3EZJofU3rZD+l/4rq+thC44vAM5fGoXK8G2neKyHI1nqU3jjQBJueBvGoEAXI36XFWB2IdXjzvJN
56SAR3ikV6NkrQS9O9jX8EK5l9q/MS2nt41qvN2c9UV7wFi/B3P0hX9RdzF8wrwM9yVD+HsRglkX
Ba9T908UyhGqQpZfe9Nq/lq4l00hYMm4CVBGud3H1fcPz8xZbV6x6j3sHCt6TcUgxeosCUFrXWK+
3nVKEtEDjjGa7ZKW0H45g9S6EZ51I3jJR3uP56wAD8lDHrpjktz0KIQ4sQ9RIax1f+VK55Vz9jOl
YfF79yV/UU1IERO4U9UTzVN/hf9ect2ULe54tF4aA+Ux6L3C2Noy8vkxhmWY7XbPGXzFrCEauhOM
0B2cQBRTxjMLTOoOW7b5EyrzrCJuQkxkzbp6BGEK1Vv+HlbHJIvV9WNNCXMp2fBw633/zIk5wy3d
vgViZJaHuvsLRkYzGYEr3XHur7HfHfqNoDF5ph+2UQmO6vz58Z2rX9fxu4T1ixUaIheF5m5OILtg
A1Vrjd9wSYBqkg9nl7sUP4EjHyaexLgqX+NyWwH4WpgXfH021jg619yoTBtCgyu2tC4LFUo3To4b
pz6kxwscBVhU6M21TN5A6sTfnleBkWtiX7J/oN1HUtXuXCrgt8KGtMyd9h++IR9YN3ZL1mPAKaLv
Zzp1Ru9Q9cR33TjeEm21jLlKy9pdtijVrY6yCaBR3y08YhDMpNry59H83kPOAaetmEHTivjVko+Y
QV6QqzMhMqREU5QXx2jhRfxoJLOk4Vsrb4gOcP6Ed4IheRL8BFXqkYHv4mq+XJojOPm+FX7Ce3Ww
VKNpKLxPbSjYYhRnZ/bUa7y8hOL5vOvufJeGlNe0Q074GySB7UNE5X6p2tSCsZQXWd3M4LxEhK/h
JLhMRpxdvdTNCnQLqZXabjpTPo9KJ2iFNHnFwAkrDbukF9287ijMEs//hovywJmf4vzlDD3QbtS+
2usUdsv36/9Xkp/JY6Q2stuwP78D7Ir+OSmuh/W2rLGyjV0fG96+2zIV0q1A21B7V7L5yX+D1QZO
a2FVO4oFScxEtqC2BM+4o78NgdWw2xoYgelCqXSLMByKgDFDlqZxsJwnsPxw818rPKg9wfdwIjzx
PEQBNR94bfp2l49KsoGPswU5rDKwtpp3Hx5e0q7LR22s2weg1ZvfUYHdoAmcjszY5sZjz7d/zrjz
iJeuhvrAcJNpUqGHn5lquHhnlh9KO22BOBdu1A4Wws8NsiQe9/H7JZaJ+2KrCN0vjZCTMlN2Q2q/
yxI5BmB7MoeDt7ePJ1LSx5MfV/96/a7yM+kOY8aVYSAOvZQADAOIEZs+TzAz51b+XxieE6rs0EZW
mGO739fCys6mn52dr4JONUMPEclu9dNSv0PRapgwGXNlmRKFwx1yMHmf/aIZehish/JapAqvQr65
Wf8pslrKbMZS6U108EglcCFutlMub/O6H4TJB+nSBEcA2ibZwqkjWUVh9SZS58vL7uKijq6NEnpp
tJj9KbYGPwS3JFzYt6WxYveqsocq/IFqfJ9e2e52nolnqQPu3Y5PgzYqMcpfX1z0HtI3YKyrT5TO
jOPCytH3yFFEdd2+yHO9GdYYYfxQo4HJt/8XKzSa2zaFfVBRAYPqWZeJabOco0pYyf8eiKQJdCv6
igYlqXqPqouDi+83N7K9D/6iGm7f28tEnYOEuPmEaC07x2UW+xxbAS7yTb0BH11aHBpiS/3pDtBw
gvBwvMxJP8Bu9kVaZh1L/k//RVpOQl2fEAAVkUgJ0Y5r/g6HEV0VICd6A3uuT2NZ87XcFw/qjOOh
AilOr0AyErYwEz4QTMhpa+4z6Umqlhg/90pMdxO42DOnUWIa886OIKeK79xp7xCQW//1PqwT65FM
p9Ro8PayFGMoxmBPp0Ztuo1+6zljpbPvn25acM9OZyXys5LPkpzx2TBFdUhaReZaRuvC9SG3+w0F
AWQhF4vP78ViXwGKD7knl7Zd/ZjOPdoqu7h+TnQmr9frtXvlYQTtMTxMo47LuJEQ6Rvjw6gXxluT
2T/ignxOR3OHFnHR6sB1imMTy3aOW5EdytuBl2+EUacYCXu9WA7qXuaqk7fqWFPrzuXw/558wplk
Mqqz7VqCxmcJXyq8XHK2+6kuwFHvo3kNoVPyPZ1cUg9G+Jb5Ml8+CMa7Uo3sxfhGs+NENReoIelZ
KiQeAwGzbTyE6azL4qvGov7Wydo0y85f15lMZqSQl9+cazD6Uc8gR7HcqEvg4hJz4ZrTGZHOBmh8
rAuUJ5/RUdmyhqyXxuPS3bkDbYpsXWpw77n5LaQciuQSwtVX6BnNtA02MP5KXWWkCVK+zRNoRqr1
YABeo1Nu6lbOYMPdK31sqf56IvQR+qTCy6uQ7VmTnieU9qPFtqzOpSur5rIMjdMM601kY0rwyJXg
Jc2Vhr5uuu/I7ykjAMIQvtYRp5QSnP0MaJ9zVtXbd8961dUxb1FmNGKCFp4NG4IwA17wrtTaEpLP
OIuKxZEEeGMyY/HxO0IfQ7LnPEzWN/gnrXItodxs3NomOlfAZey5bq4Fm8OYeialWS32ZwQ8ETw+
rLXwwwr9tzl28CnLSZwjagUG6hxblfha+nZNeBcXoN+dba2gdsJJLFSakHJ2Ucdq50v3HO/oLicA
PZMT5/Uh8X40TPmD5Ok4KPE38NWkETFY/pR6WWgQwGx77WMHOolvtYiq5PIshkQJmaYG1gWchuJF
eRBFOXGKnPGb5458dCcPfZA0xxmrmefVKk4B9TGwZWEKVNkoKG+c2xFdtkTl464wt2tkJAZN/xdk
zGSvmxI5VPcZ66wfGfAi9QSyAuLagi/iUU7Khat4OqpFLwU/MzO/TTelxduz0sCl8XAKZyB4ImVa
QV3LxfD3AmV7x+8p21bQhM2F55JblDTnt/Aw0DT7eEJfbDtEEr1086u6Sz+rlCvzFc2YdrOX4VyL
XCW4Qnfsh4vKexZ31cB7xvzk5FuM2Uukb5EwI3wAf0uIjqgnaMFbz8TMOtZTt2RHZAHopQfd7V3j
z5TvxOnXu907MBRoE0IgMgdtQIQFTm5nJK3TkTaS7WqIf4UTnBl4Mz1XXNyQXaGEOx1mL6clRG2U
l0L6HYaqivw9LKvMP9/MNxG/nHFv1d4IYa3Dg1sUrGeFDgcXYBjG5v/u+qlnL+Zatc5mMJ76+CRv
5fuV0TfxeoFensaJWwNby9daYmeoLOZUXZ5KXBIo/nIBMC3NYev/nl9PgPwkxJexrxPZjGd12gki
ZISC8KqUbFbTOUti1odbyjYsiwMyhlUWFlmzNHz8IpMs6KUO089D0qTDW8D/nwMFYlsW5qvSBAcP
md3ekUaxs3+NDHR5woIwpkljAUBnd31O6E4UjMERP7RFmolzziufOTivRxTBzID5pBnNw2QMy4Uf
bfiWJdcFauFNON9Bqkhc2ajo/1wBQt17PH80Rdwu22pMVHOh/vLwIu0VUB9By8kpnX4KClbZUoku
PpEgFQNPjU4UwIzKGXwqoGsr579hdkN/LgGgC4NEBdk91Uifr/vSetsj5wL/kagpP9HtQ0BkeBVF
fRN6LoJku5Ld7ygganduO8sjXYTV8c1QlLwa2lmf+hHlNVzCPY7aoNncq1QV0Otj44nld890w5BT
gfQajPQ9tmPjLamJRxf2a0DBGdlT/q/xR9nBV2Mmk3dKiASkhpI5AF5Fd/B0Kiy100cvIhCg1dPs
YI5WYi8KG3GMDzuGOh4RNyCy5Ps+t/lwYkTMBopu5RrVAruhUw7WVzYRFR8d4NMJnrYDGXehXQLe
X8a7k7LVvcTk1i+55pAHZoHcu3SVEj3kDVBCQIzrtgMhFwgjqftNqqlNJ5OiBBl/V5V2i5QE4fXg
5KDfm2eq3XbcDbmufSoy/xAZXP4QzBSG3kuKVURgZOhVnHhcekhafCQU+6DBuAey8wKQYATTDWpZ
2VODwqkoG0tuFF2ToIqobHI5M2fiDJAZGoM+h2QFDIzeSag2TDD5TFGbH1yE9S4ECZn7oDfkN+jI
Tg+gvxAbr/i1LzCw+6av4bHlkeZIjbpCBNJiC6/184sQrvnJyAVsnD4tyxvuJwQOE13weXkmuh41
dMThaNUJXRjNH2OzLTSLb6yZ4P8Qs5JY6m5HqIXbHEppfHtKgpqlrs6LwBW9c3R+XHF3K0G4Sq52
zjL+h9lhPehJ3U+W0AawVyAEKyHsydX/GmmP2qkoUrfEdjxX3rOyAMDlDZa4yhy1lkvYAQkouLIb
lkFu4BsjPqk30TwAQhrviccRcEc3OMdAq3BLo/SiV/dCr31PFAyxdeWcPgqTlajvNCGcnh/T+QLK
75YT0x+tnvf/4ZXiVXWS6bL+vIzkFGOFTgYWOoo+k4l3A9e2cj/5lc5b3IQ8aHr+cepOwHjzApvE
/iwGkPFFnmHWQVZ8wYae2nrh2TbEPoaH09OU4hWfQUMOjdbxxseOb70ayk+8g4C5y0YroZ5OKTtm
oDajwOJnr+sugxf0r8AMNW5luoDktTD/yOvUBzgWiAfvv+SHtsF3PoiJuZ1Iy2QbXBc4p1JZ8Z6u
pXNMn3QeUn1q9TEKfnBwVByA2MDKyhvwC5yb55UlEgV6CXg+U/ATt+SYjwRiokGSsB32srxNIgsh
9XEuCPKDjmwmCxnmxZCqupQVTZXJNvi/RmGpMRu0DQd8KQ4ToGilvXNK6DtAq+TcZu9Dn6Sbzf6a
bzCq52t40Z3LGNbKwt32zbkT3AmrY6/jK6Vh0jIHP5Cf7Yslx8KXPUSCRcu6j1pbTKJGDOexdgoI
fiheRAhJ+WzYlzEi/rrmkoxNqoOEMqOIwQvhcs/LHQ2a+Jn56OF7a6FS7OdeuAfT0sk1363IUbDb
W1KYwiexKtA36MSZtoEmWMKBljee+Ofdaq3pTAlcwSIXMLJ4FKeHJ4JDlQummtpf9b3JXYLFEMcg
x2PnQF/IOjjkJFGfsrWcEYoh0IRYFuKsnc8vRyO/VM0fFsAmhh/I1lmVfAOrlwSUHayJdVPokC1d
haceNelAKJzYYKrNCnnhsf5ATEQx/Mk/q/rDg+Z1XW3bCcEMT1gus2fq4dmdx3DmwrJYnmUJL8d/
onKRLWkUN7VOQ0anXcNIhBMbnvAWPGPxYPBfjD3skytUSeXCXJLe1zf9PpnydIhy2VKUSCg0cgqe
FU/FtOqUDWIq1BojCkwWN+Jo+d9samZGM1PkTKhmaOdu9/7MmKTzRLEnRMqMzQYUsdO5p+jplUgI
bLJXyRwo4esXgBvmjxqxIokqpB9ITZhIzsYafwQR3i59l0le1bx1BXsVnBpBcvyGDyBvtt289PQl
OS5pzOkENFF5fwOKqQuvM+gbnoibke5LmwJCaOyvWdHsKTqxI0UZ3UpQnbZWrYD/E8ojkzhESWkP
jDyb0OMidnQs37DU0qwhoS884Iz15pA+9gvJlWhPJmJfzRD0KctqF8Wo1NOOUFJkQbz3C5wX/CMk
bV1ZSE/pKGGV6/4cACMlEnTYw0XC3rg7WFzQAe34X47B0otiOWXDmMZxgCM76y1U6b1UMpPPCE9z
N+4IPBifQBUEelGR5Dlrq237AdFMGKE+CbNLenFAei02nWOKWiw6+CWjTQpwxwEFQ+l1Va+C4vqM
YosaP19yxJKg5bEmpQSqU2u97ux/9YFQo0bn9slsPwH2jGrDGA+SxgbCD3TNwqh6nNPDGM0VZbFP
TjJVRvJ1uxV0OqNQ0Ai5L2gFSjdtbcZgzcvw8eDeQrFGEa+RfpyzrbOBLEE8xz00TaKNvXMo95K3
5MUg73O16DrxB0vJbFrFQFi5ELafEdPrOElNtwBLFiWQur63UYkuNc2iH4vNk4fYslGN3nmhsro/
8a59GMjwVUlshk9BMd7XJWjOOoSVpNzkQ1ivoBsMGvubLFZrgsVw1K3CQdF168d5QQcNttamp90k
BTG3BH6+gEC3bVQoSmosSGvqz3OQ17ZLYcNNXkuTIyRZqmaU6GLSDZdBFZb8crFefD2QFhQLFovS
bV+lnt6tu2LOtiUdV1nFBmCNufDlxa+zACfvsXLvrindZMbhtVZtjICfBRmMmrNjP85sNQPLBbGs
oPHUpDoUxFeP3VcV+NQ6r3GYOBCDJ0I5RIP4r19eUNxfCwT53yyikh8y744a6zt8od02yTC5ZU2Q
zTbEogoIqityoL0EiPv5N1bvzx1tsr9cTVjvbic9YL+iKT2E3XUF8Ol3/D2rj2M3+/Xi9rIOeOqe
PoRo2yvkUQ/NrLaPPQ7Ga905FXMfY/N7we9T+8WlyoNDyqtvO2vaHitEDiqdDjGcMb2fXxb2hXd/
p9IpJNO6OheJAcKpaY9Un3Nk0BJYatvVjZDOXDasRAbzTP6ClDkOCLPGIVf+6YCKZV5rMZLKXt6u
LM93O/pPCoMrE2soF6xNwByuTIBmQkzScn1O66qJSkNLQ/v6YMAml6RDREhiCGjlKWRhvOX3W8wJ
Al1PnXFYdA58KY3XiMNBnCISFlFhfjamGSlQqH5dJWvgwt2Il7RGeXLGE5hP3xxyKzFyB3DALBQr
TrC3QLYHgIgbCz0C4DNFqQujeFf8avL8j2ZYM5NSNTz0HRA2Arg0CZmfVnxhGjC6xB0ab1hW17VK
QQDFjfZCQLJoYpS4nEc4nSbs9G8jyQL8Y3flNWK7pndMbUoNQQ1x15+ZXE1Xne2N6CIwQ3kso03i
QJMcfdUz4awN5dX2Y1Adm/yry83NocJSEEqr7w3GvT5ZNqfzvcyLhKP7bNeXFxSA1smNrlG2Bt2b
Pbn64N+D+vERPrz8CKXqlFO1wxlwqSCZ/W6nxduksPvMGvEQy2zqX4il8E41yU+WL/6iaKr91jEf
ahD5jSNmQL4AkJYO4JoDrTCHGlPPMX1EO6/xXeXxLqkAWuUq5tlnufXKsEiO0uvzs+uQTfDls4iS
qQixjujZJkFDy6pS6pw0WU6GW9B9b4hMX99wCAovlvhmJDpTummVU0M1dRK9X5I7f8ek3hrrqlGh
jP1sQ/GguaRooffWR7X7XBg2nAwSLGjvShPDIRLVVToYZGKKD1t18Cce3vKvUY1Yi7MimJippOEQ
AgPD9y4kFtpiqEZj2mlHqY3hPH7cWrTY1v3pb7XpISlEVbOUkkkl7tgfdkO//nRgXKKxbFLGqZD5
aPVzLfiyyZiAqi3E+Vl6NkvPO1ozGvVigp5UpNmsq6o9+fo8yNSzA/fMJqGtEwNdTQAxv7Rpplp6
TYxJqP+g/GvOrBisNGr3yjD5LZr5qtM9Q+WMoBoaGWAgf0gd44dd7cz+Vy4J8O0M1cEYmAyWdwOB
E/WEi7bmFRzIeNIB14MB6ii3jGaSyri/2QzNFQaImzViMYdS6ZmbR+H2c8C/dHcI+kMZvf+Qml4Q
M4PMgPAThYHuYBb4BoOLLBbov67fBusAzfAUCebeobAx/xxeJqV3k6W8h6uNLzUGD0dyQ+mBXE5v
ybP/ppFiLeZ88DVYV1xGTh2mlPDhgnKHxOHgtM1ciLmEIsflaJydx10gcjYuDrPD643j7c5UqQw2
uw4+jrZA9S32ZCDif2RKBjZVMCPT9v0C9+msLCK1REnSnwoMIIfMstOCP0OLygEZu1Ftm0kQ/ZW0
TSFmaBlY/SCHGl/RLeR+NeAX3qn1s3AhnGF7NM4J6grSzaDBy5ZxjUXeLlV0Ad9FJW++gdMoS2Sb
xgGCPVQsSQoc3bL3DIDkJ2zJBofPs6Uid5s6TqKIafshLgbzCctea9yYNtKXhJNuTYqOW2SBJawy
eSqpfHXzYpBjVy6dc/Rl3b6oNu8kOownAnqc4RIzhGF52Y1JbfObgnesxKUAyeCkjClXHHBbj8/Y
HEQNPFVQn7/ctIUKpKsBJ5VRaaoqLNmIvZlQPOvvan1HNfgghqjhMOiDEB/ZiX0w/AdsK/Rrl5UI
xl84ElgKepnsEzVPjckH6sRcYMegadkPQeoyQP4gM5/lvxo2XZrwyaB9O8g+7uNeWsG5lb6RFiFG
x3X/G2s8hRgmCMO2bKDurujMsEXRkzFEnrf49wXIjmKMisuqcaTwD4Czd7GpezQVpFVwX9mgLCP3
Jh9MjgPox8bub1uMS8ZtbGR2h2rcyaFoS1EREKa58bGv5TcxYYbFuskhaq7HSiYyb/zdH/iDB51n
w7/WluCXei7bZc4vh7zqgeiWg91f/SIthHPpX4pbnp6y6mr+TNp2KAxu535FrYvuf35swgSq1RvO
yAKqF5qyIu6G1J9ZaCACOT+qbDjFzrMwYV1KadXRGGlJRzIkxcVeM7FbF1hm+YrNLsZcr2pAwf4x
u3oy3kjuGcbyuXlMwysexIGv+JPeLncECIk5haPlB8SaahMqGt2qR3Bd2uBIY57+mhByciSCB0io
xSqsbJNe6pI1S3lxqTH705dEzrbifJfOIwGpqp7/QNtzD/B95lke6NiXOCQx4ECWAUxI7H6b1Upc
+YTgvgjcRW+VTLbp4kau62e9Vhs6q+9+aK1+f03bq5H9IhkisJYK/L6yXaqXfSKSKug295GG/BXF
EkfCY4YSVU+i6+C2SNL1pRrV20LzHarRul31B1PAACVmUji5ouC3KDk2V4rzMhIJL8nqm3/3MVq9
t19ZUvpbHBi+iZcvRwIgZoMiX8tJAtVezqsWlJExdEUC8QSCNPhlNTnVtkaTjE5sg/PUL+QwL3lq
o0vsxJsf+aol8n25LiaCct3GUcK3K86sPH2hGiDR4Jc5+ibErZBHNn4gfWtvCCGTYFoC+nFOFH6X
LB5fPyVvw+7xZnFkxGneGjKRi2JPg7e0ynkCGJbt0N6nMNSYleAlDUI9kQ6bRz7z96rgbM9KeMpe
vgSbTPBE544sAxpusxpByK/JN4rxNzW+lweLrI0CB0M8qoKR9IBiaVnSzTm9WdtD9OUQiH57bUrB
5Ga7aAawXftDO7kxGSW5Hq9Pc6JULczvShDZ2SVvyCtaamwjcxaVJDx8T8OdWRwO+SxBKH28Db66
IbxDte9VH8ta5eny5kGViowPa3sweWyDEwHyo6LT+iZ65gcaCg3u7O01MwUuoRvI3WZMngBtHhmM
y75VPiEWzVsa6rI0F+bTtmyZwXOuiLPsyGPIbFEcZKB2bi9dlFruJYLieXHirRCNFv5LUmu8uCXN
piNcWXYSIyfix8KMs86SwU7Tr8LNLXzTiFNu48JNBdWA142pZtT0Fillhfv/aje3/C0Db7BGZbWH
WPpQ+N07H88GPP0O3y0I3MMhQ4FAzBsDGaqIiIHQrcl3qt9V7DgkfFgYbguWUx0exxeDZ5zJri/G
6VVACOmel82SmMI6/2XkjdDQaJt4JfbXXMW/xef1s+ddnX4wYgcSnOL6dhmQ+zOj26pebWpsDuxd
M5oiAPKEg4cDc6jWNLQ8JW74HjSoS+J4APkPeVKV5IzvuAmF6Xs3sA2Eg2AvbnOYrgdb/reMsdlF
6sh6yf0NCnR+KZ5wzQQRULD2pVc8ihpaDR8q/JBbBpBPHKcFtiDsumyp9rgl1xf7uiDL/DN/SXUI
j3Ko1eAeAmjrR6AyNCgLi7klBz+kOQyVUMdDNaUWzrA+ygKdfiNDQ8dRtVKrK7aRuuTi4I9OypeO
IhvBTMNb+w4LCAnEIRyQFAGz+v2CiozPrESbTBNycTIWSEv9Kq3Enr4Ztw4v4Cax7WkRACkxL+ly
6JRTXWOswl/ii9BUHFEN1aNOoBtw+Ne/n9wagwCb+qUqwXaxsXkRNzyBdCKIHyqpeo83vf5v7Cll
GSEilzm+2VrVCiRNZX4C/jSLXgRzOIC/zNBb54aT+9MhXOQdOmo3V6vCwrxOq+7ruxxk9mVqkhoQ
EvSf9MXeXTmgAvGJXzNjoRAhs2erRoenheIvcQbi/ASc3fXN0FybylEiZEpEgPExQqYgw5VUwnRk
X2OmJInefX00GTLooN5w6pWvXd9oBXYGTbKsNenoTQ0wYOGMtDbXeVhLblgYQyafmFuyPgvlnzKG
iEKucWPKJc3p6GRfa61EcZ9H1BqQaTr5GyyT9N0FKn6C7iMZLG1B+Xbe1IAXOp2TxTLt4L5aTWS2
gK/v/3FE57f4Z0JYeE8G1/OpJjg68PunRJ/3mJjbWE4gogkuLP3pDoR1UTHoiiHIBAKDjMntIsny
n8ziFVjFqVAwwIuRfIgrF2GTwyQnpTZz9oFuPEIZYwsVNIHf+zjZdQf55MOjDxJDHcAyWWN5Cy7u
esWKmidgn9FOsk6v5iBzxd3MiBFVyEs8H7Vx78GzBgil08OjwXdKDtpX6MY5ckvceHoS31UqAdM1
QDhgFpLiru/+u1DHpCUrk6OqXSNI9GtL9ALra7uUo/oVjhxvuYJzk4EIU/ZKcIQRCSagRZdWUDcH
3VhU5kdfFHUEHYXYaOgRiXLH0KnRMQhdzNRpepXwn0yoE9F9nIkdPa8KYL5Bcqp8LINKZqU/WWp6
iLDak/m1NytbZtRsE8PwlbaHFq0lQUMTALSIyDLwleMonGl6wlNgmlBgEP5jtEKCOdCJguqZm61d
jBzePTc/37IVhcmrZOU/8X71/0R/nd/isgLCg9B5TCy4VmASjRhATWyFgWhhc116x+YOjzvR8zJu
Ile9IN935F5SSTJXWpuM9z9ErzNXZNLXT3h7tUHZ7Ct1RMmF/HABiPS94vqmWc2E53y4VeSNtGRe
wn2Tppd/hDoSSnV4gUBOlrA16Qnszd2sy2/SLRsbe2kX7Ad1tvXx3mjWT7ZBKZTTrZBhvMTuAbqN
e6OdHdgTBGzfy0l4kd34sOX7NabguNSKIcMlwdgvzUX29J3gP4S8alX2FL4OvnmO/V/KFhBeRoat
ztm0R9c0eji4eNjaD0AVMyeoZgsEJobBV//8tD6NrUtToFdeWRDZRHF3moZqcnW9CyiIlwxglgGx
LkpMyFyIsA23GFxAgraQG+n+mfUkDxSIlCwvKvRl2bU88ND2iaFpw2pj3SwOA/sfOoRtwU5LaLi8
BYC5ntBj4xhz+Hha+93+YgWsuprKe6S36pAoUxFMeiG2PrtpggZGPz1RNhCb9QRaHiUB9qaJb5TP
xyXP6Z9jFFwq0tlfhRc+CYQIZcY8dWoqDhDqTrnovuSX1KoUXXfXIkoyxOKgav6dOZtHz3IoxdtF
qvDIkBQE04wiXykKmsgaFOsK+f0uVxL7fXWX7OkdTDD3+4DZ6D7FPVbp5nLhWoSohH70mBCu6Shb
mRI/ooD6FtzRTF3tPht2Ttyv4fFKABA1qUAmd311LI/MpU3GN36ttcGS4qIpTNmDwCwoQF/ZTpgO
jvuUuMG/5R9Wtwm45AzHmIi6iDnjw+JrzKP4N8eaUrol49MZtC5tSveN9BCQGz8+HUDgeTB1fuvR
wuMSN7+0B+s4poaKZmn47oSDwCiqtMIFvDd6O/hD68sxK174e9xBWOUkllWbv0yLXc3KDPbefW0b
nFRIwZi3gZgHcpB5RszaUeM5ySUKOaJH3SBrptQyu8wnfnmzcOamZdhL4RdEdvPrR2OWf5K884sY
MVGRfUkUWlxj+VYdO3r2GoUw8AIHx8jnkdSTJbXu+SzOBuK1cOJk6Li/dBwZRiYwt0kwDfUY/jPR
cf1NCdzgXQ27XGtLHK4cMR7OBMw/CJKoxEvd1NdGCf5wS5p7fQkLVu3bGWuXJR9RlOasBKg2rvjh
TIC2szEtYSk8LSF7gm9cec/EYqYlf6PCBa8nN8e5t0gp5iAjjjpuLqZUdlFmUX5knh4y1Dx875Bp
i0i2DJlU6G+tBuI0idI0O2rS3Rzg1dsiLrrtrLzetrWY/rj7xCwSnAeglxA9LKOLy2L1I9CCDEz3
qOjXY5ZugNh/gAYh3zLrFsGC09UdkdPZ1e9Gl2/TNxpor6cSGQAv9eoxGxE1Yap4hNB/Ph1hPkm5
vkN2YAgD4OC6RIxN6JOTdvIskh7+yhBfTvVqj+WElsUjhJJO2tgW/8lNyM+TG2WmecRhG0PxObXz
GbBx7KaUo1/pTggV5FjRZJu+iJcMR3JDGsL+imv/JqfbZn35mypOCDvXBpNkIlIvU9rzuEI/PDHq
SzaHeRFQhsoYh7m7m33PFxsG5d4TdnYBCX7g6H4coMOfYH5rMD05Wfeevo9RZOeq7OwONPKwTN+j
K6l47/nnY6G/4tIOHwyCy84KV17/VU6W1sHftHmdy4aKxVNLjI4MxVNnkDg3LwD+H6VQxMEvPzPa
B+01r614lNhX6RsSUvJxWOuVoAGjfmpULhaLGkE0HZKbYd4F7HsE/AZORqyMDJHeEq1sN9PYKbKw
4eCFpU4gTHdz1eNn5nT50061WWZdS0oqwIObxOrEi+Mdbmyj3zG/rTztOD5ENcBxd//8ND4/0ANO
x1bRrZA8LFZOrfgx300HuT9RkACS7/94K0KvVMWH5r7nPkfWoFDzAMWXyTQPgmQ3en33ksIezh0R
0ZLhbO2KIMqOukN4FgehKHOpcr4qFy4EYxenaent5JJJtyMsT7BanuvlYBNZUC9CY9mnj+9mftHf
ExFJa+21BYmzT9nPidPGP+1kwpHHmEY30dOTqLoCMRlUizhFMPwOvE3QIV/MVzQs7Gaa8l6im2Ts
J8v+WQYKqPoP1K+sLs404M9U/Ry19BxP+Ja5b55Pdq1QE9eDzRotttNyQgpTlN4LFPSsUPlIG52f
H1SOzRXvfgU/vhFP252uG7KVri0wgKjkzQ1Z4zWKf+vqjkySgs2f8KjJPGiokoMyTyRBdTTsu4Fo
2ap7nhydokt4P90HXaOnzngAifxkNNvbdeqVVxWljA8PhjDwZY5A0Cp20QBWc4CNSE3K/xCSvWXA
3Ggxacz4QlNBN7W3+RcD6YHNwGRhz+R8kzaJMPABHRURoLuqQkwmvj1NtpZjE1hBpEEb7P2xjj3k
jRN/4NyKCwLkUEzdJTEQ0IjdGj/0VpvNIVT8oPxflYx6p3TWEyx+pxq5UKFB5Z8oGGCZz0MDXPa2
9uR449icBvWQPAjZbIQgaMpCiZaPAmETeTNvLAhGfOZZy6+eF+yHjwSLfQIe3M0Ul4yAam3UOsfg
e2RYwYCNer6MkEHgOzO+vpfka2eVxlt2fv5O14/swCddbjgWFonjB9zy/HVa8O9Ulf7AyrVWCsOF
wU7lQFcI3DZhBW7/I1tHTnSQP6x2X8D7XCSmxK9jVb97sMYqLAPk7gBYpCKcq1mXs8TUSoJoYg1d
hQDxHTV7cRqy97zRSnGsXRhgZOLWnNnI0WMPNFIPX7w2Jd8mTB4tK6hp9sCoVsXp3GSl0eZ7aJZD
/7Pd0y5Mf3UoN2Rq6KflvHlBIuGDzzVm3DRRzmLuTwFDCtO/EmWghFxEwQsoPnglzCGJK1Fx0a6i
N88aJcqbjZhh5u1YrOKxD1Y/D3ISahCWwanG0DfVnzIoP/2bgxT9WAYxqaZfqSwrWrr24NxRRhSf
3p9sL9RCwyRoMfZgIDeNKv4a4sRB8vJOmoZ6hKq2yOND51ZhxNO10tDBjD6DodkePXqg72K9KZp+
ToH3TNny/MvU9gp3vKGtN/8TamLuQ1pd2aHtYi8JitAr7U9yPkJIHw3JS5265XqA35jvSGj/AhIE
csOJvHJBBG+Qc+MR+7AO6IcE5ZU02pMFPpgRb1Di6TJxqvv4EJjHepCZsmVSLGdf19TMsdIMWvID
oXO/O1vpLVutCuCG471aaJozWeiqNwT3LHuzjEQxNwTdJ8rlJhCxjPfbwfdQc2c35qegWr1+Lj5U
0VtUXaBCaxPMlhTfgMXIrs+saLHC4k71RdERNllMBaQMRwzDBy6KM7tOrXJKb1xW9G7Ns0m7icnR
9aAEBslFjn/CougRFtTN5L2xmtOEN9/I5kRKWhA3OTES+dFQ/EIpBPrfoXLyNowTNS6NuKxr3S9S
Y2CFtLcyExB0ZO0vHlxHuZQkw0UFWFIJ/2Ytg3zRuHMAF3+scBuols6/0lhPq9wDJ5iILVFb/dXC
dKTL/yB30lIp5scv41KO/iOEPolyFBxCTaVCakA4VUJrsBdOhs2B9r0yYI/YY3O/21kZVig2+Y/O
vRLrtdTlWR0jUSA+2OpTgztHBGmYcQAaY0y77GFdVwoeQt9/L0NS5FcFtd+fSJGi4d4rGvbxbSty
0SFxfyqX+XOR+eDYW6NzB2arm3eOwGObgDmhfgs0uuE+edxWmVgF0EkaOWjq3snffRc7Suk9hXfQ
T2loyz62g2G+iJWnq/8QQfM7cjY65RB1ACbsLfVQmBF1EnDTnB8Z7onZeI79dzmvprZ1O6rvl4/z
53SwEhYZ7JMYhu6jW+6eOZBYI5iW5IX7rFpbZBHzp+5/4xuTal/WQY88HcVdQlaVcPPqdmXznD+s
PsTbu5HQQtopug3bI7zDdp6nJeHp3ibcSKgIo1StE34CfotLv8CuYvdCUDUO4ijZLdiR2iG/cdC3
pzVqoUl+14QScNKwZxjkYOH1DgSwNUuLUOpeXTVkHTiiH9RU9cWn8boSCojWEqJzZty2tedBJbjg
L2OLYbAhuV39lAO3gTNmf/ySemr6ntvTlxz/V7UZ1OMjGJ9uGmQXRhkJx7ugFkj4Th3wzKQSzQO2
xSeN4ibvb23hxVJ3Vg8BoOqlHQCe2vT6m53SbXuIihBoL2YGpO/T36PVBGKgetFfRypsCUhCzIa2
uxIjbEL8RWBRrtN/emqHZ8dbmRV2HqRzJ22XxZdMnf/haDBlEO2+GdI+IWH7FXNyf+FMpbIhFFvF
LY49KLMb11+VwjKUnabSmmeR+auW35tCleCgmt2ZzuY+Ln2DM0QxC7+pFMyql160Udh7MAGtu/o+
xtcSjF1hjHRAvdf7Cn3L6NO3TubU/IWj807owkE4J2wgYXw2zPbGZsv7irpPjs2lEALxtTEHOcfz
C/kGKZ3VlXoma4lA8ae0wiWpHMovqoAH/lDa/6rhu/lO4EHo58GLYLL5I4Ghgv0a/lz8Z5ZyEMc6
xj8kXykSr7DoAzFnfjSZNxAvLxe7LG7D90D76Z6S3MWmGfvY/xaDSmiJZaMPWcwzuNBx0BT3i1eW
aiDVw+uORV8v8o2tq0wVAADCjzT7mDzMfMLa3E/oieIvwWMrWl57Pz1tBH4If+67VkKElE89Kfg1
u5abyE6i5X+iIrqNn+vLudMKeVN0ze487Z2xhXYwJd0HmKK2hjyfmMpLvnMDIIJld6PZbDaGSu0v
az7wH8fot4jQegCV5psmjt7WTtNTUkY/Xn6kbtOik2Jfu8GoVrxI7LYoojjUq41BMs/LuN3bjSEX
IgMzttbrFpc4jB0vT6efsh1tAaeAMUSsn+xaT2Yx4vE2tEfi2IsydOZl8FvgLGAyNOCtUyRAQGCn
MLDEUBvAZP/Kr7xK2JxrXPHrUxYmDMsgwdcx0sgYHHWZ/KnH7mPX2xY/Tl2dDg3QcOtGTj5pppsl
xp1vq4KOmBi7ufd2at4aaF6G/+Z60ku1IZgr5EVQgX739rG+JKBH4KB5vcATOi43O23YDlJ9bxKr
nJclYFD/NqSSsfpU1Cw4or1jUEdjB9gVzQyJlo4leZRsleYMHdCFm1mPnj9CiS+GycGQgcwm9hCF
zTCcLeA/8mS1Py4VqQzzOv/LvaUlp0uVhxCETwJEE21NZ+eYymRKF6MXDzvAiUV7saO9JGMothAX
YNk0OzdlA+wRLBR1db3moEYILuQ/23NsbwehTnA01C1iUO4Bgzh9DdCj9K+pDUgPqJAazqHde2Qu
shXesr1ybqt6pzh9Y3A+L75VFjEdt+oX2s2nZn2ypzg0hTDunbWHpynxJh+LH1xBMQR7wbIW1iBm
IfdP8GPBbAvTt7lshW/IZM7ZP8OAyA4EW1pH/oTRXA6mF4zJ7+Ws0VhebzHIY2/fIdFO8R25AHqM
LwplCQX12xYCLkNb9bCv6OdSlkWLnTONqCu82wO/4jLBOdFm7JSS6GWgYa0N7M4I2v+OBzEcDqkG
BR5wsFhlRp7cqUCY/NtZ+nyYq4gtRQoSuPlOJMPsuY+/VTeHBsQh7sIVcO3ExRHrcL98JMECf9+8
OxsZFejlh8V0DoMEERunDIlfZWCKmIXgdEORhNPECszhzSuLEFVwZ/oTNAZTIVa//+maTYVDKMn4
lm/V28xdvcaAh1any03Wv3bxQ8alpgYptkVJCSWeSKbEPmNhjAUn7hJ3VPem6hxpoUeF8zcdJm+i
5RtlEJdtUdC4OCy3Iz5kkreAxTyQbR1YB34Jl2l+YIJams6IYISA2Jhagg9IXk0pc8bhhjrhImF6
Thad4V6igjUgR5CMxT2f6IPyJNa+B7PpxLSiSX/lDMCA479sGPlzzXLc1xCWHAkw3nNUnoRAHLmE
Kz0CclFCTn+IxvfxX0EdTWXoXakO1TFKW7i29j+Xa1OynrOd/3PoPXO/qzDYqwXQg6aIWp8oqtzH
fXz4guY6PuOGxny+30wzsEyDpo8yp+U3K+o7vFaZBAuHrLrlGbDLDFCtMr5vbm/ankPX57x51ck/
e0eX0LI6HAnN+aP+DZLsgndF3XZGikGLF47jI8PQ/bH3M7vchhKXoNzg3alCI6fEiAA+u5NWzpai
cmFPPsCnd4kVzfc+/LXwKBczJxCa46oQK8mNgWvQKKRltAHWxcNJAWSwPDFmXPvTzgU1pdpllz+0
OPWR+TKkOejtor+/evatmA8G5l8LlCAriAAgNnZNFeaUNuWBwp8h4loqsJkINGe+FgfuEvrZMtFV
KwZNsFnStRg6hLnTFS/LVycHmqVDDN6qqTze1veAaQ4wbuwUp21ECjYm8UALjMcxMlNsxsSP1WLd
XoQeC1e4pZiCc5Gc6YjKNBMjrPnKWZd3wQbxVmya/2S7lkUvmgy6ccwX2wmgsbhZssUOhiaBJXBW
UOO5xXI49R1C0YHUufGihvRluXEoB50TEUYkn2AT7sk5AFJS9JIOhHwPiWhmycJikV0v9uxd0tVe
8csNzhSOtrSKlh8lDp0Qi1hq/DUgRegGb7OYL10pxKy/jbMKChWf3WV7OSMQ+dCGPPJ2EJSEH9Pc
Uvsx8cVCf3p2qDPZkWyTm5qKuYKdSxiKuKzPIxFCxUoTfWIJKNoPqZ5DsvgTVms5Jm+ZtHJ5KZGl
xxQUQHPjcOghQvtMs7rT1gvQPzyi5FGnDZHtZA6r961cPh09M0XcnKDGo/Dvy7H/qZRvWKRI2Izz
EbXQHRSH3jJfAcjxLrQ3m5HDojgVkQgDmadUEibLCW4k5wl3eVtvyP/S/dD9VilncHuTHfz3ZrJ5
bIcaoF655MA7KjHcYUSQmUe5+rwXAQfUfuyC6esTgoKHfGM7oVBr+yhqRe3/N9rsKozm2bIfQfNv
BXiup4IVdiwPvyD9s6DUMvq+dwQzLIHfXQguVwISHE/BKtXIis4nkhzhRXmNaPHBfFi5d0Tf2hj7
PW6KFxKQRNHkplpJcKHdGGxc/dEGs+3r+bOlI0a4auGjNl1SYPkkzk2mUfvF7xY7XYO3S/3WI0sL
TDFGhMdlzn3RNH9pD2JJpbVbKzMEE38tKugAG2SBiy35xWX0Y8v5Scc2/UgHXrUnK+lC5kgUdXxL
IWOEey5SZHVixXwi0obz34yLMDcqSvx8+iFd8p00sm0E1uPcQbuZIYHWM6ynBHUfnxn5rVnhNRuJ
yl/kY2v7Wki7SnEIsPiHyLsFUVdxutZoB+yKEeAKwFf3yrc5x5URBAriiM7JDn/2mvV9dJcRT7Ut
q4kRD/zdMFKmrBR8kJsoaqiRIjHHcoRYUxq5ryYlY0EWpIE03svK3m5Ixu9fGtIlCNq3m5RLuXCr
3Cl7LKOERugkssqY0MbJcMlkgEMUPFmfPKdmmPduE9YKcTqOsWB2GpwQry8Gg78BdC/3Wp3aQwnp
Fuy6Tr8a4WQMy8QWv+atectFrg0glJGKN+/9ZbvTgWkQPvN9x97gUCDE/G8xhzRqZQ3OSittu5wi
NfF9ddLVfAKobQaB0yhfE/WBkKuN++RfU9Z7G0JH6K/dfy6BM5X4jMsS9iLQf46rTcUtJINl1OTg
j1ZMumQAT8dY9IvQleaCt6khPWTiuwPkCSLKIzCLWx2f88Wjf69Q2WP2i/nuB0/XrkWvL7RV/8F/
3v50O8vwoHcJwtTK7sPjbKZUF4cK74Jq+BYTHbLKT48dcJ3siuFM/DszEOCvezvXZKP4B9934GLn
mY828afOK1ji4B3gLIk/p1/N6fpY8KNko7AEWq2DCgfBAXT5UkQkuZWCfF+EE3q7I9XlViGW/cO0
RO3G/Z1jHFTDgg8I8LoBjn0uZQjUDwCsRjWjHDlFdQhLOQZtCe7AG0raWaGQGWww+gvZDcY/gnc3
AXxsKE2DPbkwG6XdAAqLL+o//vyxTW1YWI4HVaGjpcn2+by6TiAlEysIuXt1YpcJ/UJ+OgYKLaov
r77JYFRXr8VJ59fQr+kOCswuDdLVTJM7Bo52Zdz0GrmI5khkAB1Fsx3b3CphlgCMnzXEShNE1nrs
g//UD3GwXE6Rl3UN8i96XYalopKtJtI0WA6IBB7Lo8dvVxsQ2OfD4w6Bf4gdktnnybiopqoGdXAM
1RdfyOu+ElCcHf70fR5DLeH2FaLAcnZZGkBMjiv+9+JDvDVJBQ6EYp0wOiRo1iwRbR0k/BrflJlX
wYhcT17nG5dbSQN/As1maDaxzUwk34I2aS4Cjo//TJXP7ZyMP1tu92MIl2h8HhllzPTO0jiVxlaP
eVSzdhjCVUvlyvy7vhLqHt4dlw4TY1zATTuwXGN0GL21EzVpoDwt+9zCWN1CWJ0ECqtwi/ncozLQ
GeR2FFN6h47fJn8N1qtmVs/AKbn+7Are88U5a05ZXFFYTKG1Zg1hcQc6igR/IOJ6I5JxBlNkRABF
YTrIofGvWN54DvWuGqQj2pu+KG2nAhBtJEPDtBJB5vwgpZFvQh+u7kBu6uLtBCv8z3h+lC8Nt9N0
JgPdclU2LHYTrkohJnANIB7A9xody1+HH6yIqOsxeMklsKXBjukBqgMZY/DoyRo6rs+aXF2lNIhv
oO2cGGPqbOfWtuqNgrHrAUZX6Iir8sahUTQu3ipeMM2s6M/87jiWS6IkULYDzQIsELW+aq6oLZXv
URsnh0qHhJrPyY4hrvxAtpylfBz+l/7BWV/OSKBgePpiLIXRZW0WBGhHeFRwp5U/VlGLJcvXZC/D
gAb17ViBCNJrjd8amvp3mlKv1kMzni3CPlSZkKyALzxLUMv4b2ln0hTaxkiur2f5/pBHRjP06VAq
cXJ9YF8c5FRJ4XkRSp4v5cTnW52txRPHGiFGlykZE6zyfObCjqY8rdPNisoLOGkWJCUqAziB8Lrm
yAZoKPGjcH9MwsLuIYnOVTreUKXTjtL6RjQkosnnFgfEcmCWhxxCLsAOLz6064ZnK8eLiK3QzGtb
CkNQb/8i2vFnbwLefVYzFcgmiFjbrOO3r5R9ZRwWVDMiq3fYduvKwj+V/4ZnE90J4m/xkETifNXo
VAIZBMnunOKPW0LrCc0bpXmpzkd8PnUWSHZ3GKasN6aHWWge9ssvNG15NF/TSdLr7InhqbT/VBcr
7eRoTeWuLnxIW4wHYc6ksVgeG3nlzvBy+B9Ei9afLKTQ4h5sXYmDC3oD46oD+KBISPb+0O8/2IIB
fz1rGW4A3qIOU5NLqYP/fI3yYd/1Q13JMgaXXIz0RTeN9yzzy8jFDJQfEB9krb9oNoXHtGEOxUzQ
PBA2ZZyEd18wOp5befvKCDAkUhuTa7h/rHAnEAksvPVYK2bkkarDe7lWqhR1Dv9A7cbkzN+/ZhGD
H9xbOtiR71pbD2VFld4p2HH/uDsCdjqpf5vtVIgN8b6IHN4pGjCkN3aWkrLSWa0s73RDWILHHmDE
//ImOl5rx3nLgSQa3pFvJvnziMZMw6iC2DNIpXq8UzEknHEcNFHsNV0PLn6KE/zBdo6a/ybTZFyc
Hwdeks/yuo+8eTRyRcIIg6QPcDHCu8IG3ZwulD54662WVPf8BCXaOWXKm2mFhl4dCocFUu4EycZv
faFpKfhN+fS1dsaa5iNPrjKdumQ294OVWALt6Zp/MnCv9tLyj9OOunSYRaNVEkRvJjz0/LoOfzHB
8X7c1tRN51l5YGYHWDgLKIXzKgMqWG7XmxG1wVK3BcY4nuBSYLJNyWluTyIyyVNgopo2DPUEp+Hr
Qi46uJQWdat0ZXalSLp7LqpwbiwUfGGdvHGAN6POxnXrTuNjJBwdp5P0eos/Q7qnPulDqav7/cUD
JygGpURjinsEMbNTYirsoDf6m5WdSPRFgo7cdQQgTfVcBvPzLgLcZseKqXU2mGP/l5NOjG+t+O1W
cMbLB+TCgaLLw6zHrQcxLZVd5OPT07+iG/aeq+MPNogK/21r0kdKgsk3dpnMGQivP7YbNnJSzjei
PrSGQi1FDNrMf87W24F3N9VBdO9ZHaDnO8Lc9br5ojRWtHZ2kd8p73iDwYleHJYzwU37dbgsy0Lj
Z79lqFeT4CMqcODoi4PkhCw87bULRUV7IXm3I1WX7Ab5wjrZEatu7iizerwhFtYFftZEHHXHM9fL
VthDAZ8pluZrK9Ge+sklxiDPrN3F9DprkUhj+PA7haysB+a8qSVUVl0vxeWUyWOZf6wEvtkp0dDi
1L6kp1tQ5eYjHCqX8x5+kwSQBm7eB4bJ4ezSrWVtNA20T2x8zVNIECzJOEGQlUCvrHcBNc1s1yg5
GLk74xKkMvropqJ7VzBK6R+qvjDorgLzZ18FkE9HYwUHqxkPcWnnP2O/yh/DgYjiawrgZsdCEYXl
r3ASmsqaf5bpxTYn92s2jvPeKr4X8xpsNSXAj2z4zvmNxgSnESJaK77OqURN4mjA95zwy/k4A22p
kO65BJ46aGntvWLjQOZMab2JicsU+1j/mzDlLr2T7+Cr1NM/O2/yNZgFuJAT4Zh1En/FD1A8HXDA
phqa2+tZaEPhXssYGEvLWcuThSc/+BjDug1UUqiVahROlV+pUi6imrPwRe0U5D+Sp+mbxPPLVWMI
XZN/D/8AtJYJVw4+HDK9XaCCa/4wmHzP63krQICbfKctNvOebipM6KnWJAaiJEDhGjBg7B/n4hO0
CqA0GnFY8/tw/llLas3Chh3oi0/+KGlu2CgfKcVkhNqUmMNBMhTSh4q4Lq5c7Pw0rOU2UvGHxeDQ
ahhiAwnuih9rFQbboQbL6LBbxkW6ZyZgauLow9ktAZsT31DF9RJ1EU+1kLBtbIEA1u9Mumd6mxto
ThJyowogX7qzp9mSZwj9eHI2ZcORLc7gydtNpz2e3NB1M5YWaZcXpP2qTRlPvXA57E9thVUG7GGz
2bntHS4tE79ikiTfdyweX82OjqzcSZz+EPY5xiM8PvVime8JwjaGDWzW30FAIP60h4iEuNtSYMS7
K6x6jBxpLHj/LGQcnXAgd2e0oJODOc2L9+GB4+4PC4PgS3ySx202LVFy4YU0heCxwhthKgfog903
extaVDfybktHOVBrcdtt8l3EpxHKPfSj+OQoaYisMSJ3e7VmXb6TQzJsgDneriX2LT/JFSVS4GuN
avg+sKvWWJE3iZp92TdJlZf43GKhw4Ngf/XlWMYd6Ab5ctkNazhHgd254QhzJESpwWBVIc8M/IHa
HiqEaBxTsltLHJ7HaQ6ekQXcM7huekpWT/JDaJbhfLeqY87ffXsroURVB3zxHV4TwdWNgs4JnH1A
Id8ZYNkQV0rv9q4i3EKhnzBls6IHeokzLJLAC58DoYCuY1GXtaj4O9Z1P+P8K8R1R5Vo6LEA2BVw
2gz2kQwWoNYg8vdEyAatqCs9EQ15LTmGR7CwExcMasXq5LcWsr6NWdqlYDonOux1uwxESdAt8mK8
tsY3LtPUwbz6RT7qdMT2/IhSg3agWif1fbxW+pMd72pz3i8KIfO1SKM4IxkYNnafgT6RkY5+sl0j
S4USNVAdVBqoXNDyiCXronXwGtNpWDKAh5/y5pgcl4Acs6bc7Ygwixj0K2ctTv2rT/5Fj20SCGIR
2H9BtrrCrb9A2Iq0ThWN2x3d5NgYE3puD+p340by++eHXuVFHh2Gq7r0A1faKgWwrvphCXku8eJB
yqwwiTQVpkIQHxOniJA9YfUWCAHNhYgQs1EEtWH97ERh51dQZsX/pBrxuVg2UAbY2zLRmChUmKuW
CcWO2G2XbWyWmV97kp7KUjRL53I4ZmDpC/1MGmSMTpxDK1BjtzeDjkU2tCN1+v5Rrj0yWlm54+mE
yOfwDf25/zOBibYpefCcrwEJ9RiQJHByLpZmJaVs5XRzVp3FSuAXy6B/WOTh3VZeFpcSDUY8955/
0FlTzGLoQeYCEboKAHNNZKQAhBj0ZVdIU7r/MfX1WQuc0QuOOXsc85mO7ZCZBRY5LCLjfw5ZaMnK
/AvZBaju91AcU2sinvKyNAkNNvZqxWtErhfX3KU6yUHklKHeSE0DOKY/9r+V1kHK5f9VFUcw30lg
wF7O1WX3uZlTcDh2JEVvrsWjoFIBH8BIfjOZrs8AhtC2k+Z3eNNs5BIeQCFVkh7qSTKngGjOhxQm
SrCdt3lN6e19DXS1sOU6KSEuXcBHGRJckUqljpsviKaDyGrUQQSgWsWyxeIs72rzuDJG/uSfMNIT
iYhaRYwB+PsvfUqd++wrDE6Be+NyVqZUuUQr5cRU1eYIow7ztcYZsK0W++AOQnRbLmVtslSeqFKS
9ImQpYHE4s9adFnoDqdT8uo3u0PdXMIRSitc3TmWk/8dyR1Ws1tC2Wbb6iW0aaW/ftpqU5lkXJEx
52ZdT+AWJ6y5m9QxQczxmN7JU9pqLLTcrZuvAtB226qw0KYguXCTPnNnsxv/Bbc05wVk4hB+mRc1
aKkaNVuKrcoLtsl7ic7z5IVAFgvmwBkwc66ApSyO/MrfG4U+sUoictTGIIO3KWaey95ZWrh4aLmx
Bjije0O5MfdfpMF5tQ37CONsGDJOGovQZ2MkzmlA7gP9OF/HLG/2KIt/kMJ3KnCbGft02hbeoE6J
svcuc8lGbWWYgnGRMtCFuRXOfYeK7/gJop1y1vwdaIGpW0hbYjj1uaE4paWpCajsRA/M0/GU78u1
Qf888rcBroplS0UHcXpWXwiv0BqRMN72PWIBYYgETZ9uNHxaIOe0OGnE/ck7ssTc4m1exH9K7Z4A
QRmYoM+w58u+GYJfhdtGCaFbHDLcQUVFgQe5eO2jYrZWmqFNLh6tSoZs5cChb+kG58qqIBfrmM86
E2uQhsX6YvqK/Pmmt6yx6WfMlE9GXw6wRdOughFqXWJKoSA9Dz5iTY5B/yEtlatwguJ3t0/kgaP8
wNnzy+aUXFfzkM4o9lNPJJLcK1OUz5pDCCqSCnln6mo5Py59UtNGzKHtFRVArF1BG8w1XXUDi/fg
8JSKCp3S1ZWtwLLLF5g22aWhu1n9dlSPKqRVFUU5GvJ6NhHtcD3rXID8YqL02qTgTk6cje6oyxjx
lE/7ZEE6uzFKZiZJ3cZDcuLlV89o1ABFhgKKtNuEIPWtxL4EKXgs9AwNhAB9NZo4ZlAxDKxJB6PZ
BQIYfgdccq0tHmln+v9zOVR4LrgcDNnfZGtwlpcZh59xzN5MIATILtGhNtuHU51lWXMuPbL7UTfJ
YpnQHdVS/RieyAg2MvEzYCmst3S5y2ovjbwjwZF829u0xHwKvVv0lYKm+xo3+iEyk+u3CRST8TNh
VO4CRgUNKkpMn+ZLh0rcG45+7kcUex9LmD6jgjfSRchnP4kxX5vaJqgQjTbh0uJ2szV7YnupLY2W
EKMkJAYpCaS68FGfEnb1JRcWoFzvuu0t02wFwCY+7URE5UJ2+9lbSFSWuM77XnBzOzhSt1WSBoNe
W5VeRhoSkSOBCohveta6N9GpGjtm94nOOKBa98+TNAbVmtEk+oY533QrPNMyvL5FwKows2SSfYF+
bFGrVEY9+jlsq8sPGmFWlbnx1l0o+/TN6g/zZanOCXEj3IP/LSnF7StJTBMhTSFBgxjFanb5/MdD
psXLcs1hk6AVYu5QEI2lKsRjMMsy9umqZkI+q8MQThtFtygBJUP2hnL1h7StJE929Q1hYnVmEAKh
6JC2oUvoFXh+hMHPQm5vdS1aya7z5ZJ9cTLEA6CR3MaO2SpVHgeH+IlrlDZowjKWt4hjlb6JMVoF
F0TpSD0EBQq+S+Q7/zP1X60gduvynqmN2FnAoLYLHrJ3IGet37xMDbNtMQPBaveghNxiSejSf49e
JtC/rqruAUWj9iyyVidD1K/gH+PcPpXtD+Dx6QcYI5UNP5lmsjxZmWHD2dOScIN6DvJTQ6+Ua1yp
brveoWdSogUcN+iwU/gsht3OwGNbOtbsCSZO+ajKwW6wVJDf5DWD6FrkiJBSsREfRelkJ05mhjW+
ipEBM6Pbk4BXE8iNQk+wEEmq6pCaHmKEO8s7mGXKmLuMleQaUyeDbFszTBc4Iq5AYykhhUE4NbwV
pY48Hj3wPoOd/T7DaxSxlriDSEt90dQBa8YURXqZ+GQqLHb01e3fTdz3UkiT0G8bK882nuwmUS0a
wLo4DbYbT4g0FQSxyVH+uii1ScY3dN5zy+c4l3YveE2CljnKEAcziYdxy+zfqWCWFLJUzhXlXOk3
JXAHXs8bR21Np+r76Hi47iW+3OWPT4JbX4ahWfXs1ec44pjfUdywTsckOMurCXhhQ8PAQI0gxLoG
jdp+CJWFRdyHiqhl1FmTrEO7ZX6JMIDIUyg2MacIqGVcldoewSQp9/xjE5lQwDANsi6DfcQrjfNL
ANg/yYyFbCDjE4IVUNo87UC5U7V8JfNutWxPzn74bRzqYOBZbu5wgqc/anPy1I5bhR7RNpxHHoTS
lFU41z3Wr7hiP7XvuaB2yQfajOhLSVxi9ZZIaKyl/4wtQ4goX9XkwZ86FpgHgRBclTHYFLB20eJV
e7CEWyzjArkEOwlVtUV6MKuyFjCBEBecFFg6zLPUpQV2d3uMqEQdqNDFMHJsgkzLA1kIwlL4yaaD
Q1E65I4zgDYbom7u5yZGkrdLdMQLjxGlFaQ1J7D7PyXBOnONWj6jJrnWeT8teKBu9cajR9U8R9cT
0l7Ihjn05eaRvqT0GBtupPfpNe3iQocR1Vokpywgu6I6ljaNc/sQ8wRpMYRgKKcI7cqF7jBi2Xnh
k2wUGhWe9Y8dXbDOwiephnbm5BX5xhiHS0qVgBIyu8fKreE/SKeiR9Ph7YAv46YmKSPRLK5l9cxW
QmoFiGjWAFeRh38tWckJRGa6teTQuaTx6tqR/aL4XMlEY2Bk4itUqJaNnkq+4s5hUXp8iyo/tPV/
HYR3cwNqZu8foYOR0rCmfr6fl6OVNafLK/Wo3bZ+zvfHcaoob+PF8kus6mqHbXl9kkbO9e2NrEjw
+kfR7/e2jhuSP87DdQsTPpsMyM6IaDnhAY+wUfCPN4YCnjl47LDQsF2i0jQmUXRHnrhoZLB/aLv6
8NWFcmMbIelh1XozScJ16GkSjTyxcIUrlWwKFup1+DVrfmQDmKVhRO+ij2sntOnEhHQsLCpUabPu
92HbXG1j48WJLN2ZsfUZCVyPFsGbHGRxWrUZ+dTB5eEwuoOx1hwptGKUJpva6I6TBsCsUHFMBzYM
V3D1nS3WIrHGNu0iF42tNrNuccs/t9nDrBY0N5Q71fGenRm0kSqUPOeLMpWaCi76NwLqiXSJDvXM
XUZVitXbY78mPJ8fbqWTq+2/7HmXinCGuYlTNJAZOp3mtl+Ddz9YdrJrZ8Sln9eyp0jYNFTL7VMA
c0Mv0lcYiOH2dJ6fnbBlPwiP1cd6EyKl0MreWCkHXCfPEMKW3l9FGwDGVVddfqmejndJsBZyYvCY
iC3I2h5gcZRLBLKkj36epqPQx3lOjoDklmkMAslvr1moT1czDYKvLzr09/YHmcyhEMbg6q57u4YM
kGGe+FoBh11inPJo2rGOgxF0PeBCqCU+wKxnDJ+0L+Bv8FEyAUN3r/1tyeLK6X3f3Ppu7S5UyFrd
miUK6PMYrY44YomnQnxKNFRGr6/7YWH64Oq1tl1r76hIX7XBRkkpzhVmSeNGyVci7HA9cAETo2UE
IfroHq5Ikv4OziWSEITjVcLPN1tMgVHNAetn6N2dY1YpO0tunggnT6ghRgdTiFSbV0Fha23cdOQ3
Bhj4hAiIMJqeKkDzj6+Q8j2HorO4g7gpDFw+TyppKLMtQEzeiE34NajYZCHvJ/3N8/tCbPUanHWX
xqEUy9oAkN1op/WZf4ncyWT3pUSoC2hRgJG7JKoo5MQkUM9km5i3ier7F0k3+o0vH7IRZbx1Lgdh
EhvHCtrqf2evjgaSygYUfzt07hshlAQ21vo+s2cR0QYCE4w5qX8Y9ncjwtGAfuL6yE1f52EWxJbK
Rt9LDANt6732aW1rrz/jlhatNHBVnbm6w4UQ5w63Jc+X4n7ON2q14Yxxfetw14kcAB4f8X0iJdP+
DTwZssb5i4eA6LchMovH51n9dy0kjKfSLr5ZQrXvzEEzYadnIVtRhaZd68jtiK3WjVy4IhZpRb6p
TM5SBcVJBke5GgCr+3k/a4d0tu32UCrXCB5ZI0yzZWU6TMwM4vJ0gMoj6pFjfDxxL5sIvfQGsRyJ
upBemjzlut7OKKnOuIYVcyeuKM5n3+3sc88Yg8qvJ1Kr4M/IATtf6CzuPjclxCLwgFv1bL8JiSUO
zhCRAjDk+6jyIgH5HGEYcwKg2XioNgTbJ8WS1zMXMIihAkcBJ4xflmc+sow4ksWJaXb2Ds/CrKOO
B2+iSuLwbIO801vfAZrMTLXAeT/4aeLjvlNgsOgZU0TiBOqBpm3bvw5C041mB1W1WbOKoUR1m7en
+s/Oafnj+a7LxG0wHmGHyGHTbyOljO6MbHCyFDuk2dSmPnaK9q6PJLRbmZH7eB9d7uUttXEZbrl9
iES45Ep5N6GuOuTr7vYAEvzkhRxtxj3NCVJS0L0gwierY2Dp9K+fU6I4qoo5pDnbOh503223zFuS
HqCWoHX74vYpGtwfkx7VchFrd0Q1CfAIrNtXqTvGNssNJwHFugJrpCptvWsygZrQqbevnO0nLfjf
XU/4vaos7aGEYNiy1ieMmDcU5zE19Dotd0zq0+/XJgahmlZOWZ6SCC4VhYmPEGnp5W/n8pYInSTV
F+KfiHMyNETIFB+b5PtLAqxsg2YN1R0b9bUVWKowJEtO/VpejnBod5lr3Xh8bu/ABj9wlp9KlBuR
2qaLHYThoabxCqzzvlgXDtJUtzRY7fFBuXME7/SuzK/dnu2sRRkUrtw/CyMXRT/3VPDcWdqhd1Lf
26bppsW6OEK7f5veopF+u9LPksdwFKipkKLun23/7HZ4NLy4aL5AbQd11AUCzQVv/Y0WlQaS8CHi
kK6mT3dQOZQQTWM//kIQjusQvvibjXCFbcOWAhzMrxKeTuFpoqr6qB9DtUzNb9852gXH/Zb00NyZ
lYg0vMFQw342YqXQ8VzhfpU0xUfANwwM2jYIvfZaAO/aZo3JHKT6B+xOgm04pDbqorf0ZUczjh3z
AgYo4+WAiaPgm9YqeJ+yj+gKL7JwC7hpGIwXClyFJmQGcPVMi5nodxn8Q47SkQUodSAmQHtihi0M
zlRP9tZOsQ8siWBwcrqW25SQ6Ah8k6ynVBFgqvECCvotBMrBQcIgZtJ8Ry01xN65/dqFWTN5juNg
Y9i0KX+HhDtbAA8QalexHV+cBZmrkMH9RCL9Q6a0XloaEYiTHxAfFJtp9LjDbgYAtUvCPVATwjt+
DV5h9576Qf0P7tfyPetB5Z/P70e99b55Zw72uHaPAtK0Onkz2Ik67g2/LBxGfTPk25tTX1v/FzsI
p4Cv1w6U0YfqdYFXoZdvosCR2RZP0EoI9yeAaYOtsUgVG+/X3jnSf3JKM2Zwf37mU9P+6Y+GlwpA
a8kYgAsVwJWEX1MD25ASloqVdrCaw+tqMRQ88rHYb9h6ijQTEdeL5/tfUh7WN1sfJbJkfBLhuxZF
Mp4XBeunv7J3b/JL1eQGnKJC2tH6K0ItwwZG/Kya0J5v8SPtK/43speRTYWtXjzepz70Va40eDIn
LQDp89Kt7Pbd0yZZ47zgqjumcGkR7G8A/iBBrfVKbVqVZN6ri1aNvc10ig5dDTs1HvsUwe5V/YgL
mLw/IQzVsAczvrFBh8YX6DBh5dEHx5Il89eyJdKXaJoCe13wwzR9rYvF0lvrVgXnumwonMnlh17z
Acd9suUKsCXg6EdTJ3lPLCS6RPISo3T6Ld6SY7qvXieIEyJXH9DaMcYJgtLfTj/QHzmBHFhsxGQr
+sL2gTkvIAEFf/IEA5cgVUbAE57WQoZA/ofg5S0u17sIHHlGn3PObmlKDM8k63gtsy8Tu1QB2g4o
33oTOiKDUZ3ssm5Yup33/V3saKOygHM0+ja47NBxERkFiCKJ6H8MZsShxRq7zpO6lJzuLQCrRph5
2F8Qat6rDYcpyrG7iVLTQL87Xq/NwE4Ndmn+4rzqc0PExNn5ycydtRPYPjHyHyTjqF01M4gY6yhZ
xX+GWJq6Z4Ov96Ir4Lt/rxgkXvwDNpzUDfbgCStgY3oGoIFEaSpnIDAOFzGRa/hrFB7+rmDLR2uo
X93g7rDBcLL1FwRI3HpmTL8idRxEmtx2PaKNPe+6SC4RTxucnfJ0JHjiOCIipeg2PjFu/+ZhC5N7
/hSBVOMGzBYvQrmphH3PIhndagKRsBikMCtkEfiS5Tx37holkBon6cTqyzPurjIspnpJ59z1VfOj
mEEvVFDNxLfLFSnBUEls6DmidLib+jfcodWLxThMeZtvOWGknB/6xXgH+EFtqKdVCPPwdwUjLJ4D
g12Al3O9iKHRJDd9MSI962YpfYnjwu9R+spSHPfhoo74/rTAAtPraKbMQV0YW1mE0P2J3PIl6bDa
j1p664HT/0piaOL+KPOYRCHJTnVj4tFU66gtki6rp3lZMiCv+2QY7QEbVHX5bXtFGn+RquNqRXnu
9DGE5zd2xa2btTTj15miamIibeAdmwA/H4IvmL0Mw2jj2qsbpDF8xdVeYLFIEl6mRRQ+cTEVFXCP
3mrv9CxCy4KV+ykXKQisJu5QbZujLDHgqUD4HsKTfJVePHb7VZEJTphozWbHZg6Vfn2fAAb0onKW
4vkUf+OiOX2M8JXNM1rAWDlalmnX4D5tqaIN1LGHYAQBFj0m+5naJAbqMiKiL+ibsdXMlrXukou5
2ljhbgubDEIU4/Y8ZbWGMq2htwKu93YbdDFgEzD/5HOVEv7EnzysLGf2V5UjMInbNi6Zd75J0rhy
KztYRhyseGRcBU0AAkpHp8ii6TroAv3uz1sicMBW5h38f6RhzhG/XH36+/AVwxGaEGo35LCQZ7aU
wKF6TZkl2H9FGPtQeCJBI2jf+Nw9iIEOEylkOQB3cml5v2nUsw0XwjvRjE/Q8mgSFtTSpZAdYgtH
U6adcOgqTwdUCgC3gz4DoGsNA6A/1iAjLPGvoBlp39Nv725mbklgAbMebvBNyMUCYdlQ2ruH12hN
lfFHWqTqSCfHTiuhqeHUvV0zEMixYkELZvUOHJTxMe17urssXyNq+h1EyPPdQv9aC7plR68UvIRw
fDwJPI3PzKshq7+VLIhRHfFf7qqlFmAawTnarLYqWd8aDl8qN1GpPba8N4+ZONV2pUWUlAS7WdNl
JEdvWzqwW9eXnv3NU20el27fUtUDEYzm4RQ1phz4wp590hTNoPA4+Z9UnuHVmk+gbtmmSxQMQSYj
r6BKLfkWTfXoD90WcmENccG90bs92phD+kqt9ebtrRtrQdnQN+t0tTmzb1Hgg+AfX8QFAnEqZL8l
QdKLehNhqa1fy34o3iJbBkoqZu12/tqFSKOce5FK8hzt2D+W/t82mLFfHFcUftcu20lI6sdQqfMY
GJdPOs5sakH4byMTsDdU+N/qpRuTHHK/FQU/UtMKBXw+9yc5PnH+6F7gg1vuH/6sxj3uOYquTv8l
z0KTdnWnK4Gg0C8bMhJpiL/Zan7f73CEsRF9xJWPP7be5BOjRBdgmY8BmynbQcg1J8aMqVOz1k9M
JT3rkzdyeeI9GTpD2lIfAuKJoRgnsq+iH67z1yNR5avxFZyOIBm1eOCAkoI4k1jP7z42G74k3/a6
xKPUkZiuMEki3OLNyRXJAtdi9dxT5OcdRaEIyvu1W9yhrQK6c3Bry1jxPMh0Q/LpVrRFiIVM/N3c
rKsJSC/Xu55/PePPWuGIrKYqoH7VV84dIJuq+yf5p6qkTcSQSwfKk//eJT+v5NIV1SbIUjiQLD88
KUkDk9RRh0b6nEy0sJ32xqvkLCv1+jmpbtBlWp3+i5PecjsRuMsXMqC0skZ3oZYVwUS5J7dsjdy/
jn0boaeNHAWD+PqPZTclqZr+URVEH3dquBi119mIXI5+xiDVyA9OZtJGyfhuY3+wIq6OoUEAgvjd
BI2Ce3bwu+6xZwAHIkr69E4lZfs2A2X27kMV76Vwixvq4AG7EjZWZFETru3ilJvNBCF+uj/X3v2D
P0umC0oMuj4dX9JsBuZNUhfqo50N6r++JM8IWsEiGGrHTMRYlBV2e/SBQBO29mZRzVn4z/ISHFJB
2naozVGXfX/1ztLLib6XuEGpRqQ9hadvh616Rv9fRcU31bYHxqr5s3Gl42VmemrvxtJuc9Nc4blG
1tfSGVxIChlmXeiYUCBC1eVEqJ4JymBa1vkf8sQnja1d7TdShWuU7G7IEYVWmIhLd/Yxnq+JSd3t
Jdiawy8g+bbKKSSbca69qfu2jT/OvB4p+FSnKqyF43hLx3NHwznPuysaB8oIVDuG2zRiIYgx+u+e
tjH/2NttFxkl0tDzh8BSG9/Ob8pcC8M1l63q8Z5P/pu6f2QH2IHf116M2uZ1Q0+xHFV6n1stHOaI
Y+Gq71Mdnu+Y61Xqbtef5bE5NqW0/DM4QeHFs1naYQEV91yetPMQBXYML9idStNostPUQEO2xA1s
QSbi2o3VGWI/QpPgIhrcNW0YGoQP62LBWdHGoyYPqT8BKBsTCdOP3RCpd+RshAsMERZWkkb/IZxe
9B04tQ+qwZZcR3XkdtqMmYqwBQJQ+Hbfwn2FLczEGpyEEnnapjRzU6BXG4cJBO2lBXGYjcnhNNFa
xU0q/RIGp12wATe9Txs7fSsDSy+8L/MICVmNcDnpBUotDI1eWo+d1cRY58un6zfBLBHtf9jy3V9c
XlpCv+EYzYbf72JNr62KE7U7bo2pTFN4WNN/PV9tCxWa7GvjetHqn6Y3PZf6XOOZy8PkT0/6Gf4Y
3w5o15obVy6dBy0jy2pamyh/VrPU6yke0yHhOvDPfj4AJGbTWyKhPombS86AiOZcEkzdHYf/F9nn
LNy7cd6Uu6/2j4d6HznOXAQ+4QRqLDY+6F4ccJF2yTEJzgfwtrgd6S76n8Ngrs3Jd3qaivytWwuh
BUheU5hlnzQypYbIQ/l13La8GPPnoa+mOf3By+E5lo4/dhokEueh/j7d5NoVJA+w97VHZQ0KZUpr
jYM0pdl/masfkALOII+y4AovYhtH5EolcbpgyaR/zN1dKArAuBBMBaD4UaSaiXH6y6ws5IvunHEy
c+zUjCVTl/XKQFES65WdYAK/Spd9Ujw3LMfk2W1SALzboXxQHyO9j5JeGDp6C2AmvWTUGeKt3mrH
WBSLs3YLDRcC9pCxg/Hydf35HszH8ocbEoV3puluskPkUfYjc8zxrV8AT4oLzt/yKt1EyHzqEW30
8vy50Xa7oJgyNSVbfMLZa8cCxP1oNwbQ5JlU0DUUTdDy3XYdduXu8HCTXg6CMr69PMAkrh7+3Tbe
Ij6EfHVaDVtLEAXMVsV6KyQaQecTGRKiBZsmj6XBfhkK1Chg4In145stqyYMpwJ1XzCTEiQUpiQI
9gtNpfeR3iLBNmMNuE+0tEb7QgitpO4SsaX/b0PH1T0+kfKV6rHZ6jRgNvWJTmk9BD9HiCE64oDm
6mAf0jz14oR3cLNZVMdWgPQwjas9a4+UVC0YCr/A87OD+HoxoUxQUlLJLxSlcUGIGu9+9vbnqyXC
nZ0mjwCoT6PoFcZlfLKUGV6Oh+Rx3F6xoR+6IIt3TZ/F28zC8+ai7tsYlaiFmnOPOisfbTDbeznr
kq5twBuAysHPwgz08oE3p25JH6+ObtNhZz8gRYqWL2zI0a4n/vCQyQ8BDHOHx34JwgtxBNl+ULQu
R8BuIJV9RcIdw/k8t/+9lnD6xvn/P6FNFs4cx3z713dYUIX7+VOhXwQmDijHVuzEjQH6WYlrWuJd
7Q6j5LL7ytdbq2mcm5r3uSS8KJFLJbC2EWmwxdSiAWszSUQ9sOjq4TK9yTdzbDvVQBfgENOEwQYZ
uy/HjosNGFc6wPm+chy7jsWpEEit2g7OsGzT570xUUwVcQA7D7uJ4YRdHIq0aSf6tsGFSEaYz31B
DV+eoJlxcVEhERBpOa5Gn09QkEUPioubgM2f+iUclx/wIxxLBogCxYBZdEwtyVk62V3oknVMJpY6
LegN9yDclH6ymjc+5cHBCbmdc4grlFTGs5g4Abi11iLSoK2NudsGc04LvFK9CTZTY2liIBWGLIss
WAanQJc7jX12sBicLqj96qXkpi7ZUFvUUdbSkxtU9nwdoEgTY9NeCgpPXzfQFoE1RB4+P0jhKGkc
J28dV+AqHloHfqZ24U1ndtU6BxO9XE6ySbykAmLkBifCaxDw6vxXhh17x4lbuwCPRtb8CrEHpTdY
0So+hWfVXd/IP6eKLXHFx3l+9rmb09JdIwuRO62r5v74Y/g11HGsEihi13uDmayjq6e6RBtyu2g2
gQqpKAglE3GmQfHWbzDelEyREEcI0GSmBiWzCgBOR39nzXt1qhl42QuhIJm/WQ4xpgNfZIO87syo
X0nez7pH5KJwBJSSo8LvfAlLtIVmKHKLLFIJuzKRyG5JeORdBKsDr+UnYliaDTb9CmHS4aTMUiTQ
Chdi/WulHPFJXDbhw1LudyTlE88EI02l7YBw91Kmms6PFDpEsAeZuEKG7agINo4CBlo6Fk8Zjivr
c5cktqfKJuXe08Ep8LF8DfP2e3xxDR23AvMm9eRbZe8mUfeX9GZ3MujXfXN+caH7MGMOFt0xXsna
4DdAy1QhkEaHqj8bPmH1qXBNz9hB4Ae/CMISHdO8i9G1xdhQvadxXa0FIX9VSpkK9ys9B8OvAyN0
r4jMJmfXbTMIKOK8z5ANgRhIdFVgtQZL13I6ke+2CC+O3tKz/SzoIScEiYHafl3pP6LdQy7GRBi/
0cinuvzb0KqAE1bY4yU5doiVcHscBMYprDXZxnBbt/NOZDt50yWTqzlLJmZHgEetfHS1RLJVvW0L
TaismPV0CUli0d3f08VEvx6J0ve2GyW9itis8GQjoQujuZC08odBrhXOCYVFzrSqmnllEzlwLc3T
OkBcwD1YQtQG2VMFI7OOju6NnxLsKvmaqOQi/1sfxv2VXNYRJkv55FxtIfVCwkBfuuqZoxkKi2bL
cu5rDOtv9s0xf6xCxbA0owBZh4uPVm4uTVtJCl4/aHFfdRXqv8TZiq+7Wt2GS/km3se7XH5j4sSL
3eJpO8J23aFlAD9/DJK58AHWoAsZxT31aX1zP2hbL5+8NUWxQuvn6iZiM/skIIeGX3nolsyfqM5S
dQ4PXvYbOIBmh5AakaKlO65d53NTGlypQOkUXndvsUXhQIkO61Qr45vm19wF+lUtKBuemQVlWOkr
Lcu7nvVoc0UmjwOVxNAZWJ7+6+etpFWAknXF+BgVLV8D811jXelaOpMYmjyvlJ5oxDQn7mVffiLM
iEmPxYMGQLqvoiImfmZrEeUnunyyXVmtb/oEyuLbeZ1FcqrHF1KglBG6SGZh54UvZ3CAVwjB0BJ/
TqP0WysC/2UfLE8+tBKtnpDTRU2tNC+wZBn8IVt/RBUE008apIQBqfjByrYZKwoymxjUtof2E62d
OqgMhxL5TL6P/Bl26xsuMITEm73XIUgOpo3LIjkt75OJ7AjIehb8lgcsz/XEK47O9hcNaDbN/gx+
PzbXtQCNhOPApP9OvK4Pe4AZbbNaIK73RzLAaFJs3RoSbwehdwT1kGuSfp4lnr4yxsS9y/mfyHHR
vVUgMjHpiE67RCIsKEGWHW3s9FsGOa6ovMMEQHc41m2/azkt1Jpx5XxgAALcsj7hlzLemfAgRDAv
r1tytr5JPYLpNX8ISpzjFJJN6Hm1/kS0b0pjOiqOnkfGp/x7iSxQxiuANfifKPbKJD1zVNWYpXn7
YPD3OuZXGktLJDrr2bCUxiARuOj6RwVZN9NKFmDoucYzYZV8X16GSli3zjtzKpzFvOcdmnWMkyz4
yJZRLS3S/WvxeM81FZZ4xFrb/LHUjV0gzGJMgO4tT1/sQOi88f90L+7vFY7oa35OJmVkNPU5pnh8
Migk4JDkgaE6OMKfaPta7K426Dgg1DThg9RWu3emg7ptASLLSinEdiF1ami7BU2YMtK8Px9Cjw0O
L8kErQzH6k+HgaSv1X4HJRgTsn04GeV+rzKtMYIqHmA81WgHBxEZb5n6J6DRp8TJEvssoHf9N34m
DnFe71LC0aLra6lyJb6iCKdp9pDuHGStOFiTqD74wbuYPEpGnXOEufej3j+o3SVqAGKSQTl89LDp
qICPYeVx8BBOzUVehb6yVkovttlVI2wd5iTuGcAJOLLabvpEBwlfVgsZQQKiwn4r7wdN6Q15YiWx
WyjAsH2djqIPpI+b0xo/iNOJ4Ftu/zGlGwfuQJzCgWX3fK8B181q8DPwqOlkIKGVT1D0xqJvXZpb
vgpSnuCBPR/1t/+w9wm22wyMm76p8pV2i3cRfcOsWrpKkmxl74qKjBCONBC2pTQbLOjv53tYHtxD
YR7SdxXt+tSl0sBvOXmFtAzMSFmrqMJ+jlUF3kA0W6c8HqwwXIrS6Az/4shwD1IC+QLBhq0b452o
JiOfUMqXVSPpkQ0dF66nFK1Qr09p6pdk5YYp0XICFBi/K3D+GgVVqzAkwq7B2hG9L0qv8AY7e/hJ
zmynFEcOO8YMj4ELr6JSOIuHaAD5math/HLm1mrv0giseHGSCoGkkPoy4m0Fwa75OXXUoFnPJNAS
M9+hIew0eoSDSMJHJ7fI3WGFZldQ+35VvaKGhMyf3Jfo+N8bizowSeBi0AlrrNkzOFMt37NW8UnN
vMTt81EkhEEzgiKYw7bBKtFG7eioLGVVBs6ldpRG8qF8DSoPx+KEEsu2LcYzrsJ2N5g7hxQjJzYN
CAMfN7+AZwmwFXMq9o9Dd6PI081QOxjlHo2I+BXKeld5LqbeYlY3zPw61+/vejzgoa7REvDw7oEC
o41xqhw54y9N5hXNtO9rcltfUAUWOJlWAPzP66LepSfrdrngvYQCRJS8tP7wI5NskWBBTfbDclCU
aPshL/3sD1mVih48Qomzz9cWDXWRrNbXkXJ/WuajJAikat8etKJ82IJ3fml1TQERE2mfs5fZzaTg
jCKwRRC18MzfGSICtC2FYOo5X4w8vUfdu0f+Xw7iDA+/zqrVEq2xXJH2HiMryLpCjw/eBRhxp0uF
FjIn/LjC1lMDB89CBI+rohMWjkhD+mUMV2EuFvulU3hxe1XGR1P+ltZDRPRjLUekVkrrOF5hId7d
Au/g2dulVNydDeluOAFvFU5lUH02jNMMAQTJWMOS5VClonwyjB6R/1cngsKlOokKqifr5XJKJ++f
tHQUJ8LZU5KlkDMy/AP7ZGXUeMWKLnXW3MsvLoX0x7mVEl+9N9UFSEs41Z7Ia0ZDvj0vjGFx/H05
KIE2FE2Pdijm10Fb0oAHnzSg9x8QNFEjm+Lgt9/BuVlZ8OsdznFxXK8A5KtAlnH3vAf//2nzO3Om
+u7G6gGcqXwAlZyBl/DAUNzvXjCUFn1HklA8sw3Y2YBSMjCArzYqQ0i2fMmruVf1pYIz0XtQI15P
Wb6YX86K9ZZLhvHX1NdlQRK7WqtaZPHZOQHAfYoLjk+nmxNilKySFciA6NBiBNkmOOIJabW6gOYu
6tDTZ18RqY9UU0s5GlmbDkiMXvSvA+7ePreOjZUJAojO1tDSSO+cNUVlBJteWyxkeBVoJbytEia6
TVRe0mjeUbIMGlHJ39DHMQQQYcJQH7ogaakjwy0F+xU5oRg84s7Hti9cEdC6CPfwoobAjFwXeILI
WZ8IJT+hjekWby4gXYpSwjZitKKGLY74EHJKq9AeAC4H9jBBwuseAtTf8drBZvFra0DOef/7GFGh
VxLaUOyiOpS5pXhAfg4AWC4iKLDxdnKarYjB3+q9a/7m876v3t4O8Wxly/aMUC7qlw1ULayjJ8u0
AnZzGek7qzlFoca8avFGGPFZX0559vNfFkdFwMbciCP3vDJOKaT2qhBPgMI4TYZL/DeXhsx87S4O
Z1LLcGUjDfoW2+bcSRRGNzeFa4gD8v02ZB2pUQ9/D3c+dM3ixanN/2JuqFlQ914/aDXlzsCsqSyo
D2MiDStl/UT4AxEukkOLUmxpu7eOvFWVKEEPB7o0GWGr+i8IBSW20rNg20HomHQ7mLwcJ7NP3MJ3
rI/DOmrMkA4sNsiPik8PBnZLMibAkKYW9o72Z1pWOss3ILjWHDVTfs9irL+uUbqleMcP7vFPynv6
1mm7B8LxcpSnKLderUDg6XUwoS35/XvbG/aQmq7W5GDHLN2dQIZz12mwP4qjna9syhQpaz/qZWYs
A4l4SGNb05c51SeMDhXMPimFG416ESKypo3bgAxxjx6mqAwVIUSRdeR+DmuwRHd1K2DPjm4dV86p
ZczfYIM1EcLzIKu/a2wytEMetQ317QVHwuc18fsjwS6WMsdCjDvHsMs93F92bVoVxOIBCufdTPJT
ZNkOGlkHLA3oObM5OX+9ySHfs4ByrjXj88rh/Z0GZrOR4WzgSDclhuHoyxSSY/QH+/XtQwmgR5uu
n0RBVd6+V/dKItTaCM4CrHRmaHzDMRb6szgWNxOTXo9AvoWZyl1BCrN8Nrpg39k2nWt0rEuo37iz
AYCs1+2J7nWQdc7ERIwDVzOV8f2VuAxVUe7SX1wj4GPOUIXs62BZR/n6nhxKprIfzkaues084l3b
Od77FSLn2HOPgrkAxKVFH8nW+N9ROC1b4Svn9oKcUj83f5McWQkjvfDvcd5j//GCH5mB6NepxxBK
+bCD/uc3f/sv1qEgQ4WwCDtEk6Xflc9+lksQfpEZVAei/XOv/RDs3B6EAZvcIRqdZJrv/tHaO7ho
jpYHTwNX5/EUCPLNB35/O+evzy0LDkfclfQaIMyWrUxf4mFidiJApOgim7G2UEsR1EQWeYNQSgwi
/6icrx4qmf3PPLgsp7wheQlsoV6fM0KQ9/Qb7LEt0LqXzrSkqHJSMFGUEcEDo+7CVPcyz4U7pSve
nQ5+ZoHNmV/r/j+QJ+WA54zjNebvLqNHhtzLNV23Zys4Wm+UP9LMMejzZBx8VNtuHpQU2SQ3BD6w
kbmQz93Z80kzxMO6fyoj4ggWBq6S0NaCWIq+FWtQIMCElXojIDbQ/Zs62aMrV1OZmU/Csi90dOTi
jVAaaI1AU+5O2deK9+zxDWZlYmqfs3ewbSX77QMLa98rS1JRF3Jz9TN1Z4+kHk3fCl9FqNh2BOnc
2FuEfby3eFhoqEqtcpCeYBwFdUb+hhzKNCYWs2NxUbRvLZTPwa5HKM5/yPllfVq6NdJwSLwzpddb
26WohprLOXhhf9sojCLh/e6u80mpVHWstIQnUH9wC+bPiu+i/sD8rLy3bC227iUxygJuRcYUHbPh
pG2hoogBDA2XPjGx8b6i82mZz6S5Hsx7wbUf/uT88/IaEtnYhxV57awJmu2iFm14YvUoPZfzHE7/
4Y0KF5drTFAw4/3XgTOkrdKMxAPXrERn6w5kyuq/v+/NZiZWj9/9QpQyNPc+vpZaayOCvhb7SSEh
v0tqLi3ik3VYxqAA4tcAvBoumLbb5zs2VGdZXJLMeaP/+NRRwg/7PzfQMEmIDg1NilcwanHmEsH4
6wdkCiNqGMtWIs0aJTHZzuyuZOBqPYv4k+a4HTc9ZAMYBGVHDoL/wSV803IOVnNJPJ1oMAVfQcnG
psMk0kXm0KINzOCGU2EQoAL+WE6ukburUHngVgJmyLgL2cyZ9RaVgDcW1xUxMLm+mAXZYoc9+VlN
n7zdXbLR+6isLQTUN3u7pkez1iYradl+1nNw6Dil21LAyjv05hzafAClulyVEuuxHY4M2ttlbP4m
cWtFQNXn4Pnhz9ZB+ARoeuw7aQZXmh3tjO7tCsSiD+iQTwsvFoTVNrotla+pjVTZ/EoBZn7p9Ize
O2NO8cGCjyDegGyQvAO31Ih68DCk9Kl8IrqoRtquU5czNPGDbc4YmhCCifO2ZQ56YWksIvzTksnq
kEg1PG+YxbZ1qzDvaL6kbqcS55XXyyF9sjT5sXpmEFxFv/dWjzNm7eV3dp/8iiudQCjzMZLzofhD
KQv3AGzffX7B2jFc3Ak7gJgruxYQLUOnFSy9KlgF5YRfRctdMkXtU0F1aexm3AB25Dtzi1NmhWZW
lISAGPk+nzMpe+4C3uwu3chQdgDlnq5CxYdhuZeMnLX8uDDP0W0d/94/XWEKS13QUsQtNVXvbrjt
KqPsdJaX7Un3sTNJD+RK2IsF2WxGhXnGlEza1fnUJRlo2VKy/LR6zYOFH5t7hiwURP2Sj8gYBcxh
SfdqTQM/luB19wKyptCBGlHtAJ8VzVi8Tr1wkgzUwgDFlXSIPKF/ssDdCR8MXdysBru1yT3Ycqgz
26E5dCo6YjZ0X9v1Z7TeBYF14JEV2PAuFzwkB4XYZcna883cWjrfL1p4gLFmWHpk/57rt57MF33R
aCLn/pZoPf2EQd0Ob3Wa5i1nZrc16MqOvY7PeCTSm2woBrR7uYppwwfA7Zp37Wd4j87RD0ALiDta
bwbI7eA/ybWdbWOsuyXVa1/JEjSagHJkez4Y2mzuAp2rbc5VVc4GImvu6+nozTpCbYJcvqxshYdN
lFm3hRIEMTiqJB6nuCUqQPmXsECqzEahnEdoXTfbjP5A/WSZXt8bE4Y5wiHMLMOahRR51DFULWrT
2S6gfKVoHbOYJiyKkcmpQFYW/sHqd5vnyV6HumD4aXLZuAXgpLtpNQhMPieHRBme6qvpW0UNXeu7
aH58Hrr/DI13XzG4nTxNePQA9VgBaDKuSiVjO4v6mTAxwqi8SVuzmDI7afcQeOgPAyvsXvTlvdwi
ptd5PEXqYzOus3b0e8fKBwYDUq4vsF/eTCuEaBrF6JpbHvchjjO7VikpZgZORZhnZe2AmPqX3EK0
TJ6b0VT2+ayRKzv7f2gh3ub7P14hEmX0EPPd24n3jEhelNO9Wa7ReAOD3uWDBhL5dj6ur4DvTard
/yHwrhy2HdcdGh+6XLmzd17ldEoC4gxc8D5xB50YGQf1fmiS+EUrTvCVfBbJQVHjYoNybJvUT8Ix
wfcPgTUXEPJKmc5SDaVK9MaijQjYB5C4+o9FruRx1uykBzYAwq+GCjCSHd5nJqh9iN1xJnh/IuwV
2OzbtswhySB/46+TYIAAqOv8g3yPlKXsFkTlCCe49ovd4EWd2fYAxeqjXJdlnx59H5vxuNdbmiIj
ZpDIF/b6DXPvShUr+PZAFeMzTyjP6+iOE+8lGv0DlNBN/8gPPUQdOGAEdWX0RGTFY5y/I8wZm4Vy
25iUcuWJW+zgGa26eyRx18K/3fmoEluBnbE6vpXWOd40fgcVPuAx81aX/F9yOTYkPfmBv/vAL6Df
x70GsWfNID/qTERhQjiKYrpG5ByBYvM7LOv9qhwYkUPCQODmYA6HSpIcdhruJej3ESbokwOsB3bV
IUnkmj2J61oQdt+FKTEB+/JPV2DPGaO6w/8ZaxZ0X0qRzizZ+bYHipunnH9Hbt8uslNmE64kURQw
wRTXc81Z4A3ZFJAbWiJe7eRE9VCbJc0s0iK0r0AI9MV9cHZmHBF11/67oVhmHXEWfITrhVqg9/Qi
XW6pyisq61iOzgRUn+rXE9fejRpVhUEOj6/k3zTn2LitlRPXt0WwhBkZIaLH0EQbnc/YjHtW73yb
3vZiRoUPTr5xXxDShTwSisFsavpv5uIaXHS9e6BhsHazdMswu2BLkP8eMaGDNxwgJGxpKB/GvLeJ
SAhM0QdHC2e9BKIpvzRti5PZ5Z0PqY/p5jlVapW57sJE9hFbIaDlb2z8OQo63UuH/pMlddOGws72
+uXDlAR2Yt3Fu0RzndJrhZvLf6ySzCaJ6F6YjHTWtRJOaiF9ZtDon9a/VL2bBUgUxZcmBLFxsAk3
0JItozfcAVd39j+RDpcXm772NEjN/jpp7aw3hJsCJvfx+P8oymhVekOAs+wKVpib60ACQ6CPbdKD
lxMlnGOJdYmkuf93a2VtlR2AqHxKs7KMP1h46i9rFgDXah41jXUboTiWZ7pEe6NUwW7PQmLKO6+V
YG0cpXmONG2eMYbLeJY9EVbrnO36alTftlT3q3iiQkKpkySpcoNKc1C03QaBO3MDq217xtlhYkOP
TcQ4UYt4MVFqW+IxrifT26wSDbE1FXxz529Zgh4TjXJehs19CoHVfgCTY7NCawUYvE0jboACIw2K
vRr6g3xDz+hGGyCp1LYm5FVs8IeupFCjmgw0KTwwHJ6fQfIMbdYSlSPfYqUgFod1/i96AEXj9f29
gPDgQH/bklJ+oa6kRxS07TiXzMjg8ROsNkcnXWFqcq7xGYO/DtUmPuYhn13VyvHCsecQ3R5fnpzo
q3miZ9F5FIOXbg5T+GDZRQvjqcDyxyVk8FSB+R9gXE+Mq5qPG4l/oTZsAicCFXaM0S9nXxVxb/ii
xgiNp85XVuTPASM5YDlT5nxLAG2ho+3nd9xiGn5MbBdIluvQJQ45VvWnuBPvj18TdJKI8GHMQV8o
9m8MrwuqADkm/4Kgi3Qs0qhZRxT45BIaw3OmAHFyPCx5vPbHTR7G865KohQvTSOlYasr1/r5/3fk
NXSs+umvedCzu5fa0SqPNHf+OO4pbE+6rbjJupog90oNL2Z+Jy7aK0/63f8o6p7PmccjG78vn8hT
YllOeqRqWe4ukv+5vyAVDywM6aXVhUZP8Pnlrtfun6E6gIEXSdGRiRRkImeQlmUEPoQIuCYRSnNs
inajj1PzMK42KWutIyl2aqyMxHEnFcbVtnCsrVd0mB0e6Hf+Mx08utyKIH19MxAW+v579R9/LGPc
nZxvWzajajtxaSH/pBXULSklg/X/hycHgWL9e3qSwWzExPJXbDYTajYGkwjaDI1TVc/OD+aEHkWK
QPP7SjCmSP5Nz1egAwGQ/vMg2PU7DPUlc+X1PDnQDTbPt4JRa1+X2BQkyuF2jSSS8UpY+OiRG2Rp
YRzWbTPqAKyW+7WLUS5Rwd2TyjfByrJ7oAzL2SXy8RK8azuHHrucjlcSOCYBPZKkht9wtzXN3aO7
vaXmAmGnjbOgycWMkHudeRi5nOc8iqI5S3JqQibjm6MrH9KYCQIGQrBnUp20K2ao2KHADYH9QJg4
ru2xbddIQcJTbdu4tqpWDygcwgM8DBdjyJo9+v9XIJGZc6WJmNCivhskYR0j4xL9QNM7HEfAKURj
N2p27+haotReljYK0XLc96ilaHl2uzs21/V/cCCPuSAktCS5hTdZIDds527o4iMm54B9nfjCbdIb
GbavM7XR+RPu/uZJCuMqyv91lqrqVk4Ykbqc03ieRgOK9rHOBq9nBrMqJj7fDjQJCMN2GKPWGs6e
kBxwKG5Uy0jwYpndyIi5+E5SwFDInjhetoq4JUHzbMo6JCcTqb9WvSoQ6OILckYP+x5PB0aPZbDy
d2aeMN+pvk3y3ughBhcAbgSQRyO4uArxw9xgru9wDcq6UMaBiW82lfwssOMt5bqG2T0oxIWnRfid
Ajw+tX7mcOF4160r7abs0OJzIrgNptjKYlUSY+r8jY4WewJqPJ5+UrSuABM4hZBVpo2l5+bRjWCC
+D0L5SJzCoDxxX8OYGuQ1ABfkDN0+CPQ81Vq4/Ir9TV6qQ5ww9CSA97QzU175L8J1LtOqu0zzqtm
ubQhNoKkbaYuXPmo9PqzrDE9FLyd01Q5CgV1nb8iok6RlZQixrdA8rBqFmAAED+tDzUFla56TyS+
MRLhj1bmjPaCL/TLy2GhfGLgh+V0TEGT7bIlidQteXl2w0r6a0X/pd/zKXEdfx87ExhokXm72+oR
FEk88h8gujrsLjFY+4YEzxbaoJ6fJd+ca+awVsdRgoZExw2P2Ihi4Ho5BGYY1RwsidJmN17fxale
8vHjNaI07MZwChN1BA6S5AYVjMKnA3fcL24fThVlVKEVa/RVGl41C5lySP4hA6J0kaNpYucfb009
NuL9ezAuu3SEXZj2EVgaaahcBRZinosUTlCPDayj/+z4jHZZvgCO5nDJLdVPLqXFYsew1B0V69Nq
LGwy9RtBab7m6DEiw7HCUK+5bJmHTRY1LemKS/BbAW0A5K1i0oWfObDJoykK4JVXJzAgQPAbsx97
NEXwKdWrWUk4tI5Z54kB3SGsl9hu4h6xxjn4Uhjte0COCYoBea6jRfCKlkdThTLwetgfaJ/BnOQ2
NNaeJhXPjGbD9XW+JsK1SZrN+jJe4QBHT8T3+mtlgv4+v+K/foLK6eVRjIw4Hog7L9e1Ak/GmMV5
cmwOpdhVU1H5QqTloNAYnqEweJdOsf51c+n39xiIHoj+TTKMTOdvDW3eeYATQFJ8xm88cLJvttgy
TWcwzsV/nXfhrwygXw4puCqxZO0s91l6LX10TFcZ450INWZiyfhSE23iS7iiuG9qa6ZklQ36m2mk
ukdNKnoofNeYEabJE6tDkSOuzphwjOcivbEP7JjchvC933/DDkF+8FsGklirO4HzoW9BAHHBt1gD
CDd5qQyqUJOVhoS+jmiv7lIX6WNa0XIB3ZJ3utb0oB0YLEUHtpbv3JQz303ElxpUABuSW6fS6fd8
e4XcXLXHJZUbhSgfv0UQEnwPkg6o92S0vq4eaynhm+sm0jyR+vmduA1huhzAfc/fdpDYjMkMhpux
7ywTkeBZ3Xv3IHqZ4DW0z6xJ2bbUpskYDQX+Bi292DaVlI+6UNlxMw+DXxhhcYpjl20y1UB50O7S
aH9A+q6YASz4gdRi8Mkh0QbmEtUR7pi3QZki9fmy5Xo0E8sGupFz7anyfFVjVxX1vEq5cj5lwp3v
569eijUA6GPzYJGcPiSaSEDwev1/QNYQEze72DXu+CzQH3vDx+QmBmLBbNlviXSw1tydxXFVyjLq
fTaTxG5goIgxvarHoDddry2OyHhguWDBIowBwHsoboEDo7l7RDG23Z2RbeIsHwpFxsWV5Cj6OFQ4
0+zTTQ3BSwhY5oCognbnj2NOIas45ziknqSUteXPnq+d7JxZ/w5r1cIs3CjwSRJ+GkV9mQVrg+jA
YkRDLvUB1jNZHgYLm4yXKYQuN++z5bWLc1x/7EUubRgkMkIy8Re8m0r6r2KyqNvcL7x6PYD/MEfq
bYUUVHqcuNtnQMlqUJVwjYJUrZTOdf3hdf0LHkRb/uFVsobilc8XwwAUi/QrIrl3CszbpGcSHfit
ZoYHy7z973W75w7iIU+oyaaSc6taz5M7sZH6KXKf4xLmY7vbTa7+l0ic+eIlpMt1sokmZIU35yKA
nX0NU0ZNYDVsh+u4MvMblupMCo6nYynvumi2IoSsqv0tMfncSMIReKyO0vdTFVZEpFiXtDtQUPVO
rrPAQMuJkLIFsA/+hP9FwzornWZo//DRDWkn1nmy5jA8DO4AX45QQ87qYm3wR7haEYueYUJ/F92V
ST+iopVyt65G9XYLsPt8wY+AK/w+vO+IMi/gtNeOaBoS1WJ46196pVk/SveTyloZRBuAQj7ZcQuN
xTf9I58H5fWq0hd3GSbU5C0cPY5DBRdINTa59El4C9ngqaLPsyPVsLVSSeWDKUAI4cgUrlE4bGom
GOi/6GV0I8KtqgNezG17xfzO+Dt+DsfFQs1H9IySGbc7O/o6JCf4nGQt7KMEZxxcRaNBsZGoXECt
AXYiLjYbNVAJcK3yTlWNPwPbio7SgwiDl2v2ruQf4mB4ZKu1aSAhfnd8PCe9VKVEMzKg4naSypPy
iqW/1l8IboeO6RH2e9MSxqzCQDFvuaD5h7e0S/ZWPxE0L/+GzKBBQ80mcgXjue5qUE7tDKCG+lCm
6A9y6+NFF6tIvy0j+0Exmop1AXmXH0QEGTVqzuZKxUTYq6B50PwEY28QzEpbBd4qIhiyyGrbwtD+
9G0dElp41mHo+gffvjl8+GhjPlbAc9zjFXCHVcRfAgI1TTmZzmu4fXC5KfcWWsu58kJqceQPRkeO
J62QRpACy2LLF6Lw1CCGLTTlhoFc1YLQ7/S9ZgRUZ26bE4srhW86AFhH8dEdYddjMZlDZTjzviON
rO0X/G+Kcjw3H0ihiWQ3Z/p0KUEpaJFBIQWJm97+a6KpeFb86BNCzm0jjvn1BdzSLEoQXExvvNbZ
nsuHDmGhzbCzZB9GyUG5bstWePB9D0iATVFgPtcu9teuElZXgWUTsYtYEhKCOj5B3DHmumakK3Fu
GVyTJjnowe8giNQvY0peVXoq/KW6FI1oS3x8iBig8Knwx+3o9cJzdMNa9PhepG4bG0SvthPzLdE7
r3pirNlpGcB/8jSWY2VTUlgCRMDeBqxvIGDapvk90nt1widmvmmxg3NYSNyeoO6txnVuSfKo3Js/
7sHIUkkPWmfrmnWKja5K4Vth5nBzwpEaIkRoCH76NCtJf7RoLDm8LBwpnl6C27W+knVkH4x1w3iS
9qxY4qN3ud/yos+rXOTjWuW3dX7mag/NMQ6PDpz1buN3P1Yi/UCjNwJ9gIM0xxkVJB3n8FOqlJfb
Dv6fFFYFaOkYP+QpZM1uLPClvSfnxJg1hUhASdLWIORH0WJly6Egr36ehZsQtIj7hmXfDRVrsRqG
5QfOaqbrJdFj1/atIdR+T82W8xp2VJ9zClt6WF1cmzcrnc3drGe81VnTL1XyyHbw9cHJGZf9P778
FNON8/yE2ks4N1a6Q+wZzYTsFgEV9l2mRWaVXwqlCPA0Krr8004VlJnLzbhgDxrLwVGV6ZAGwiW6
RlqtXn7qXgpS9Rvxidgw04BXDBL+SdVhRKJYQPbWjp82OZYKlN2OjUyhSfuf07rRRL3V1cZxaTOX
ECzF3v1s2RJU/9w1ocLRwMYtrfuVXQFXro79IT6nHkdwrRRHv5o8rBnoW20WJLneojIn1A7glwjZ
TwIVK7i5RNVvugGg4oo4ZKtMzzz1900uapJhUHg/75ZQik3yce1sYNLMYqfsrRHZW8h62nvL7oY5
/j/VXxDGIH0Bhrr21Y67eN781EhzunWGGdJ2GaegHOyMngjzxJuq4IUUkL8XWXapzgWlA/hUJ4+N
yqf8UVSC177f+CnGqJ2+rHorL1Xx1TUUe0t9cwSbQ5RpZVQFli9+LQC0b1Gfoh8YMYtbUNWvlGhs
oufTGX1CDJkW/tAs4DzXshmsHwH22SU9nTQH7hPlIkMF3kEZb9ddLqq+O1b/2mX3EaoKiCfdEYUW
6i+3JXVu3NUU5WjMGakFHcjBexIxWkYB+ynd8WfH94ZmaBVxOmxCrkuoJxh4fQhRnjgLpTWLGRtI
OKd4VhgaJQZaEWO8EiTfXMtjyM9whDdRTRolwpM0T9U8n6NOl1/L6KMOgEOKEAsecHPT1T8O2Qz8
VQrp8bKuo+hTMD8c/Z9s12+TVsQrXJXCbqpYOdMJJz58/jCS31YwqrRNpAf+viDz+jfqYqynb2QN
OwTTFkV682KGWUFWdaGKHM/I2214h3gaZj7M9oejfxgGsICqZw/MzH75DtToYVjo57Ls9chk/dMG
M6dsEqlonaFkgXJAzb+wTiiURBV/QKcNSrhCFOYtdAMMRM0nr9fiuuMOLvVyBxlaak1VXEf5a99H
fU7/EDud+X40Y6aiM4xh3h/vp/LOcEb3TiK/DMReOnZ6NkYvEpiYjgBbZqLc5Cz61VhbSjqP3C8F
LJSKTbtY+AXjb248rN0AfoElCtFi+TTOuBfsu+e+Cx79gW37BekBRPdlP5uGAP7tUFYJq3qVkcCP
L6IwGtRCXmkT0guvWX+SdNgJ9trWYuiEAUr4TvAMiA/X6NRmJd41NUBBckkccBbX3ks/WVDghEB8
qqaeVG7MwCrf4PS7lczC4HP98NDO8wn8Zgp7vBONMwNOQRrKvca2S21g0K2vqNqH+Z00ZpGeR5Wp
8wtvN8uMk+d1+4vMMt7Piqr9KXd2hHw6Licsm/FFo8AdtD8T4TgUy0AlW6BwdTWTlLQ2zK5eyBv6
lfi8NUCWdjdVkd7ZgMGrd2aLESyFi2Dw3C116EDLBfAgWAHcjikV2m7OIUC2od6Xtoeht1YV2ZTt
AQpgoYvLqaptN383lNXafJlKrg4bLHaJ0ZV+mVxO05rYXvGp07uk0d/2r645O4F5kZDOLdwFryWg
F6Pp5H0DGN0sB4kZig0JYU8yKWuF4Cg8pGYixwy2Jw/si0GeQZKsgD64hoR2rZjaHL2xzZN3HSmR
cI+gfmWAcIrWehu2GYa2IAOWj4zz9f+LKxO/0yrPqJ2O7HTbW1NSnQotSl6xu2OsMWBbunUQJgn8
HDAOnQiJK+mffoNGimJfbt+u1dTE/rKOZ9mVlIuWM/jWHpGPh+MdnPij8YU14a9PbaJbSOTGScTz
1lsJraGotpy5uelHpjFFSuTP/+MZADrzcBsmNbdupcBj9mXX0iSBp9M9AwY9r7H9eJ4JBc7S4RuY
8lc/R6ecElFWijMgk+yf9wn21j+9bhdg6T/coj+LTjTda4jBmBqTB+5IDeiFtGeifCDelv3BPDx0
nW1AZwDbY3a84cOv+Lksl5QDz6D9nfidvNwGOQxvxIZt3iyenD6magwaY7uwKhY+IFWS/3sHmxE4
xGHFt8LX45YA1x6aQzFVUmGRSW9ycNBKEx9viGGQItJwhE0yQhmt+aj0lhO3Bn3ABLNvTqhW9+gZ
MrpuhqBkOdnfO5Xz8Bs+AZImo/ihybRNy8JlJyb5DaYHteKILy8tzznxRsAuZHk0CLr1P23Y35Hh
JXMymOKom/0fzXAQuVG+aQaHKA0ZZOZ5U0WlWtHd4hkLtvgGBJrpzyNK5H4msj5cgfpNRsWSib/S
YGL/LB/PnKZXR+RiRlUH9j7qg/TJ15qXV916UKPB03qTp3yH5mtJGqRUGJXszAJsTgGi244VMP6D
7zE6tqOwJef2wpA1QgpNLZEFkkE8AfaP2DN63HDPDRQjm30q9Vqd4Pp199p6oO61Z+122BB0tybb
3ulx++JQxGTVxHfRNZ+jYiIZArS38HJtcLclh0QY4PMS3P772XjZnPNacBxLh5hW30ty6npZKLse
JA9CgVs3BFIQ8MM92mWYneuiOPfp4j78e/438MlckO7F+/HTZk97Fnc8AazNQliddMPFCkoAgLlm
P9siqYsdUT9BdKATX5XXmikul1xrgDdAoFxlkRR0vDOSBqT1zxSSVo+4xQqCQOKpzm5HH+WRlAaJ
3ldsQroaZ/y8U8aRHU18caCxqGXR/+f8X648J9F4QB51As13lOdxYyWIk/Jcp4BeGiwAEqGem4jJ
lx5ZViLQCBMLNvObcKyhC+lI5ZH9FacTuTuOsW4z1oE360yz18sA2ux2KPSeW++9Eo9SObr/kw4a
e4yUrpAkh/ymsHZ3y6pAHA2ve+SX2BaDCYxR+Kl3H/tKhQUEa3AmQ5yzFTef4OvZLgMf88BLcUwR
TXLS3ejVDDVmFl/sFFvclrV2tuLLe6f/PqxEgHU2IExjFGr5wSFxud5OA5zPQNpppMD2ucevi+By
mxEaAH9wR+AG+UunPDEXvZu0eHS3RQzaaYX3Xo8rfri5iGpWB0R+7F9WXEGbQKSGA8TxcECxGBJA
H4IoWEp803cp6CkN6ed8N52M9uk5GaRCJOUDUTfl1DfpDa5v9LiyaiLGF+UvAxzRm61CLQaGcNrY
cBNpkwNNlPPVL6FXRefXoq9P3G9tjyK4FtxPb/+bwNK+/tNNeYGScc7NuOgMr0Qn5uVy/6geDgnl
fEpIkm1dcYn17E/Hfow2SP1LB5ow6RLo+tPL+NRYYJ+uqLIvrY599xIiOpErr5z8Y0gF92TdMYnr
T1Hxm4cOsoKq9MAP0xvZKpuv/RnyUE1OXuSmi7ghQGFKG4edGqAuKCPygL02jCIiiNSx4DSRXVuw
eyNgtO3z89Yi4NihT6Xop8l03HF3yG9icssL7+kSZiu/IhgcT2mbtwgXwVxg+mpLsQYJFWkYdbC3
CkJRiBzFWDZ5JLGgMVipv3FJD3UE+Uqd0EaMlUIEhSWYThKt6aZhj5slBSaKHoAumAXh/7GPCxHP
+m4VWbC2AvxH2WJtMd6InmZhD8Fb2H0iMAe9c3vevkVAzoOiorNIqZZmcFhtjIeZAegaMHLbsp8O
9u1HNSCQVVO7CU6x7so2jCquqiA50wTzLOyXakmUn8WHlAm+HegJe2CJx5Caa4rQttnucZSKm2lP
NbNL3FwUMuq++m49chK/mLwxPmGY13kv5W+TXFDMXh4dTyjHwZzFeHgYwF/6GAIlTvrGPzeGM5bD
0SgltCOvcn1PlNSMq9BYT0cBGOm0obaonm9iJ3odMwfg/8k9mfdDfdE9iugp8oD95AWjMfm7MmXm
yNrUy7L/We2bsg9so+LitnXfBZYGjO4tYo+3BsgcBgGapd9N80IWtaZ93igOaCNyIcfNr+lhbBS3
f/4ejXvkK/SqUDeXny4M4DFF/pg+yzkB5YpqycOM7EC2YC6+IKL6RktEeIklbHtpzRDGzdXgoagT
In+u+s3ebAAuD5B9tVtdZz9xWkrkEYc39lyk8+8+TXHvb99cJAxU70P5MLE3TKEGlyjWvoAY1zhU
CFmeTM4+cv4Snm6T82u4F+4pdhNRz1Iyt2NLz0JaxRgLYGCXleM77opldz351tNN0K9yDrQl3yr+
HDVcDOq3MfK0vBeb2VKPZBeDOhJ51KX1WUR74DjFCZuJ7BMDkDMwcMd44KHQXKe1Hih7iIaBckeS
lwAgBP1vCC3ZhdZlNfKBhhGXq4UVY5LreveERw3ZX/qvjCNFI/O5wh+rdEzhBi7VRMk1autOTimI
T1SywjgC4juZ+6lbD8trHTp/V4Dqh5mBGTMmOhq2cyGTSfcqgmspQr1SGflBFGjoyBfPaWpqM8dl
kpN86tsgt6Osu20+ESzZAab4Mw4KnFByVlDIhuvUe2QzwiuqENdYkB4HqOs+pstk/Pgaduwjd3kb
XPna3xP5imne6cITto1NvwR0Q6+rgqSzzyBjNTaZywicpqM5WmzvdA+OGeJjqSXjiiFa8zp78jnH
Viwbga+fne3pP1wJ8syglnIw81hN0XYS30o/iNkdtSkIepA34hBkLyJn/YZWAFnuuj0BLHG9psNN
dkCpG4zENLhz7asknKJqTvVe0u445j+ud+X9QEyoTGfVyrpx7A4ZpiqCISeQrvobNs5OQcsvNA0C
BrBWxJb+mBUo4RHxK3EJhWNIRhkg6V1pYO4Xc7d+7JIyMyU+Y3gYHjcRVxh1OEAgdPxlM2W4hi4q
lvMwb0tem70HkhT7wa+IVisJQfd+AI/PX0Oua4wHfQmEUpp3uOmdQM97S4SKLoJKbN99oHj6Md3D
l6Jr1NPKVWC2ZoZImt7t4X2bq2LvpdxsUQKXj1FOgEO3ihnTl5n6LnBzszPb6t3Xt3nnqyYWiLsy
vpyLd3zd5NvwYTsHFUzh29VaVngkc+rlOh5jZsrQejkKuBhXmT2YUVz9AgRe9aTm8qEbAo+qK4KH
h4lhqozT6cNHaFoP2fSxGsyfsk4vdwEIIrTt4KokcKKmWrGHxUEGoC6tIb222sRbxFZYVw+RPNVR
YjEgq4K/J1iDZm9IzQW6FfptdosFJzOJT6OGgiFrUktCAqp1+eaujskmR7tQFr3gdbvXamesMuHD
b92d6wiMS+PwVGAyZfS1rFY9VRQHrMT3pKddLwRBsyWFGdM9bsJtCZiF/sLUH/bRSSfueZ0cpTET
/ylBFykz2Qc13b2OxfQ6BMxmIwxfxKZBEa6cuJHrHUvbrbZyHg1sEBvjnIBIywxzpORGUq1rZQw7
UvkGo2vHmWIQrIRLUlL/pE8tbGItNZXTLlubHR+wpCjuO6cCui+wm6qMqsmwIyj8IN9eHr5XvNo6
ZPAaxC65DQdJvijuJERCh2JnNJAdxH8LitLxwX8HcgtnXxqYQKMgeQ2Fy2XfB0259Zm188szfLpQ
t8dngMMAVEPDh2D1GMGy3GNP26ob2sysWbpVXRtefvyXYA32efnDtbyeWP8iBRvXPO1gxmHbRKuJ
JKGiXyamMQ5ZAtHBo0fsgZcNJ4dRinEr9SuDwlBwVkUdjK7xcsCNDfeEkhXHwtqBB7d8+A3U9SVq
aufg68iLHiJUEFpnBK3weuq5k7nEyflWq1Gp1YJ1zRdGbtWvnAo2N/5g9NUU/eAbTE8RgG8BsPie
RRh8TqHlNdijig2VkyHct7ECSkKgbn+kIThBUtvn4YiZ44LJsdyUc1sAwz/tCS9rQWaP56X8O+4A
lrre3t2D/574C/6BKwq6oE9eRmQHDeGr7MhkVRzYT5RraE+VqmEiE5gbovab4F4mHEDjlhaGuAyf
tS4P6AG701bW8LrwoxQJQ0oUifnsnOrlaaGJOYMdolObi4h2w35qYRcu+KOjd43fcRmNhfoxu/bI
Th1je++ZGfpUi7fDzMmOPe8KSpgjRKqVwoaEistajYidjesnB0M68Kwy0fvc5SDCzivWQALJuWOA
RQAIV+t82Fqva/zptxcmk2KEMwpnXGwwDi96g2K1745LXymKFepMGQkpiERJ4yn3e3ShjoGOy81E
f1p2Yx3L3zAxGUJjc188C2lIP2ouUs9C9FHkDFNEN0zSqCl30h48yVOEVCpoMxd4zWk5XzKcTme9
1WlBPAV/ToORbpEcNpA/tGfPJGhykb9HzSAU+lBnF+ur/r7dUE5SB1dpmwUo5b32xGk+hq9uFvqP
DLicPzrcJ/rvg1W040Bt6o9mLIlrMVUiAnMBzATAJDy2FM1Vu0b4USA/ey+n9BG0Cn949YI5Btgr
a3Qf04ueuQEcyS79EKp7Ahg112+yU+uhWMiwZIfrJOJx+xDDklgfWdugxBjblWtlcz5WROkDdYkd
U1vs0EEj7S1wf49M7GFYsXVH7QVRaRgpClyxm7MXitJphWvgJBFRbqgssMLo4UdiaDI02Idrpn0M
IOEjE0pXFHu2MujLWeNtT9mcqaOqewUYO7RTYPhRDcX5cpYFMxhhuUlht3Hvxym9AlkVafAmGpjc
Kmf6ZbAuD7UY5BN9fVHETRA6h5LyFxuI+jB0oj5JsHwNdm3kwpTJly92x1iVDlyS9CSUFmBqRj49
y7ryJu9VmMGxKhn2y+apg6ErZbxZcHintbMqpSsJTkdodUWXm9ayRVhvbAxofnIPPd+FabojR2cs
aQEUfPWquyzKgcVhVNd3la37NQPaUxyPn6W/VgFAfysBl/gOAa+oW9ckwb9YyHhI2OpSluhKBozB
TePiPDyTwUGeY7sBdeaeXM0D6TPvw/XTLAXutmNZPxTHxdWFxPrHR8S6fTi+35pyJ9l2PiOnha+L
am+utj/bIkCLahVeM9cdk8ySVCrh297LcE6Ls2rGP1W1+h28bIiRgoum42VkvZeeMBpofEfIdzj0
1P1vG4D9mtnukUJrU0oRSBB23s5hcsUa2SrdTvManj5TEF4KimgRfwkWks9lmMuv0c15y8V8EbXF
sj4OJhVyDqQRYnMZkpL/osnjY/w1XgytPsq90PeAFtU1tKn4n+4nE7axnEX533h5sHGuCfoysxTI
M5XrV11QsIpY/j6lbI3QLXiiv/vD6EepquQgryQlE3l0YpQgt6FYFDodAqrGRw5TU+GR2ficteTI
Gj//buBCdGdUH+vOUnaU1vOquULl9mosfSKZfbiJGAX7XAPwAbexyfqrpueOXK4gfRTmmdCXNvw2
Ime8e5Oo3haUawtokc5zBIpGpxoM1S9+HVemvTZNdylNLjXZfAlzb4Ab4JZxXXf3JZWZzNOLQzFz
/oUbY9gowLuJVnmIzrU4qSnRNeDv2vj4fljAbs47e8ZvT8equROzLEUQIJkeXckRboUb/4MVZFtF
23LwI4+WzG598BmGPT68UblV8lCpzDifp+vDJfmD3RhLx8c8Mc9uyr0EAwkdpTpl1JpIPfsZjz0K
+ZH60RaYr1doNRFuU9lkQ9AXJQJWYzrSazKiYjef0ovwh0ENUabJuxoMMUUnw7n4Evhk40Bw9CyG
6IYv3ZMWetJNbBMOu6S/NYTZAxdnWGZKJ/l7lutWYtnUWGEAtnt5VgNC2l3syZcLkegzZjNcWoLc
3o+Ch8bWy7/w+AQW8LSRJ8ws0Y6neZA7ZTRDOATM8EGTzZRmXDC8w5cX5hBmTO+k9TTidCfUyzLj
enymqoDjfhfKdGNRx+iKvfxJmpQUNod9WZebThKmRXoMWmpCdH1vKaiZl0CZERzOLaajWhONPnT4
JxSZ3sshoU+y/h7TDlFfKrT6Yp5/rZRL94nLKVdk6QqnvZ2C4gvvVHMcMAorOGLjE4WzCWU9nNJV
uSbVpElzFXTOorqOZemoxZrmjAtHV1sVDocbQzHUOdUrn3Yr13mj56PkutZYJTfhjqpmi3IoTxoH
WH21Gim90RlzHejhdG92LDQQ2nfJ5OUCORpVxdMUn2y3NNjCPG99XLcQhoGkXrPC42P4HxHiOofx
sPbKB1j+ymQVpAwe9aaBJwJiCttwYsbkGIxaMSxP0uecTwejAbB3ecFngPkFrGtQDdDgukcqK0WC
mIFKziDFF1O8pgcStx0LHz2zUV5jBiyvL64U4bDSnEoUZFhpZhQePFd8g4ZXmjm5Q1OG4Yjx4yA1
NTBzSQQfcKu6ZZo7aauj/Nknh7KVAKo2g/mZmYlYJ0j86cl1E4U/yP0EnM7hZnrj8RSNznWtXQ+O
oKNRB8yDYev0G2XWix9dLnyT0Q+YlKU754UNlLpjUxcuf+ciI6Qja0xLnKBDev0rreP8CLtkzu35
BIxmwtnRq3ovhsaqODr+qhMRG1dJly84JvkgUXvjLiQg/5jRvvvoLY1hC3FAURq/KrfpfmWEOV1w
vWefLIX7TXbjSCTn7nC5yRVPij2WmGXf0u8kL34XaGdGgkXcLgVqIP8hakXxAISlUC/shmSQSiZD
AECUy3/S7/uFQb6NBRTmCR+PTJkuM4kKWobNd4d0vjZlERoFPjYmKlQrC+gOIF8Y3j4A+8PkWjey
evAExa52GfMVxt98Y/XyT6mnbZ54e15PHCQZfDAFqoPboeYyCm1KJMaYxPw8N0bncgpDYEf5MKYG
fkbTGYDU8JoJvBRE2wFKq/FmnZ6AP2qB3jhZHiVjdIoqa/XoQLPzs+kmGPATpMR0cawQ+f+Knrie
ybclrO3x/WRGAY44wd+PzUPuHHbRqtXQQ3GL6atfAi2cfbb8f4gcHp5giADyGCGO+iPQIPGAin/4
cC+p6EjUIndVasg1DUC8y0PwrQ+hoWZ+jyu1JIYVzh20UCUPbFIrI1KMAj6S7dW50B2SmBPuewJr
oOIA0TqUKyZe9EZj6Zp/M7sLq4dNe5IrMLqr/j3dMQwF5Dggd1uz31Ais6DYjtTMUL1dj1eLwl53
5EuHEK8SB4lQ+C8qTT1PWJj+qgwtkAtiSijv+nbzg+PWpY66mlZZloK9DduTxv1yfj/7/85jQTLD
BGRlD3zLW3qBjbBtZmwl9ra/VEu+uqyJzK1El7iXk2/zrL9USteVMXgR6AmDNhwspHisXMV8uy1B
T0brqJWqH7IeZW/HetIY8N2cmYjONG1P5s2juBtfJBA40nRKVAmC41hD3FMKG6og/TDVUqe7eEvp
B2OjqI568arMV6wtzIdZLMaKV60DdEODiyncET1jB35Z+bugOQ5dLygPBAYQUOM9ofWBGLm6nC9R
fIQVkuNNwcMFP9CFchytuDa+0ZglqwxifzHbe4kiUo8fxiYi/EwYnFi5kUHnttDMPhTLdpmwAGnS
OY6tWcp8xGtZqdfLZ7Ty3u0PjJ3F5OiSX9/rN3zt7mMbY28lmSa+asV1ZJc9wgOrS+NwtoB45gc2
VPqVX5PvHBv/6GXZY57IshmZ4l0jTQc4kNhlZSCgGSBba3ea+wa4WjlH8Od6lTir6MYAJWTSSmyo
174nwR8uF4c1txUohUg9Q5VlL+CQDt9rE7hwE/CXJ/mrX6tyPpluajVM2mw3zBzByp+YCAnmI18y
DOzyqvmvIGSppgb7+z+z1wyWpgeyoNUD+Xh+vutTvaaYMXbBIOgtkUuT9BegIaxzkc1eZxPF08JA
ejRQ1r+BjndqwyeVOOaUjFwL8ljf+Vf8jJEIkT9sphBrxxB7LbhvO2iraDaHGCo38yS0E+Pcn2W0
CTx3ExZhBHCok197eV81h/TAjzEMnm7WDJd0E6qAT0O1e9P6E9ANc6+lbvAcdfNmFQTRj6ecSVoz
kmJt5ZJlzU+qY6ofjGgEjtzHbQyhxacKHyUJMi322AiMtMdATJiXQuJ2vEAjnOhOxvuhHKUk+F5v
8Z+BcDNAop+J72hMMtzkQCGpGSUDg5fZEr72a2sxvqzlL+4CGrWattyuObXKN8XFB+JB1r9t/rtJ
3KmcVzLXyn0wciT4P/dwGaoQT4j/g/5lOki8ecqq0RyFqHyhRJGVbPe9Kzf7WL/TaMpmTPAw+vZS
+hgUH5ayf0+QsQwVIyhapZQPigepg7fixR+Ae0NWXpuZaIuyS5QuO5M8qtIApinTX6UBUMQTkkFZ
7O0N5F5dyT3ww8QGCzmyg5j1A03FkjR05si2uaaRATEeHhAzr/JU1tYC4tYH1tGJG/nGzF+3uaJc
Wl6CI+xdfhU9mnD/Dr/FYi26wVl2J5kmP2LB+LSXmfDAodlilNEUqbr7Y7MNEzum5j7rEgIhtHFr
BvVWHGnrG82Nf/csJ7hT4ph5xK62MXoD27z/Z4BG2y2hDx7x3crCX9w19VAFmWi0XFJ5caAWd9Kb
JoPHprL4vBsATgx6w+Qk22/u1baK/ohqghAKsPPneG7b+CtzpfMraGbu8EtH/UHyPEvd+zF33j+4
2sPiKPWzinLA73g+CHqhKxJPQg+nUJQuzNnxRBr2GiKsgol54ilk9s/hWf3Oy+ZmElga+YMzJ0jm
NMU7eS/Frz6k6Cl+ntxu9LBCHBzYvkg+SRs49730mFL/Yax0FfoBhhjfZYuCamEc2Apxj6e/y4Nb
4I/sA2LFfNxzV417lVD+pU3/F96fCtvPoypZvwIGRY2QyEF6aO/QC3/hB4K3Bf3lOrP9QaXovL+Q
zYHtJiaTL7aO15LwGIoySOrWeCyQWHIj5KTwcsyxfp1Ttc486t7xHekJ8pjI5iQ1EBRz/iamyQmY
AldFbS2kBuO8uLQVfjTllhE3TwPdWLagbEvrXNO1rYWEr4OzCUD/uQw3ckZQ4bXmGm6kzRApJiLE
jLGBaD+5EGgnxKnof++kQ9qbC/Q481nxLq4j/Mvb3UgLDkAEQtfZMf+yFuEdRN121JyPX/aSag3A
P7FA0Y88PYTDhayNkwPTzxc2qKo57BM1g+qECpcfJHW01ss99tF5pv5pbBapYroQIdGUXrpa+qo7
2S2ZF6D3l9+fdFx4wYdV4VEB3gn1hIHUBWwbmY7KAycxIjkDfxjHMgYh5KLavEOy3aYnvIngRY9b
Tvk3GoZGGNRqL1+jqTyAWYfr2Q9X4xfI9apohCPQfbTKYJM4lk7Kveu1hqNIsQ28O38Ps5/M8Mn5
KbdOw8NI7iXSaGdYS8I/Xz79IpWlY+raEqJi9ods5uehJzTl5K6CCE9k4EtnNN8QWhgPg/DsS0Rn
HKA9WcdHBz4b4oyQm5UrJQY865EePXLGWuV0VBO8aaSdNmMWbkkhx1a72igbBygX7jltPvGXMQ3f
ZRYDPn6gNcYlcfDUaDW8LOGqjCmgyLn2bJqEDjidC+yi2V4Pd0pWPcYxrCE6Z9Z7N2mVC0tuLKYa
B2NA24bHsTiB5gQ82sXho01U+Eh4PeACbq7GvRUJb2hZG02AlutFDf8etxz9zPFKHwMU9vYJYZlf
i5RnQoUVX5vd/AwO+AoQit332RQmfmXgDPVpDjYCm3ZIFDihcqHB5neOi5OyJI5YiZJIt+gvymqv
LXqkmVBiSWoYHbksQCwX1zfjGrZKAtoxB0qaJIjlzu03IqC2/jh1KiiM/M37NwodqqPHHlkJTS9Y
8GUydkxUrh4O6USGt+jwQ2ZG72ixra3YL26rOeJLZqx1KuYyWrI1S9/skrSuQSsTvakBJbBMKO+D
R09WdJi2aLZImkHnBnYlfOw64a98Q6sq2hr2Cv9ATfdjjv/xmxkInsoYJgyEDLXe0+9neROBUzJc
RNaHptF6Lb0p4KZA1sQP6+K4lAU2Kmk9iOpFcu8ltV3QdeJPX6wVL3xCyKqzu9lfLEDC9geAnL/c
+Hnw+WU+sTPw8HEzBHqK0DCCJ2WqTyIgvrtTMaxyo8nAJvdbf+ReswWZnzxNUUn+ZWfQQsuZQDMb
YVsPVxbAQVyoQQmv02AWAa/SsN0N8n4xf52kLJnajiQKe8rKO1yIiFw+vW9Ahd6roqnCnmymo31j
jNG5ga0Gw4K7XINQ7pxtnLB9HVRyHH04RfL5pK8lKZ1exrRgPVO3U5TD06oNL9kgNylZ8UV0uOm+
IbTE8Wc8FtjCDT6AOTxk6zcDgfN5kW0m1xqWM3XttLKDZJaUvKkRU0OmbeCGWqVre0wxeZLF0nHc
4ldrGNdZ4GlI7UY9XfZqttVG5R982q6FZ0vBYalxHr59JowhGFVpM2UDpQjY8O6MgXzMGmIz392t
sL55/V29FArOaqQ13r8jkDOccwnyqNoPH/1G9L2dj2pGtP6xADjCwN8audRcnWi9XfRaEiZjvZGZ
4biQ6Hq64NVF9fb5u4K4wwqhlf9NGK+pGIaRJ7e0VOcwnAAmVvGj/jkw/g/amHqAzteuy6ubuLdP
x5ome4qOpx5wFU14N9qe8gFNXwkF66fd7Vs1nLeXNq0oCnx6G7Eem9RpbyblfSPVFsnbuc5UmNth
ANcZOXq6pUMpWjJp37o86/OXR8Ihy4XXqraer6STyLxzCt3+bf1br3JI+QfeSl7sZi2oh+t2qEo2
3yBAPmonyekutmc4a1aWE1FecqJPU5mxYqhxslWnOOyCu24heVbkcQr0iPVl00OuDI4Ta1OFhvZ0
zxV/0mxzNZ0YRU+ew9K6vL34V0o6xQEJPsj4Xwv170MZYNPSd9qCuCfpfrT0dSOucP/Dxu1OXAru
bBeSizzluvhLMNW6Dp2M5E2zyoEdDozThrP+2gzcVD3LQiXHqA217NHlSaRhf0cIF2V42KtAFcw/
0NUkS6UagL+0CIYhZ61vGIx8uGwej9xP0BYxcff32PvN47BEEZ+9U1r/ty7sRchstDYAs8Ahm++I
LZSg1JyWFNWL9JPMofBqf0/6h0n1vHwO+h1bNViqaN7ixnoMO0KLYx0bBa2n3QS8ZV3McPWoJyVS
hX33vmPMJ/4fB5uITxUvn/x9HponUcWiYNH+E/bgTsYklMHx3Mq9G/WCFG7b6BjjNuDI7A7bBUKk
azatuGsxbG5j1irAj/G5nkIAcZkSZMgO7xIaup3w+nbCR4P9Z44ZnKqDFKYUPRZNv5s/8tMaG2FQ
ych9uKQmcXEvdBtN8itrYFVwZgXb/hF2plMsPxxzvzhrb/i14DfiIraGS2KRkx41VqwTOhwM4eWk
tSl7huc6/pfwjwIxHPen+cZCEo1mrWhQ3z1V+p9tOWu4T+cKK1YAgHynxK5DtPorRDcNd4tWvock
t32x1InW9jjeJAcQW5wD1lekbJUbh/L2m/DiELdWwCyWqRh8IdYnz1tLKSyoSd4yV19+vEOCcA3p
FuPtlRxg8AI9lpqWD/g8st/tMHA1f9Ynvz8BjxHm+G0i0sFwqotZspUYya7VLR/62+HwWJDovpnS
oKZxOXuA4p+ejF/4eRr/E/n2MWV2tnAcuZh+QQ1JYNmWEfDEYreJ/4OODQhzA5jGuyS1S1HS8BTB
Le2UbcWdSQ1WdFlEz2oJzp8M84XqrT8NjerosxWjc+qGD9Ge282J1CXN0rrrEF+exiCz0mpmmKWr
aX+vZrAQf1TEyf7nbDVO/3XN+aQPzxZWJiO3D5zGFvdXSeS4abEWLbqAAqYc+xxKOG5gtNtuNrV6
jVITp6t/doIgNYwOHh26bX4krvIYF2eBf8ZuEfoUzruixa+pA2RfIkMmGqKA9NfmXUQAWB5Zk5cF
+l1Y6+OLgT9MLV0OcBiLhtaLiu5eM1vJ5ezKGxXbpyKOgV+KFL4ENnqOVPrshCCPkIhrjRHAk6dC
IaNSYUo6HmSYswA4VidbXWUkOLJixc2z+AtGTQP0865kqj+Kc1uU0bDbcT5WP/aOZpk3dp9PiOuQ
85/nqo70E4SY+r5EYCNDM+LSi5cOUPCjTvV6LcCEO5vCJPSv760uVlixe9HUTxSsKqBsHt/4+9NC
+PNnWquczmm2/L2fixN7+Lcc6OFTHbp+42+Ac0xiPvshKuHRW37DYC9QEvOptdde18OyGG0wF+gY
mScw5kbpd9U29XBquo7e5u30Q1AEd4mYvXgrzClF4Nl09Cmc1HDWHiP3OqQkZ7/CPXjQFWBLqgzn
SmzDgZl/4uPVGb1OO0ymsM9qsY7XI0Y9Itnk7lsTSofV85HLqJ79d4Mh7Xymqg3cHAYnZjZcr4L9
xAUKYSUNNrKmgcmtc8WLVs4DRMuccc4+NFXxdOhX2ADAD+xN7CDrQsDSdWSTK6K2zK4sIrsYfSY5
IRohds2SRreTOGIXcIE57aWwaLcnMjwB33X+rNaSlni2AkktNn6aVu9YwUUHRkGVRX2wTyl5rscX
hne9gXMd/I8SlZ9lpOxt+0v0UTJiXSpwCCRa0M73Oo3V4XHrJSv7mAxRbwDQ1BJm0D89kZEkxgw9
7nfZYpBylPDHafXwUBlScIEu/s62j2HAvUbucCTt3wPNYYyrRjTYhUWaeXJQAfbV32cwt8GlkiJy
zvVyfJ94xb3VG9lMiNttbKjCtaAb/fcWMnzOrT5yK+KderXeJwgIBx3dx7/NpZG/sRAORTVrzoQI
IxLU3yuafkTW0WFXXWqumDciv7l2YzDFC3tpjo4jDjuNdeBRqaWL3UPOZ/YV1Vx/oPtuxM3wJ2+G
2B05k388ouJyYN+d5aO7Q+11VgGt2mjEUwD98hzq2Zi+ofVFH0Xrwe+nwISj5hE59LOABm3DIOu0
TQfs6O0o6yf2TkiST5VoyPqINsDpCVGxzPqD/ylnhCwr8TAVcuXkOessvXcIXIfQztKyUTW5hM8i
mJKKB9pYcEnfZYgCNmCszFMVQ7LRxqZUiXLDOQZuiskrrEzrfVYJbyhz6jMv9lOCzZ5ahJd39PP0
xlouXoZ7rSeU3mIHhsa9ju6S5SaoudSNTfuhm+9v/WLuEjvj5iGQSDsFE1XkWQjjXbJPKw9E4HyT
OUTfYsQxDk3L+H1306ukh9RY5JcA739KJfgIhaQ7revzc5PcWmgtbXyeIPmWZmULfUHjAGY5+Kz3
NIHUTmioqGyV2Jq6k5QRo5VHCAI90FywqgG4eHjQQzg7uAnLuMrAYgrFNuU4pXFmUijlO3ARibnK
PUsfmvSvUQm2wrb874lW+rLnbNiQA8XEx1EFAsMsqCwhZynPA0WDE73TFnrvyi/X5sSGLrvUi5IF
4h6f649ejm0mmDB/Ua2gTg43E7qXO+e4F9zL8zfpi9gUDAS9b9ezJWiBU2E54AMTKZTKiTuYrptP
U75giIJPYoI1CgN41tPusYUms+bToRo1/njW2CxERlaTSpAXpfNTClQITLCByc3BIY+mcy12UuAZ
nkFnmT16kVPLiRV03selpwRXiCa+W1QO5gKMR81Gh9NldcBw50xQrWojdghmS4P6E7NNVkO0wt9o
bxCalKWviuilyhKw+9LAXGOepKz64zDHd+AZEbr0vuLQjzrGNm5hp9K8SdbbnhR7SeIc4Xv8/Wlj
96jP7L9CTCn2zcQ0ZvxSlAi19MDPgeq6/NnubxYXrxC8WHnJvqcjANTcQ5JLdnJ2VleLQMvdXYp2
InnsQqdEKrTDG9OL20Tz9A2KjtP7WzJoZ3HeW2csQMZCfk9w/Z4Nj6eqL0Pbj9vFkE1jdq/98QbV
6oUcQtk7oImpUvmk3syg1EBOWDUmtpfH/Nvy5VVOUlSEz8ueDW1CxYuODxlDeDPz//3m7sBrMwCK
cImc3AV1S+h4MPTpA0rSpnx+qL2LQd1I5jAEVTs6mdv8NkCrpyhIwTZB1Vr2618q8LL8+AMPEQ3i
j97NmhU+4oJiG2dVNuWKSCAr4IGMdKGgT+uR9Vu/nNgJA12uR5Dp1sxbQHLxICvpqKmiqy6deNyo
0rMTmXqDmbKjW1ZJVPfz+N0Kkxd3HuAT9JmpcovVLlnRvRpzjRqE+LDQ6f50TgDSP36GO3Rzxx4G
Rv6LMgiV6kV1kROTar+vL9lWKhTrZYM05vl+x0Uk1U6ogxgcFAVPUu5SWFIOCb3ktZjH6Wb8Z4KM
+0y+djr7/vPPNQHUsiFZafTymx2PXy1k4kn6HkQQHkaGk0LN3dwJTG7GEaCcTuTBlCeNAPdmAOOj
ZUVb31qeZuRXGHt7PH1A4F9kgY7FazVR48mqvIzELTX22H3SPUDDSVhK/A6amygDf4phZjsW1amx
oyj9Eoij0rpZ2JtNsmvIug/rZWSxUl3u4Tr4TEPiG7W7RPN/YRwdQ8WmK/o+yyPP3THOOzs64DtI
M2snPTZZ6kObddAwlQON17ZTiolqTOL1TAKAoOf5Kzi2w6qJJM7w1fa2NP/IiV3LOA6xzinYGaTi
BvyQDvcJ5dVWl7jHpizeEtcl/muiWpT4oWQUCyrV2u0PJfakZTrYJE/lx82z9YlKihzz5hYx5jiT
a2/NpHjL9k3Rk78AEz/AyaH90Uu5LX8MKZijp/7Y7BjhKvNuwfHK80nXB7JiEG4pxmNpruJmLVn9
vMuoqWFIVKek43tauvjU4uFW3e2aXsEbxjfaDam5io1Y1tEdSNHjCI3x1YIRMSonDyCwZZVlUbv+
QJ1b1HtKBxC/cFbr6DS7iLmP5Zo8t0+GQWPf0tgIQZhMUCpteGc1JpL3kukVDzYnQt6ngFlJpSSC
xhVWRNUnD3wLsmCrf+j/1CJ0YHPndkVbAMxeVkcyYZBu1xA+bqW6rnGm4D3ay346aC6kmll+kwS+
WOes2TonIU/KIMhV1PQhf+6BpC4Fi4wGtnsjw1f5tAmKqR13usqlmDe3DT9tb++Q2SDrUia0QZvx
DTgUd9A7bxltoId4k/Uz9VMRsjpmpdutszmEfmg+gA6e1HzQJuC4t+sk53D6icVKkYXJ3PS7V3oQ
lEIT5p5AwF8XiAogH6d9c1B6YqOlpS+AeD3M7E+ntBn+bOQ7tOaM+26G3cJPj33OuiJyOWR1T40o
fSk01zu2LKVXsiQYcy6bsTSvwG3RpzApSAsuvqvTbaRgYpn91hDS5oeFZYFam6tR3bR5+RsOprL9
R9AxGk/8yNOHzx/x8K9eGm0eA6Nmrts3dfE1NTbLBkR1L4D+HsEg0zWqThL9KAWBBvQcDgFWis5A
1yFj06osoH/z3z6zh3NJqbcyxCyS0cVG7c/2nbMo73ve+/fht7b2sAr9Sdau+4V1s1w6cT2qnyxu
k86jCrpT5663jcVDUdlV0ZrP20rDABNbcg7ybpUax6duMkG2NUVEpFZdiq9f3GDApTIqu79j/0L4
5l1Oh1+mWrU/uCXZvWFHd6+U2NSsGRh0nghfUaURRAzoqCABivNVzprxKaPr2sTO2hK6TvRiDDM3
PuhpS3XIHkfiZEso0rzMco5b7ZDhC2D0JyTW6TcQQZ2NOpEIlkHmMepku+nnPZ39pibWlEi1A3C4
SUBk1cgq/5Jvdj3mXJ5iDsDDsvGTSKQlrkembdwB6EhlnprtX735hhZJ8c0oO63VAQWo/010ymL/
4NaDoWFGnvqGCHxRXWGNXf+9IeCWujzuzHn6i7GS8zb1S0eJK3ITKiKiNJ7qHpiLIGpt63naIsvf
TPCF86KZGEfE+mZhBL0E1PikWVvJE0zUAva+11Z24QxL22yVPagWGx0wMbsm7O4kKOVlBnw5LM5X
qaBDdeXQBEz0AKZ4NAEndeB0n+A2RgH/dD5K47LZQByTUW4XgHAyhANL+ZWniATSOC63l9Vn33FX
idKUwbjsqNBdtEZfLsF82EQY4XSK1tNt+ddlj+bpvymcXCVmu+gBqiCdKVXEpsyqcrBSW50m9fJN
9bD9O7OSf8ItOPynrQFM+NNOpR9j7MHdpNtawwwtCdM2Kek21C4fXj3X02WKPK7XDZMENaNvkk3r
O8jUd6M0FIAH5UbKHwxejwEBZstu1dpriaw6+C1P1lwupoWj5amSr0+rD3sLzpQWQ6ixAkMQznhn
gDDvNpnGek3dl4aemiSrcHAilQ62Rfhlos7FKIltqLpA4M3R1PagkRzhNrABsd4vmLbDCIlmKeOX
kTNaUaIPPc9OO43DVL2pbf7829pzt3DI51wfUIW/MYEI1b8U78HRYmSwBVlkCan2TdGL9lwEeIZu
bNyiP0jh5SVaNsvhQDABxA47f+ilRxLcJBbw5H3Y90BEn8NQTgE5/Avu/x8W1w4yCYS+C9hRg7DN
cgU0RIXxlpMGpgL+5nMkfPpAEcsmDene+UIt1f7wlsTBlAxbTxOmDgrtfw/0oOOSWmycES0sIQtl
C9hP1Vw6RMS/xxt9VCR2E16rGyf5RvAftYy6iC+s/VtaRh8Df4gkWGWHb9Hhfg+gOjp9i7b5ewYb
7RYvO6hCdcU3nIbl0tuvdEwYN74x1N+T65hjOqq5Mi6qC9zPNYCf46g83hM1bpAeitcDGHw5MudG
O0I0CsjDg1aSQdZy5Dahv2uorRJjAPS78ZkkoWXXi5w73jGbh4wubxTA1kyEX/8539W2jy6oU9Yh
mWNUVplvMge/6MyX7fesGe8XArN/2lRKVOy2juh5WGCfHxJxyZCbT9kOfscJrATzmYFyDYAoPaHS
a/qFqRIgvLeDZ8YGy1HRv3c3enI87Vow8FI93GOkMXFuNEqXavKX3cRu0ztz9Na9EaEeNDBgdubx
dkwbulJIuYECbQbC+e7o9Sy/IjrYfRdXsTmHOJZWhUk0FkD8fQnv1Cg7Vda8GbXOM4HRM9gwS3hH
JYUi6+jL/Gw3wUYdOtdyMpnsenHbeuKYra055jM0Ywr83dcIhNYA9LOmq3z/C31pVBbAqBQAmxTA
F6gbRuHsKUBjKORZfkpv21BhbYUHU9b6QBO1WNzbs2sxUKEBJrw+XliOfoErIqyvYHZagylevOKB
1TpRAZn9pRiy4YuwtdINYtFCKPxijY2QV1AK7vGXhNYHvtTuVSMrtFsmQsjBz7WRTqPNLYJGzaCU
T+Knj0Kkxl4m04wVjiUZrVpeLZsOaUdprkCHiid/WjJQYFui/N5S8tDgUsQoJWXeYglZg0nOTCnp
2ASb6RFBKcPJRoQmqV6LH4FmbHbVHIUTc8uAfhh9khFxFAIsMfg8/78AuOin2qr9nnwc+oUL4SoV
sEGIlwgk/X95F2QDl3Idh48XRUw6sizQwCRT21k4iT5D7LEhA3umQKj0Y0pJTmR4N2Hutqc0FEk1
UdmrZMNnfx6Mc7r/goo7fDtzzEx2aSgGhZopiognl63Dl+IAMmaopuXM8nfJYp8V1cbgIlLgh4VT
gyirOR/Kb0fX1o/OiOxJ8D58WtuMxXXOiBBVZXS32roJpr3edaq+Ixw2N2EXONmK+JosoFL62WEo
wg++K3AbNmMYUzWQ3lywLi7E2ILdg0Lj5WCaEw0ezmNhKUp0V3uv0jRn4X/tJItvZk0iWf9tNAJq
G17oqFCqz+/ubXZwZsCK10C+6Ssm4pz94lTYCp6F74u1IwTCcd7lRFCPYRTYi4QhkbjYQYMYWMoQ
sg783Qp8JLSPVySdaTAtDqwDdU7b+/q2Po0fhn2UAeuayQvdaNwYOrAFa/2UsKdfKvMzA2TeRx0b
DXGzGalOyay1X0J25gBv2DPk7t5QW24v+w+o/n8u9fuP6SEfud+hS6ZaPRKk5RPCt6xjYFp3xITW
UCruWGXbTv3fD8aKXcEa3mwE+BNk6GWWOvjwLCfWULU++tw+TmnTobjmvMZeTjul1bvnAqUkJjEZ
t3/0lJCjPmi6nPIlhJ0CKYJU6CHUcQLM++nUN+uMEHaBq3Z77uNJt6U8824KGhsT8uo14PlWKbb+
qIdkeedGrBFLND1eS6NtIcqsm8ty3/rW4diqKTK32xS2OSuq908SZvRUJ+2sYQVHXL7oGhLWf54P
jPoCyX/br/V6nQIgm6x0SBwh500GD/2nlPhyqkAykcKTCj5VWPj04ecVFsC3hylQVtYv9B/yrkrv
fLuZdJE5LAN1mDljjqg+uWHzCz7A2sLyk8ZTgtyBJMynD3+JN/3qVMmLi18vHSWmogQhPcPBS7ks
jAxAn/Va9RdakJyuDpQTVPH+XzyoF1sXiwWHzNFuBVLup28k5+frev+9iP2QkVNmsKvIyBddIy4q
Yz4PX++AmGljeEaTjWs1ZSzK20n9iLHoIhcex/t0X0B2JuGFqYNfG18FZgxkNxjzosWWyoFBGu2c
P/epCzBJW4wvmN10qnXBn8GeqcK1WMyEHWr8N4zLWn/u8HOp4uE29mErIpPSC3CK77e3uILlsfEt
5zg84KGtBRUsZjK/Vqp7a1/ZX2XRlW1lt+kDdvwRqOxHM3l6FWJntvUsQoUCq0bwOl6+H2SPrjNv
dkqboTyldcVykzfgsoWS5DrtaCTC6NpWMb7i/CwqXNVaVZsaXddD0t+CIOjO9bkYprJv/+v/koSk
cUOkZvMN4ksxX3CGUwF7VK5Ua6jthPXU/0j1yIP0ff9oaLRH6pIH7YbeGgFGsA1xI35GGSUCKnbc
lLSVv3BU9b/wuJal2kuWfN0fouHtrgWTvrRUOYLdqe1Kc880oQE2VRHjb4h9SLzy+DmP/lWlmtZR
1j0mdcnk3d8OJOeCb1uDwMf04HOuyq7xWe99lNzSqWARpG2FBW/xOwdxPZAmdsBydULYhXpb3KNK
SM3/8IeLb55X2uaHjYwgWH8q91cr2ybA4uBsgsOOjDdnfNq7bFpiAerZGrQFLvsqzLeus6CUpnah
13+ldoCitexzl3k5eNmF6wAEmqvrg/cXl0UShFbF3sC/aaOpnLXZhMAeFES6ieFQcjcRkSIRRRb5
AwoOsRMcp3vC6ENTQ0+50yLyCR8lsdOoAHHga5T11Z7dor07NZS6YWCjR6HODnG/jTvPB/v1NukC
+LQ9/2m/ZfEQcloBGxTpdnft02nu2AT2HmzJsPn7V9vJZ/PwUdo8qIwridELdJ+cUSvynyemd9qc
otdbnmMvVWAOhfHHXuMRJXWR+tLPvpu06BmejxR14MaxJVFeh5SrdziS5C2HDuoXbaNCGdES2bMz
HA2/AnTSCdHOghTL/pLneQFUa4wtE0rG1qUA7aA1Ca8IMSadglGKntrR/GWeqWUrmDDAOnzrBuSD
vDXZEjL6cfZ0y/cOPE8ytVvIzVy7MDUz54qNUVF7xDmXXlY+P/dIzwBmYwuKO3Jz2m+WXwSYrXjp
M6K+WE76XACYKcykFJlIr9XMbDNF3fgje9tmFe+YlRhfcK5sB2GGBKJNAr0YT1q1Vn9HkTa9vIJl
jbBgFmFKTOF7OIEfmEb8fCyfk/iQ78C+SA9VFkJZkmDyqPjBmapyUSxqRAXVckJKCfds829Knigh
Qw/wA2u7FK8bu9hwuayLHb694gDaFB3VFXHQupe+qLw6vw4I5JEoQxIpnMrvNqThQI/rvPwQwcQu
OIi+tJc4MnSAdjPWQPgnd6wXIxjel7Ez9e648BtyVyIqsSQnQU7F4dbkJ+K0RGlgv7CpgymRoG6L
80/D2yhUEb0Ng6ZdSQmxWlgx0kv1JfGCAvN64qfQxliy3FxGO+J9+BuyOCnc8afDppAactQQjmlW
80YEcTofgE4zdgMLqCuHw9eD6jZOAFZDzhD/vBC3JBIoeLy/kP9KL+jyAGiMtImu49lDvjCbx+qN
Fs/25yHdjEdPw9ojBeOE9h/cpSl3XxMCfzeVAH0IYQwqXfAcSk++VBrsP4WyzihHz2E2fWC9fKby
fpKOMN8Np2D+xzkzj2wq1iqY58WuYd+OafiN+5uSZCcdP9lm+iONEKBV7hYg5zmvmvLx8R1tUVKl
f4S8S2Llq7UDmBZrsvLkyOmn5ARTjcpVoXngxI2QfsiDBfq8AdaF+djZnCgBdAL6MgdyCc/ftJaQ
xFlmyxAI/YNIN8pwApIRo9hA/FI1Zq98i+biq9JuBJrls5aOHgPpgdurUlAqFq+Ad/UFpgnguAv5
1wXYEYNIzQS1o2hWbDUZtCVgGAwyAHY6c6h81z7xyvEudRjnqZOF25Q/ByFqX1rCeFrFp2YAM3d/
N9lym6G0cfB+3Ek7fxcUic8P4qQIdKqBPcsg9D+HDWsv9ZKdWJIIQp/Er0Lm5mflhhnkS1kI3zv/
6v8SrEzT47M2wsGxoxkRlQ8TkJkpEwuI8HnEDgfNod68ziHvhtVoo+VU2g1KeVS+TCZI73thnpdX
SwT4FrnFOwlLggCblDxiA6+CJu+gZjV74LLLcfIkETsjTb2cHu18MbbW19c8Aaa3NtHvX+9/GP3e
csUWCYmwHDkhSrcmAl9VPZKDS8S3ULeBb0Z16ewSRDWyn9CLL1Jg5FuemQKqe2mdGQfVhjjUrBvS
WEKrbjcTD1mYxjYunPN3gKR9zPtBRPYobZPnzb6UqeBld5L5kk35yoLryCfoIO++mY0YsBslJNvk
PXFtfV0ZSfahGZTqGdZx3rrOzPq71No6sGIyX4ZI/2H7NyhaPk2sK5VHu/EnTCJMuofYFyB7BxQa
gH+hX5uUeX/QAVb8klFVQbvyQ0vCnMW3ZNoO9qRB5ROhQ2K35AkPPCYvWwjO74QU6fZF1diJ5ATP
+HZ8nflGrOKBnxQz2c9ctHnBM0TkA8rmgkpQKR7A87H9V37sO182I5nCQVtLdTQePY+AXmkkWWMe
ytAjXtfxXk84Hhm/7DQTpb88hyAJm6xjrLyfvFlFIG0XEV9OrNvBE4JuQaIZ5nKfa8kq2UwxznrZ
fQ7epBbVnhrDaeFHLHLfaF2WGPqIxflIJ9b6ajwHimojZYGXzCP1FYqFfga3z/YJjgZJXYjsHroB
sq1n2GU+bWORdsD33a7PD3uh61uybwDAO+IX+ReNveuPFwyeJpV/q3cRWIu5UCLHV56XRz0NRJmI
dd9/vMHvLwyR3BE4aTCsCJzR5U4+06qUp6KE/BZTT2juh4qlzJCYmsosk6DBwZqVSQmPK6/egtkR
G7rWuFsMRnCOexG3S4lna0iFQj9HbvIQ+yqNmOKO3K2IjpgNxC+FBwkh5obJ4Y95Bu5Fd0hTiJYm
cVE2KP4C6aSzUtL2aq729wrEL2dSXXoBAPp72EMuwJXqFEes5G3uo/e2h2zvTmeQJh45aibbRM6L
PeZMTl5kFx1Fm14cKrDw0ggJzAwuRnA41bl+le0yE6mPObw04gzfTyF3DEFm7iSk4+aoP5/EAWhM
1z5s3prdiLeonm5fP3JnBOm/VF6qRIKsFwti27zt6dYbChK/ddmc5w0xD17gBgHMKgmr1nS/LZKA
a4B8nnAJOFrZirnTZuj1utNM4EL4Sf6F4YRm2RCCfBf22BoP1OZh/RlhdTiqB2O3UEMNONhiRH+Q
jjral2+r2rfBqRKreNNKSgA0IXjLpAe7vOBXduxAY6qcMXS5fjVk6hxi+uJMubjyQ/K/SObiLIHq
ZRkzWIlbMpUzuByov9r/2e92Ssbod+X3mVkLna91PqUSdpQ3zgqDsaDjB5o69pOVsBPuo9NRqvNf
FRbNzQ/Xdx31ncmL9XMBhTrMJ7CfcwB+2FiWhsx4TXzSR4+5A5Lk6aVrLzTdcW9U6UdFJMAv/Q23
MlC64DDA8OpFsuT5WmuYY97thUtp6s3F80tqTP5HwGe9gL91qtm0AYWCbxGHf+fRxqS0eyv/8WXf
5XX33fJBLcawZpgNlY4hzH7pgyk/5VV4mWw3Ea6Pg1MvjyMncG3MW8L2crXadf4c7NPrhYhg8R22
ZiVAQkhKJTeeomaQ1XgSo2gBu98CxlQyonBAXnM1EWl3/cTG2iNWwaFpZI9eI5H9bRDvvtqntaak
G4RfynHVg941YSY2uwhPgQ0/9RVmkZPm/xnLDQ9VtzsSf0z9bPBx/sv9CyOQpe//zXwRIeCCQkAO
Vn0m37daxZ2ExftNf4NlFhwEhooco5ahod5E0np92IAQ8hVUpf02ZFKGyPRbpnBmLHL3Ry+T57zC
lT7xsGEMnr7FN9m7VkiX2RVQGTC8bN1HtqojCJcBSFU8YMlS9XFxccnOOb6p/knq1NwxzSLqHbpO
MjaXRm1bb/vV3ryZ1FgmplIvErTYGuBHo0OmcjhASBDshjq+A7Fes1fjUMZxpmS4cVFuimaskuyQ
XGBlGysGVmHg/whMRUnkyncFER0GbVnfDd5RSh0SHmvHdU1uhmy9Pp8aq2lfjGoofwf7SpIGK8W7
vB9Kl1GAzQvNRyS5DIG7zQOVlA4igAzPVeIsCT2Yg6vKMdupllLWgxAjGh65B4C70urAIhtMaAVu
FOg5NahsYcEJahljjwNSNilxp0bzAHhBxD0slQq25xrf4xzIgorcHSlc5kqlBvEO/ljS5zHK4ENp
5u+vWXwetMZaMhFuHd+Nidv1+MYkqAN7JnDnKUPzJXBwhNqo+WGxQx8NaO36Vu4WoIlCRfcDq1Ny
NT/qqSSHtqneIl4yTcWgdShX43K/OmKqT0YYgbIHRCwhULyVLP6u6tsSbVBDcrq8j9nvyYbZHB3J
LuYxh04h+bSP8wOJBltbitH/Dk0bZc4ni6Jop0X1rjrF3BdCXsl0R+vloii8Et2zxyxu+UY+OM9I
buWOee/P/tW95LYWmhvpkzbG3aKT/CxhPEWfe6bzv5COALGq4FNQoPBzMoJY/i3D/LHDhZ+u+eTw
Aq0dHTSEcZtgdsUNptA8d2XZ0CV+vcE99jxSWstYMiYvNjR2fE6xDvS/Lt0Q3vyJKk5moPT2MqCc
z2uRIHnK+SdWWSSBwGKDq1aMGYPRyxVbXdh5Wxqvd9nLKOeWc+FlXb6xOJrG+aUDamuaK6wz0uqP
7lNbYrocyjq23FEqJqS5iwt56W2W2aspaCgrjbHmNuFyumYX6URpaBUSZe/2UU4Pb6nviguy1FZj
HqAxIJQSnupvqyhhxOX5EkhoMVTlnDyWfeX7yjOQRrisKnvxsfBCYwdc+T782z36ylJU0IWt5sbB
u882TTqa9V9VMJYPV0DXNtAzLY+4PtgyBP6wj7/aU4Gc405wWTh5jHDuWNh9xqkJBkhAfXRVdk0w
bAO1jRITtm+nnf3A3GaC8KGyogyEdr20wBX6cDkykXiktkhULM6GiolhrTLDAz5G4BaZFBbwKNAH
N7nld5gSZ38HFuxgUeuh6rSpGZkL3oQcRfjo75rwEeqn/BN/K7BaIspVFuHzahiFlrvqXUNADnap
3mhhm+ewh66Tb1z9gi8P3CgbP6t5EmKx/ZlTHHx/fjYc+5tnADT1zNT9VsckrZxaX/Mz7HA7TAfR
11cfXhWq3bqdVR43pzfKAwlU5Cy8L3Rj6JrNSGxJwQ0CIb96uaEZ8m8FWZB+7f66wIw8pt8G3IMW
nvVa6KDXsUuAKMy6//TYam+9ouga6SelKVxSmTar2ap2jfbGBdFEcWj8sgAe/lg7yXAOUWyb35y/
0ZqamlvWiMiNGkgf9871FGWI2fT48H7b/EV5/qSKE21Q7HxsDKkuzMNSZ+Xn4xcgKwN/qHDh1/06
67xnI19sMpVudvyBR2ugwGs24NXmsUF7yEH0OWy4d9+4KT2bKDj6qgIOtd/EaAx8psuYlfhZJ+Oe
t8ypNteHmOY75SVPVATj6J2BxQky7vPbuxhUP8bSB8QcNXySCKlV/DPVa5OXm6ZjIAi4IqbDemLm
ksCYJVYDFtwyXVT6d6cwweVpns9kxofc1HOLi7Be93hQLg0HVTapdDfbvM/7IVQMO4kg3cmShjUc
hDHzU67RjlqWxVSDTciJDWJvIDwL7a/pgze9T109awBStOPmQXOjoA73MdA56Ky080cTizEXiebu
MyUqX1eTVrIyUJk1VRpS04lM9D4iYXEvTrIAPcUgVBGUmXtM85NbTO7NbFlgZjb7ZvPsPiC7cGDq
aTafMLFtoD4o/c5b7Dzggy4r2r/f5MuOscEEBaetZCyOQ157keRVlJL9NQgKGgr6j7dWRT9p+GOj
gfEGaiSdMSa9aZFog0aE7oAV45G/4DFUJ+aGCG0qhNlaRXecsPlUYwZMRv0kMDYROcuTUBKUESIs
6Os6MIA8Y2Oa2PlVwsdn1lvGtmu1E4JojoRV7LlmzoF18oOIIYGtObhG+Dv/HRoakgrJ/2Y0kPo/
adBLhWIvsOxwc/i0RSAmmi6iSF1Tz6mRtY0FyaWjaUVEpd1x9GLneR1CDYVcLCd2AueFDod91Tu+
C/JHJYzMoe+VNow55eVHZ0IPG33w1457JaeTFK0hmzhRuUBjE6cfu6f/cklVXex8ZUvNUKdW9cBv
fm2Jsb8jeIGeoCatAZuu3m0rrk3REKAhgjRVdXqpkvcHhLqZF+Wnp0IYN0W2NMELtpCtDXd2cM2n
zMxwS6Ew52NedkDFvG9bnbEaq51GKFnYBuidHIlrwQ3Gz0O3014pe22pSZ1uSQDvXGBbkMZLayYC
pc7JfzeMmqru+dW3LsZNp+wqNA0uZsRIpSnSyMcUKZFM7B2n1sze4i3T0RPq2PzV3mdNubBBvqlE
3uBLRb1NPuIkvvEUqWDL2iA73bJ2cLMj+xzI0mg32IUqb3EkIx3qYGtpAFzLiN5jQBYI2ku/1oaS
3HMP/z0E9DvZZ8uDc1qsYdJONK7Jb6fWNsRbspbMzVf72lY5UdhImiINrvnEjlBubnJem+XBFfnX
vo+GJBoOYyrkIQ9u56nH7OjpBEas8y3mnnpKKR9r8GVnQLRK/5YBq0iHt1JxshU0cpngjl+zDTkv
SlmqTjBgWxr5F/RmiXEoZxkfJ+jK/gdVhNJ6nZ8AYGlIAGZIXybXkrSBxD25OmcwQMOAuOMVB2sT
mzsp+m69HDHGJPlGkTOfymNUVP7jznpH4hjq1ljOAEzq4xTxZA6FKTf0Pn2XvMd2R9pvj8f3fnQT
hltbR8elAc5fWawZw+dzU6p5IVNxK15b11mFJv7HoQ4c3/kZBMrkdhwidnJt9wi3w55PQeaOZEHr
EdGjqIvbbrkn3dsNNH9LGGRapfuNPcf19GqPBCwVZ/myS5+NyK2SDg2OJC98HNjbD1KrTAkWMVGX
k3OYjf1t2HSh3EjOG4uX8nBFR0yKleiV7s8AjC2oUzLa+lzhqbZfb3Ww51H7VtnYXvP+4MN08PX8
E/yfMSyagjmO8STqju5G05s2Fl+cFL+t9c7oqcJ2zSO2QtuGyKzASxJTcfB8dT1q0FyEftSe6iln
6P3Xy98PavRiasRvspXuOWCtZD2oAXeLQnGxIG3Q14MJfitPBKjV+oDGr6Z6v69FCJrlaohZeEcl
abfKC1xRd5oJwa1Lvx50lksPNF5BjbJDqbDNEB+pViFtf16evyUoXqSlUEQl1c4+TvDd2jL4sx3H
0pZaDTQQe+ktgEaB1t2N2anLHaqP5KZHxDcwBVCSFNaiXOzhnE82HhEBxP3b1OE5FAVlmfvqbnb4
sv0wb4pS7AorK0yJtosn/IraHRpqxN4KuX52G78P7kLWxbCyKgC2kwo2mxPgRlGiSo399aMMqwQY
h6XfCcErLm6t55Gc7WqVXwZCoLbVUXgBYJ2R+s66ZOZ/lNIIqV67bcDlwEc5kOzHx1renXfOFdmU
xCtB54A9WbyXq6BZpkjnmMd4uidT5O0Qvgy6NuOF2CZ1AB3RGYA6BPh/mXD6Rc26TEzHw7/nrpSh
4W7plbwKogoQ+6j6hbyJS5j+xxAJ7OJAjpEo6JUfIhZIfZulGKsOljq+ZC3kRA3v1YNQtph6YEMX
TloxszENzSMQ43hGeb16fBCcDRFy7M+391X3ByxdvRFTVRVTF9yXe+W8EgNMAj+J2HIu87FFY0Wr
DwWnKyrck1HIkHqjICn35F2uO/6o8L8M0vrX9NN3OvKJgI0BIYovMp1/fTlipM1IeuH5ogRmQf8T
0gUR4H3DvpamGChCC8p6QAcCByv4q64qfxBaSvMofUF6shvDe6H+V1OB4ew3rvyXwR4zBUQiOioy
7U58QyZN8lHd/1EN2X4rnfPW8NWTZl4N7qV6jmJYPDbOMRL7NlsMjHL6q/B47A6rbpUN3P1pdGEf
pY/rxyowxAtO8g22zAN1idzQhCPdGkCbN4zAXCmcOuOiH1APx2mOFmF0qKAiQsgI/Pbvt7bA9Y6T
Z0MhWujtwVw0xIhUZerBMM5x/5VpV07WrSkPnaCq1/I+71uGFdT42GdceXSNjiu41IU7Fra54AjS
YD23GdcX2+2ej3fEl7MrJCksNrfAjnTQVSzumR1qok7GAGbBKvLrfSbRTp2V9CaRLNARgZpmKMwG
fJnNjD0Acff7J2Mv6PbL3JHTHtxNrhMS5Nflz5LLU4LEhRNrobfvCm9UoaOJeRc8/GS4G6LsR92J
DJ1Ymu6gl9Or4ik5155LBnbAte5ceG6uypZjFoHqzQIga5ZKi85NrgzexbmAhqemsOFGmgdXc6xu
swVKyoBMZk/LiCHT/O1R4u0FDfG4Thz1Ggy08OYBSlstdyV+h0CLa8MNKhpmE6LFfsCpfedRqxvv
loiVQm9B63Xyzwkk53OE1OXZ32GmLAi3ej/fyJlAfsGskf1tfagQkU7qqo6T+sqx3e7MWDmxPJMI
LgWNpgtnwSADh8FLDfsbjgY3o3B9CNQr99noB7ts+Gk3RjViv3B26DRRJ5EQTTjvwXxIn4IQHk5S
Kgqjc1rUHWIp/vgrq9FGPNrr5FM/bWcdpopQv5kY8i900XrlCeudCyL5NgHduduC6CvUAX8RYUog
7P3SUd8EgFeElBBtfaha3cFUuxEv5jLxzYfMBUCyl1BXA73V+m0GvWP+9lBsLBOpppGrZODOc3Tc
0Ci6u5/kU8QTSvO5rzRh8+v6hHDAZjdnH5AAFnQNmRdysBm+qX16sLnWo2c33Tt5dOkH04jMotNZ
xTUDuyJH97HXERoJJqxk32WZKcaT0uV5o5d3BB7g0LG5pizCPns1gsfIsNFI4PnsFtKq04oUaaw2
+CK7rQHRgL0VWdQOnNWNOXIgzoQMBTj1c3D6lffGDbfeIR5VvJnBtEUVEhK3ttoizHcGXdbfrKHA
gqSCRAgBj/ZHuKpGleX1oPlhZZ6hQPJcUOMNts/2c8vcVdowYtZrrWMFzfU+mYMkgWOxTM0UWQC+
m+QmChF7P1LBc8lPVifG4eXZC3TpwjkOzCaqLQfEbH3omSaVPk80+gRQU81WZ0bMTQwXxz6a/vk3
0e3tGjldGq7JQ6Jl8SQXD2UXKX8iQYBssr3bkdAuPAOVyKyo5VgC+Vmj2baQtQPZ5H17+1nYiIt4
3IiczkZzySCpSuJSKheA969dIfbWmDGe11wHIbq8LZhmiw84aFkbza9aGH2SaNBAWcYEgzdYzQv+
CdZUKWivUfEh+WVzTVBOFWdvaW36hNCHJQqbx/HTod+gR4LZ9+X47BmWSFapKXOs6CD/f7JkvvPH
rG5WpUdbc2wvGiEc7VmoK8AA2IOwM+zaKWxNaa+EmmI/44BHQtlwdDpvvOw63EjJwfJ1xO0oRFel
GJkRe5JTP5HttgHVMw4scEVJmutjfCAio6gmhl3ma+W3UtUzc6WquEv1o7JIwlcHkBOyAhYk94Ue
rY2kp6I3Mfb+2EpBXanUGSqhDiz0Vjgb2bZA14ui398CfE05cL9XE3Bz+nHY9ZJV/Ko5EKaHY7jS
YH2txEtf2EROZqwKsuDlsTTz6Nyl+yL+pHIpt/kQDPpte9bKbvmXqaqTbTkpXqcu48nTtiSEAAf+
GXvw2R0W3a8T+np/stZTDMpv9W3GUOPRGh7fVBl+A1TcIP+KVYk4G8lzYnRPLvptlUorJtAQiilq
Z18/2KQ1pFOarrxDXfOptIVmFm6xwSloFp3F7flx55zoFTDcszRPzl/eZMgtypIUeUPCnXZxO69I
hUCGhxg7DyaUMCxU7V+Gl3tped50bZb56lhW9MUq+j1HkadOivr3orxRFkGu/p8CtEz9o5FoKHYp
5ei6BGQPstD+x8SsW1g2JNMpEXZv98FY90UoNv3jvByg0Eq0mwWU/lqBmsIHUYsF9P/mxcxocjzz
VCWK3AneD/QfGKcotb6IyYjudnPNrYRdNxAd2yYkdTFn1KRjUszSZRLdm7OGCT8waVww+v1DcRTA
/KaQNe7VfLy8fTYa2COn3jk7UeaqQMQIh9jMf8ps/EQJ1xhkCzQuBRgstlj5Q8PFjXHFlF4k0uR7
6IYkO/LJhLO704dBRygakxyRJKNClEfSwWk2uTWjMI4dsoKlmxuxRTI5TAr8ngBH8Ew8R+Vriui/
7u6CSE4kdXUvf97wACbDg+8zFbiD5jCU1pOrEWzEoTVXa39j4UUa6rvq03u1L+GyxQAAE77Z7aOJ
mUqHqp6zKQCPz0aLUEqZFVkGf0brKL/xawQxICXOZQLaNLfVyE4tSixwMACj+ViZTldhw+UagYVr
og2gGq5T3paXRp210QIqsUymSP+4i1uESgfsfUxhdxQ3+lE0HWRoiGnWibZUiQCXN3Apl9TjVCG3
sG1oMHRnTxtoa/UvNdgYD3e2MWymfEF52RX2pCTF91C7SEp2GZJdjkHHIfgjSh4lx5ydEla3dXee
aK0KjyIOJEeRUbmQJL/cE4BTr+jF0I08MM1b/g2ooLzS/u1C37qSb+XIWTwUB6GAsJ4omLBAK2kP
CaAMUMMczijoYnC8KwVuiElk3oxVxDsyra584+OaxvSpj4tTpdklwfgkKveKSAzDuxtx0qLJE0KB
woMdkLdnF28Gvuh6Y+X7Rup6KE5H40FgHAR4jcsrIguCcteq3XW3fen1EP8jyV85u/JdgphMGZSL
RgPfhDoWERVmBYLkfzku5uL8AmBEk0J4nseHZR11xqciD7DELdju/YMekK73SUT9H6f0CVi0tq5F
Hx0CurlydDB3nsfx0I0Ov9PjDBcOGsOTHVtU3aEXk9mmRc6n6hjpOwWSrfsVcgeX7RJOXhHFRi+C
2DwFcXEI3ayXPsGVrwCeJi+33CzElZSPNOAeZeKX9mGxsutLZ9jP3RgmZ1D2vJkWTeQa/dRJH4Yp
Xs1ZnNBXlB5C0C4VPiahobS+bLmdz+vBgCERQtxKi0dfvyOJV16hLt1EgeQinz+GNh5LDJrG1vE9
T1MNqKaTV+tGfejytVNL7sNpsEyAlSGmIQ9afTys+Y96zK2ArTo+O/JBkKKXx9r7WMNHMHRx/yUq
CGLHM24XM5Is67EVwE44p12WMAt2fUQ2r2RNanVEEODxOaLlC3BEc5FmkECKTOK/ZzhJPJewCg9e
clL3Zz3INHCY8k3QblRXVFpMs1wMHIadzO83T8UwRVaHlyP4/xYsE+J0a3u7zW8d6bzb9eW8hBbG
KFnE6fKtLXmy3pepGP4E2TybuiEdL/y/Ryy9sx2tXdIe8YF39VoqqAxLoP/gzp1ueZWQsBUJdpfy
xIbJQ2TJz8S8YB8w9FENCPna1a2IOf+Fs0sC0ayWTJex1n1zOlXLxsWu3hnqJeRIaw71i2SaSTJj
9eRffTb4DGF4hcsfPUA+gfX9z8nC0UxxiJQbb1LPQ0nRDCZyrB1Mixun3PxNap6hdphLkYqVMEVT
xd9EMlvU79ELNqEqCDwHTUqdJEmK5p0yeHJ9rGXq2TiaEcvJbaGWd4d2ViIRePElDLM65wsmVBeB
qA4dQIQFg+dPsVB7pybxDgqdXhSJ5WIPVQJmx8uHoehNUL4rTiNra0L9zquexT8NWLuoN5LpwmjV
6OFU2Nf5d6akwc5N13Z9od1ICEaJadKUEDrpnSmxVyxzQnhZZBB+cqn//swiYeautJbebj8yukTP
SziASxLrYfcK75jpTGMUgCdcRwYn3W4Gcedhgpczy93lE1qa/4HYzhajpSvYZPTbyLqhjpeixxXW
NlTrhasqqKV0+YX5q9V4YyczspM7tp71bnN0eqp2OHbW0E+TmK25MexUIw0XNz9rrgptFjMvpXZi
p8uppYb2uAwIaJ4Z+7XZuvp0L414VE9QbbwVY6uot3vjvhv5e/b4z4ILllfMBmH5Yl1xM/9I6qAO
HAAZXPq9AICe5bKl4Y1gXh8rB9/KQgBy3Zh9YXX12asAqk57D33iezdyAagcZK8LbDfyIkAOK4Ye
TUULEXgdrX81OsOLVMclZ3O/6OzNvMrj1jphtAKbnUAl7bdhKlql5lqjCYWtfaw0bKTgy6pVPnU7
Pi9Ug6A8BPMPkfsbu94gBI9Z2UJeRojOKCT9phsM3nMq/eAn6muFqtnOoPUUJIVMH9Ys7qLIkWPc
j3YmDSi5Xr4qsl/JjdgXJGiVpa+i3bHxpdjD+iYyNwKc0D50oZIEJrMhid8GfVpW0ZKaJRqnlkLy
vhkFqGvKwCkIeCdv+/Rou8r/4Wu/ZpIChJvv1Xiez7D1jyvcShLyyWdKYh8MuaFm7dKXYpA7uMKK
I5RHSuZe5iDeDt9oMTPZ4+aMkfIdNwuGjB3EPBxq0V/+rQ472QOHgKSN2dL8S0yD21QafdlnyeiL
ZOp830Dab3P/ajIA9DITs3xL+DaDoooW3lda07bB1rx2d66g41vVWgrrLHSml5CeWfr8mp88z09A
aU5ZBxzN032+3WOJRSQAPzJ+HME6P0/hPuy2v9FWfg9WFD3X204/W4OoOqb5Mf4uflL+4Njbje2/
YZphrAc5ivkWvS2eE8lqJhZErPUR9IXcLd82gnwN0HgEjd2l1xyx1kBMcWZq/2xIVBfSkn8EWlwH
z5kDibiS7c4XBZtkQKjKzw2f9x1+K9n7D+BD/3FLsPLZ3Ot8ueivOOZbFUy5CDq+qVnXTd2sSJvB
S9vqKw2T4z39Dy/sE7MRp0eYd5/EI40XocdmXC/WOC2Ju4UuRIQvUqpIzFyorbdYStDAaWnz8tpm
WK08X71u04VjiSMydvgcGs1+rL2lWJx1gnypOOKZKZ6k2toTDKdJhoRva0EcS7Zz8s3jK5ceSc28
mRIkY9ECGYb2gBCqn94yINszd8d0Mb3aGajLVrnN6fhkVfchaKz1VqPck9sq76Jh90WvNHgfJjNd
wK4lum+6KIayax9tudKEq4Mz9nsHD3sXu3ZYSsPZRAt1DFIKCS0fIhBH2O//FxGHbc7iGmAhGqa0
6qnuD1QFJG5YlOq7/Dk3n463zMMnsErIfEE/O2i8a6ajwZkjBHOGZWnegnx9d+mGDgdTBC3dDvEV
NN4m2XLKkf3c6jW9lVnJ7+JvHhFutazhOfAg2uFA1RqgvoCBx7ix4O+8tbdhOR5d+8sXyyphxJAM
VHb1UqpwlejEkUKcJPWI7TpLRSJjC/HLntGhYg3dradYF4Ns82X8tgu2GJy+oaIjhLNrKa7tIJ3+
wp+7GUSPoJQjZmJQUjjqdqDiDQRHlh2rx5to6gIQYefqXrtXID6bE2ZW4GDjH8qJJ/UH6iZSs8af
UxDtTVxGGRP+nPn6bawXZTY+VpD4JHB805MYI+xNh9L8fsTGDg4jBEh/ZnkK4bA7ACC0hcYa7SVB
KfY53kZtEtOFvd6hkBjlH9PGP+JHydcTc7qN3PwV4KhZGZcEvyDVHOzl6sBc6cZpPc+B8ul88VnJ
vv4/EW8PiEQHzc8WC2RftIXpYopsk8OS+e/rKh1dJgI5DGVcfbOquniPSpiMqZutG8CgyOQqW+jG
RokD0E88+LiRIJqoZLNblct/rsbY/siqw7iQ6EZ1Jhn5KjZ8ulpqbnrdErNpds8kHoUYMry4uShN
p9wAd6BVvZAmnnjaD21wr1sQBzWuqaSbHYJkt8wIuY9e2z9ebcFgle87Mbb5iDtOBI/mVSnUFNPR
MBQ7EZ/NMV7tBlqyUYLvESniFZFxbZ7Q/RuAE6ZCbJoltmMFo8r4YpV7GglBzCLTG58/WwoemPzr
2e52h1B+ahDBc4e8MMtKUEAobvPIxkgG4lR+6CWLG54XTCkomY75ZpiZ7oWv4VZG1PYn10F/vPTk
Xe/rS1oj+R4KT2EKmHX7ILF7JE/hrh0Oxa/Q62qyZCtmFhSqHUIswOibnaBCIHZfLv1gy1WSETNl
HE7I52D0vYfZkQciBS4zTFDzRB5JN7+L/jEWHl/oC4+HhEfbdUqXPPbJzCMxNqKEQQldbTWvo9dS
xvhSpUDg6bIu9b1SuNd6psz9xQPFz8jVil11xSM80xDm/H+Q/NViqc8Hg/Bn0GRq14bDdoS6EcC4
G6a+VrEcNtZSmQaDhNvAL4qGt0kB80N4bdiiU7t0P8Ud6TuxiG2RnBwPC+Nb/merofvwkHaxTDKg
2uXW7qx0AHb2RaJ2ktk6bm8TXoRBQnmOVimGcr3IRBe99117RNDJ978zN1dhbPMqkb7WCTS6FAv8
fr5G/Ekp2gpTSXWcUaCxDG5aZEl8cVzCZO/IuFviNrRKBhT1NtDQflmctNzZC4h4Mf4Tz7W86U1X
eTauo78/4umlLZBTUQRUsfZEfoS715y0fI8vWuFdGa9WKnlnalznXx9/wSTF4fGtVIbkZsScMEu3
w03ycWcl7+QuYEj4JMnQiDpB2X8DhOOY5GuBYeBSZ44wRlCyQaUJGEa2XcOT2BB0m354WaGESPGw
FQytxGT1A4On7ne9x0xUtqOZaIa7X9zyQwpfhyHXrC0HhaBuxKfdbdM0hoqwahxkK8f8Inp9zggq
eRU3yOHRQdh8WyTj2P5Yl2ZssH6oLPACY5RA35YwgZP6Gh85KO/Xu/IF6lej74Oxqdq3Lp4x0QuJ
lclGi5PFL5WabmPrZEmT83faTGAmA6PdObKfUTy/dqrK8eVAsi9P8wfn7kg7CELdHsb0BScn1FNE
IeBqcpPnuc5sdLMySpqPX65EGh8HKAB4APUoiG7sisB5kR8pFVBg8BlqOlBOD/GRuZI/UMp/AIYR
BKj7XPfKPdaBLLVPsjvtDbELBdyCR/ouQGyZL4VrbGtdAI8nK/TdBxB74kS+TejPKYu7VuBfrism
quj6SIu05SB/DmkRYKbp9r35M9urhZxtV8waQI+y6FAU7y7uRbxD4lCscyXHo2yiLQigCQzQDvYd
fyBYIOIv7VZ7mdse7LaT7p9Fn/A0MO8BdxQ4C0SV/HSFtrdAMswTV3wfdZFkdkJXW1sYXgK8mUDX
aqKYWGwwJM7zeY7f3sIbaF065jJ3+e/iuvgHSW8lbl1GYR7su06UfcdthxYA2ZMliazjjhwPeu3E
PPkTT3R5MPn+wo9VY2lSK3aNb7EJmvScb5bOYOQvopMsq9VEcMOo73VTF6AwqocWrBagv9wttT+f
ZQtwkttq8lSm9CPP0OE2wBQcaYf9+Gx9Oyhy65pt9EGxVJXJofBOC1uamLbOZEGTLVi6pFCgPzd4
W3UhUk5XXLuzOnhw1VHETPTbO7rpgWbYDEXZs+Ij1u2nB36V7TSfoC2sQ4D2rRzcpxEzkVrJ/t/j
xeQUXISkluIQe8bFGi0z+bnvObeNn+s1VFXmLRfFtQyMne0Rt95PgkFVvQHiTfgSyKIpHCeyfNGF
M/8mzA6X8yzEDgOuCxUzVdXGZ4S9D+V5dPuCFdF+epsXPeOdXacnkA1I0XA3cJl8/uSMGrDcRQpw
Ue1eLf/f2rusp3NF36/5z9/PPxvsr9+Y35Ecod6meFPBGUKrYCW5KMIOatHchY0uDUg8WeBlfnh6
B2Rx2F9sb4nXeNy6snIGwI7xxL9YpG4lUB6bA/RHTQY0M5T9p/K2jI7yLWK6dbk/29z31FLIvQhV
Bjzq7Ant4dwmYf0xoG11sBiQErdUeakmmzuWwkedKhFruTeWc462n7mGgyUKHLvMlZjyOHOobLXA
uFHQ85r5R/WNLLFhK+A1gpwS4VtQ519/B1+7jTk6oq47Qy/hvkBfdpvZLmo06daPFdUVbk139KjH
Naa06B1dWZtZ0Ocoi8v7JqyTgw3Qqifm4P6EVxdSmFuvQ2hVB7wnkt7t0uODphvdMkMIZWbAzt9S
Bgk7yPwJoPUGS+BX+dz8YB5VveK3XFyp8AWHmdOjhL9iDS9QR0UbbI8mhh5ss3WeEH2OAt5gGAuS
1D/JFNO1SA8tPal5RXFOwOD1yuH46IftsWhCsfGC2VAkS4GbYDF6hcN2UF+/HpB9G7teHmkZg5P6
cnFWsagPBDMCfh52eaSY+5egTe0dxPtIR9qCzAnad3Q5/TR0MEgU4ZfRjNy6VG5NDl61S3HG7tfJ
fP3p1J90pqxjpyXkRDRwS2pbKX0col70ikChh+lZR+DgMH/V98FWwgzOnEOkj9zj+/o484tXgSex
lgbuTVne2wkmW5cw0dlZ2TAEkGnD/qmFbUs9JbvsezaPHPCp7fWxud+x6jpD5sL/bD5qN78kPo1J
9NbPjVIxGKjcY4JEgUSP7+N45M1Dw8c1iRzdVEVbr4tCe9yXIKM0CLXooQGeov7OjHB/vn08TWqc
mYPraz8XVrQ7A3Sp24kJDT81Srm1nKaS7j8AUTdJv/ig5Jxj+XxOWHfwLJki1SxnFMik7pYLGZYF
R5EvylQePe/xwRVfBWrB1ZPq/Z676XviVPL8Bufv8qfSBwLhnE2tmBockUL0kd6MphzPvE5hOiZj
92hR1kOSQ7mfcIC1KFk1zlDsS4yqGqGqxko470NlBSzddnUs1Nmi3+TdtXA6gcq5yn+6tdAZP1lF
GVSYbaxPx8Lr8ugWIG7BRU2MO8SP/44IzwW8+kVSw3LdVljPdQD5aFfvHucFr+TK/caaED57qbp/
Y0OD9I18tWPvS4bXyGwczC/PdNwiD9nqSbGIi8vAHkFdd6lsO8rsqd6kYR/bRWi5lsfn/iGgsIcZ
YoG+IxG14wDB690lOo0Ed++OqCu1tufR2fk7f5+AT99jme9jL35gx1MJ+IIgNTYIrEBnBB5Bvkii
HnXXpo8VYU4gBpIMX0zfsJ22+3U4HmayWrcSP5cGBWc9DHQqZxS6P9ejc2QbX2alWu4mf7qJcXxE
9FXCN0KoZ0SaTEGVAz4R9uEULGdfCqS83IQTI3zZfEOWjObD6xtfJ36vNOjP3mXbN6O7sHsqrNRR
/cAitAaL2we0+E0wPi1+odJdIvGYfQtByGmWBBPgjrSj2HnIMJ1LZIrjYf46hMmLoQYIMq/qBWFf
txyH1jgQd2FGnghGTmev2cLV1erW7BWyxBJRl3nWIx5CGyTgxkd929hmRRUzsHJh6vnJ+zN8n0kB
f4V3wEIRMCRo6n9DayPpd3d0KwVdBymeb4i4X5TerNaU24cl0pdb9szo2gBub7irhnOKgbb29NcP
89IhjklplsF7jUTT8ETAZTc7RCa8YBBWH1mTBE7vXPD0LNP5PAAvF017SQUHhO6OmM6CyzbViMxJ
9mKbbx1Zmr+CVtjLbOwrnMeoE8RjRfZjAqQf+0YRyZP2Y0GWOQhBBBGGUqUIDN8JPD/M7frOjbTV
6CK7NgJzHqmqTLfTzArZUC96nezW/hQ4hsjqqGws8F9QIOMd0+eQgAaQVibjST190fo+6sYH5pVC
gQduiuetB7g+q25QUhbXEnqHY7fvN39Jfymq3BIXYSq8q8L1ld55XfPi2wY8mShq6FtdV443MhOy
9y04KmQmhnpTgd/MwN4vXX7jlpUZKiXc/rWmztKesthdLd2ghOsNv0r/ndvR6wGpVY13heMwrl4G
/feFF59bnqOwAtDAOXErKDT3KPmk+s0L2g5mAH+CtesMRugV88ihTYHP2ZLf4YgnAJAMPQ48SzvM
EgvVaQLBU5LP+8aC48oS3q0ATPktkmMkFSzepgrKfuF3wwsQ1+SIr4/MYJ7qLL9L3parC3uR2ZEK
kMa9yO8OJy0Hf9rPYqVCAfBG2NywAoCt4iS6/q5PsHes7FnIFQRx+TsDQbI/DM7ZZyUZagz7DEHD
meFuV8gtWV/36sDa7GtxFOi8CjzaKHVloeBHIig52ABcQZd4Hbd+PdLZOibo4OtUE/0nAWUcUHQH
Xq1HNwEseIFdXL5Xc1WNhaQLiADOJRBG/Meb6yYQVshLMsNREI0/iVfWNgJ0P5jP5yJ9oV63HE9f
5dI8+nFKpn55QWdWEHBOxSscdob6alO+adEoBEXoNIH3J0JSCYWMEQDo+Km0zZugERqlgsFoBGDl
rJoWyQ4bMbvRO5qKInMmA1PaPH0Fp1irQsDpzk63Fj4EMUh9VhpS+mdjXzPbx1Ar5it3WmetXF4x
zkvPY7lFM2B/e/5XHw1OfkM4pLJ4GaGpegLdRVg1PIAOj2bT8CvOKujX2QuyUdS4+1x7WVpIRql6
zQMag3v6//LXNkT4//TdoYTYH/N6FO6nqiCpUq29nY/d059UfnQTIAX1iuFiNb6Jo1F0ZZa0QBcN
1p2PvdRVoV6ccWKxNHN0FI82ijO9tqIVnpEpVNHveNsKXHxD+lfAkACGH2OwLCt97CRWj6XgxW5v
iO5J9DCuS3Es/NWf3txtT8n+UZ34HuderLQShGcwOhz2NHTCai5Wey2FS5XeKvkdZLszf5WBstIi
rILSd+XuJEjxOF3n4H8HHHSsnElJj5wXFjaKsmbJbxF1s9CJKBxzFCy0iCOlVH4K7W9BAbccxU7E
RZxezj7Q+edscA1oJsekGqKUE8NYsEZxCTSgS+U3iobFAwnb7tBhKpeOoD6hRXim35bgcsmh73nh
2+E/lsXvojEu5O8VLeophZj4SbAkSUD+ZoTbGHo4BIMXEhAbYXgpdwPLpGflDiZHMMAFP24kAIHX
51Epq6ME1/XXqLd2WW66Wb9Z30Ewt1AsNAHPmeq/XQzoZdEytLbBmV/5f8HbbjlPKs/w1gGUN1kZ
P81t+hawRaln4qJX0e1NsGT3/yI8EfsSswKnNgkttP7IVsxE6sVbUlDI9oq06V7QxCSSHotUes0B
IOlKyrx/LYLi1lmNHdAbzRiVTX3QSLp/ZHVBLiht1QZXRScdge1xh8X/KhafmrsvGzJZO7OzYEXk
U9BsIZQODH4HaCr3Z4AKj6podBn+tM8guDUQjet/9HZmYf1suvMTOJiLMPvt6wslgZDoPuJMwcA+
ZbwRJTBgaXa6A7SEOCMlc9jR3EJ5vZhO4mrIXEuxlh8RJnb+hntBYHUs+YA1J16vSJMS+4TyVwQt
hF00b+mq8Xd5UXcnJGkzqFj+Zk8xBsJXVedw0lkK+n70Ta+PJLVJelSU0P2xfRyeUU4I1xaQrH9r
gN4gIzrYDMEOzMUNyAjBk2MHjnySodiRYvmznP1TvFfCFi6QcuAUHrnOoV/kHKFHUJBf9NSjRWYI
ySa98/2yrqz2ZCZdoPMKKvj2UdIEVZKVwmhrzcqDW4UiVHgT2bOpn7Q5Gcs/Ln512VP3JKbvLyCS
WhJo/pHDDkwI9kCYDMv6WQEAmoukffnYHvvMBSp59W3WIW1O+NexNPQhLQRy8s9J7LsunxZPMspJ
MidnghPWWGyKOV7+wrGzxbfC3M61rK6o/hu+bKLhaTYfwu6xdL+JPMvuRDcMRVEscaATgrR4cGOD
gNGKyvptg9ZRY/Ry+lN5gSPYt8hwJ37pDnNnt1FbhqK2/vKFqR51PYPwbdeE1pfrKJUL0e+9zQ1F
hT69NaicB3wfxyYmaApOj54JU9kMIvlj3O7vMsX/8SNnXfm0xflR1qtCrU4zhRjDlz4uCpm5In8x
+Fs9JzIXHEA+p0cPYXHmK5LpnwHCNbuzpqCl1N8+L/Ya6IJpw7XF+4rMTfysYy2lePaKB7mds3Xx
6ENpX8H7ozkccHfl4K+j4gvh5PJmspRkVgw0p69DzGWT/mgAKjl09fpfejix4GWP1D9qKEH1Zo2s
SiFeXmQQaN34EpU3UaUsI9NnT3PJx6ZcLYtkQ7m7rT2ffQszCpEdq4C05oQv3wArtEyJ5EsTiljj
zA+hQXNwEWiL2PXqEm5+NSYJQVMwQUKu8hN+Tm5CcRnbFerEpdihtqHw/07TeZ5qb1B3Pi5QAa2X
1ZxZ6GDhYMw3ccCu28Km1m5IhLYSmFd82F4JX9o5f1OW4zYnTbO6LnMEeF4erfCTYyA6zkp8nJ5z
/QrsSFNS+iPq4bfXZrxlFMOXS2VgKag7Ao5pQyYrYlJ1Uwd1JMwWpgosJiuXqhqDi1GWZkn+9Wve
iUw9bFZYTKyk3JIf4P5yaX909I3fpEz5gN4FfxBa1Hqid8VHEWWjccw7iZ7BicIv75c+wJfpLGGD
RJHL+EHL1+K5LqDgkw68ArMD8tcMWkDMckfMEQELB0ONSxpd2v4uTa1kg/OklyYzxE0/k58zyx0J
B9hBz4flDCT4LRl0BW94e2K40zPt1T1rvIFaPfPoq7fRcNMNacSZreYqivhIEZ6a1Exf3pfNOtON
+hHFdawwFx7/KYsqxozw79kewqYI4zVMng2cUUB2hC5LnOGe7gVR0Il7o2AF1OpD2lCx9RpSC96p
bvZ11oPNIIMKTRQp57IRNQS7w6hfze5T+7shKDHeSvK+u4GftKwjUzsqa5bS7eh5I808pzBMmbKg
E7VS+L7jAEwZWZ2wohzcPsEjUPB0KIK6O6FGsWvwbKR4n+tvwyiEztIvruFe4zD5IrFFXsOylM0K
bowEvs1HTJn0mQ+AMcaB3E9y5VCVDYShfQJGr3pT6OfAN2zopaHXV/hVCMQXaF4ih2EyLs3X9KP2
8tcsZD5el/RqXr81r52gcY8kc0PBhXR2++KRBLP69QigQeL3XOV+jZBg+eKR2IB9oRzIf3pCfUI3
M4CFOzzaFOnc3Ffx59Xa5NS7x9ev/gWlX84yKmZYH5YUqgmLVEGswetCVZCUL07nWcr7EN/GCzTq
AT2RYt+Ph1L+dQbG9buL0+sDWuFbgoX1+kCz5jWnPVf3NhVscipbWE7BIVb+0N1uFYfGyB58E9fN
qgi77MOxqEXq5dREwYuM3teigbTyR4akZUarTNNuvNCXcEeU9Yer81tEY3UXphdGhVOWcbadt0w2
go7h6vxM6KGL7pXEW1LPAyQq0sB7wL9rXEuDskVBvfJl7qZbnMubbw+aaxycX9Zaio1N276kGj86
yWa1Nwth4PMyAX/S1iouvB4nPGw9N10WG2sbJ2PByviMOIpMhq3X8NQ3fRXtszHx4qgKhPlKtk0A
24Mi3PDFDTiB1YbqQzySAmBhMNwxpw+4FmZzXCzMsTu0bThacnaHvvDZYp8Eu6PDoznpd+3AwKQ0
Ug1fgHputlpf7kofwtwcTWf7Gw8a0i8qYHRiqXZ+Nu9vwv7qX5xR/4bq0FZNsGxMcRSePLwU2dr7
Sxhto9IThes3IgAaSo9ewdrbZFZhR7u3oervmT267EgQGaamZy8j07xcPSAhFUIRS3i/xQl7JW2A
6d+qa/r2wKI12Ov5VEwjOvt6l58ggXJZegqaPCXJxjegT0k0oRbQy6Knhu0ugUejpXwlMrKvuaqi
aieftigTJclWJaiGzR++PRIv0uXEBVONZVtSmHci2Rp3StqP1Sq5TwPthAATF9LtorLktr+GFvQo
VHsywZBhGsD88RlgQa9vMpE2g4olacMSdHHZPfXvgEl72By9Wtdr2i7Xt1ybkQOSHjzDhMYclShu
gyWHibg/USBF98IRpAQQms30eYSG8DQpdsm1eqwTddfYeXLUz3C1bxWR9jLJtJOnA+GHVjc9Gedg
fM6HU2pDDUOFOi50paodBV1PUp5KiHCuzSz5HGzaUrE2zDaut/M6p01qLN7XnxY3+jrEWgZNij3z
ZRTYkZ5goJ6WgTLzLWkSM0MiKn+hNzp7ayZzCdfc27IpBzYKQbFD3CK+PPuxg34Q8+iO9wV1YXOq
kZYnqaFzVDAXShf8V0J7+Fm8dpMIXa/lKSgmC7IQ+hnLr5kFnq0cf5Q+kGflysH0SObcv2oRLHcj
ilhI8Fst1Uf46u5qwP3E8G74OXDw+4b6is9wjfqQR1uGVtw+EOidE+A99eW8kqN8kSXdZPUZCeRU
vkEGghW5hdPGRz9aRbFv7g/MFqmMXYifwR31eDflZZlI/oXfh8AEUMPhz05SdZIi6NZbQV8zOKfg
4mSXQle0nD8YtVMfNSPLDNKY7k+ovR19BpfRjVE3D4lbtiBEGkuYS7TZ4QGzlOyRKrQaftOGa5Ns
/aron89rSR6/zIKZa8QM8Wotr0TbEg3bVeZK0AsgnwZoRWwd/nWJtAEgFWyD2WvkpiDN5J04jfYk
+0vDDsfVAsf68eQ+FZNkTDHETXohd9OFhONskpU1Z2YLXxLCJOPc2qEGAvjzWNyLcKcl5/aIMf4n
QPB+X4v1Zq5AtGvZqjXwHlia25lqe1h7Nqrp/NfEGk/D1fso/xcnOBrY/SPEh2+efSmLKbTUPwGR
tydsCgoIsMlu8IaQ+ZlDiJ7YEqwLBE5cMKq2P2Tz0ZFUTqwP9dQzXl2uEavZQnJ9PKCgscYsG+Bw
3bHeXBh1AugFZKkigzt2rfut92YBm/o9QkCN0WiAbaIJrElVOv+k7O7NVj4kizgPV4PGC4KNZI6N
i3nK+FVNjVVswj5LDyJAFdbzGoPxTa+tFBKEpnNint5CcRaU3/Jok9fGPsCYCG5xQfWyLnCvQ65u
2LKjsndvlCXA5c+F6W0yC6MfRXbjS7wZvi6Dnr23Q9+wRnCXa/zNRVlF3ep2l54q3QyiB8SzRZwo
Bf0c6IIpahsC0aGeayD9vQ6OFX3bBd7LGMS2XFtuAoSsEdvi729nq2gOY6SWWEmxW0gf3HNEtG0Z
ZXayEXdXKo/3t9TwU/Rj6oYMDlzdVHWwHUahN0cT8oCj7f4lm4kc+o+h8iGlK4aSPI4+2yCY304d
nwB7h29TH1ELpvJEn+3Mo3ZVJlRImTzvLfwiQoYeBVGVdsm5N8Xg0AAvQK5EEv9jSd4uuXBNhvnf
GFUAtZA4L4X/flY6SQe9AynllFX3uOqebwUpD+MixAdDyiAlyhkEIp650IWh54E+QETocc3Sa5qi
RYRlx7A1JvYmWEWRQRuoLV/Ec/7OSlHXD3qD0vAppgwpV1U+GtQKJYRapZf/PxjSuMw8H4Ke1xyj
pZZiNVxVG0SoDgwOJWkbrzlDMCGH4jMqaOxsKnbNLkAFZxrPL9q2EKAn9rLoy8bNpP2d7j1Hz8Pj
/Plb0cPTCE22R2yIwgpBjeZZIeqqr9p58vp7SVKikq4efcn//PX94xaoDPbYFM+eVd+wBlBJPXVm
oVuHgUXC4sTSSRh8Yjj3kPG0SV8T9F4KKRZPol65kxGdrfFjMSGRUniORLfpCMdRYh8yRhiZZkR3
HAY72v4evkh1Ic1ubfkvZ3FFJ+9VbF08yXPVKMCnwsLah7dVvsC4KyGKvnNT+MdVgPMsksb7nhaP
byKofLyMAhzLuLM5hKdiGrHT1Lb150xLgikJMjivLeixx4hTIODTRnihr5QxT89XRt1GXbHoKsVd
xcUWm3i3p1b246USIKcEPpja720yE4QZKSi6UeeE0A8659onxUrKhnG1ZlSBmNYIQx5sno7ZB7Jy
kYQ96cJ2XNPFACDp50lyYUlMywYth5NSO2hr2/wa77c+o7n4NIIu/a6ACZTRZ2PdbAtLGUiCmRx3
25iElmOa3r3rZKXWfpPgVV1TtqgB5ZIa/Hkg4KVet2svdM/dHy91VKXOpupsyg0m9BeVSO0buebH
uoAbxMjIDG3sjRiVWJvAtX5XwYLnQC6jHjo+LPA8E4V+RZMeI6Qg6v8mOWsD/ktbBUJlyh4/JtFa
F/vdgcgeutH8rr551FF7Vo7G5754fPrVBGcqd7Lc5G0YxT4G6+Vf8C16twDxEnB6kmvki5oWqYKy
H3BalTBZcZpb/vHJJn5WmyV7w1EiITW+IK4qvFxnRfcIccDCuH9Y2jmaIn7tqP/tDk+nmUe4zWUa
VWI5apzvmcqxZgCxlVeaIOkSNBZHRqXXGijDZ8dBAraf5pIOvC8yQROgRy+D9tIee5pBAyJJ+LNK
Y+IqRTnSnQDnpCRmY1paC+7Ta2bDcTY+3mWPETTdl+tz3mFmAL8UvGLcG8RNcbYG+aHXddiFdpS4
YPQGEJxNdoA3USUGvJA9KGKnX7YapJsxEbF74S5maSL9kLpZ/ydWEH3EcMpk4CaQfGJTZTDedoMf
niRCqxIs6slQAmj3BOZy8gM+qF8YPmg60TnSOx+RjKP92Vg2AfETKfuQuTTWg0a3H28gA4VdKn5R
w9gR8IQt2tw+4/afTKflQujuDOmEjmBe/gEMe/MgqWi3mwjcxatk5hCVeEsIdmZ87kd+pEudrq63
rekIv7LkBKJTpjeCwMFolJXZj0q8z9O3ZPfJBp95dW7ahnXMeUuw3e/5sZTrGtE1GvI4Ydl/EfPi
Vlf6Hty3O/Qu8K3GkRLcgHeuLu/FMsIC4Uej/7NE7Uwkm1n4kg5I8Om+JnnT4T8TawLYuROXjUnq
9Q0djO0i/bsaOze+RhME1qG8tSlNu4zZyuA+cLHh53r9Jjd9oDPNW33Vy5EzzIGkS2vabgJoFNXl
0bgnRsXDkYmux3yYiqnd8M3oiOr6h3a/cccHOWeSlBKsaGU+tkzS395POrwYnB9xvlTghVNXZ65W
O8R49qlatkYJ+bldXKWR5s/TBMsaHWgMYlWMJjC+EsWfe/PHG1m8Y4+fC7l248RTNDXD4bDTZcCG
/+EUYNBKHhWGEYCpZKCtwV1zP5fCArFquCkk7WCC21xIzbH2FRQECHApPXYCkOSslYwL8UDxUXRI
Q1YP2xiB5eKx4Twh4je3gImoFUJv4wnO4uXp5lxbtsOF+8/kETgh0S8ICsOal2wuSSRBLhSaUZx5
Vkr7MkAGaIdMtgWcUh3fp4g8EtC/ZzGdORvtSdCNOQirH2BSd023Ku7bF98qtFJm2ND+SXUNWObH
H3mKxhh21XBtIyyFXs6WJMpW9A9knuHJ0VRtk/0gR4DhG2h8IqyGXfwWYw6/WpNlpysa0LlqPGJG
R0afuhi0OhVaNDcW4cbJjNwDbSauUizIh8/9CO5O9LdYbbR/zqIUz2p1isQuOhHVlujShIRzs3n/
Oj+Hp1ekMq4eRtpRbLpIGRpLhFqw0BeVxhUUF0sOciG5UNP/shr7dHcyeUduG/IAcpvd3s3A3m4e
oKYAzJb4XU1xIZakWsZnBDjH+zdfubSfzojYlBcuygFIg5j+2slI4soj/4zVB5e7gEyNOqrkO5VU
KlZgTtvWu/eAuPlYsbdBVa3TN0hhBfKbUEIWYIOgi9FdSsdNE8/YzunT5l5J7n1d1pGXCOKTQHxs
lQ+2+EBlqG5dKBXIIiPSZcOK2KHIScbeoctuP7Xv4ITNnXOwOyngtC/iFl0I+y74h5ds/zBX+en2
+rQI60aWLxx6zUOdKgjlL8GS2AyMWM75gedZloC8We35OJYJAg5NoIdcDOYL3hG9ZMthxyzAVCg3
4tsoParVXp4xczhb8uNiHDoyB830Q/Rs+6DDhX89T90+MAjVDR0+cRkmOfSc4+PH/wDru3S+iN7R
PN9JZCT/NzyD38LO94uqOFDww09N7CR0h+ewUM6/nIgSIgrF2MnBdv0u93s6IXwbMNUPoEumGW0C
9xCSQ/Kyl3LkBH7o/nAhJ8t+Cz6j6sQ84g7KALf6bJZfWrnWBA/6vR991H7Uu61oTz6MPr8CQqT9
isaOJDTPpwx7decb4BgU+1L2oIipaRsTkpuk7JYuHNHg6TqCSTcpiWA2mdLhhHe+g+Ll9FFHlbtS
JOcOcqaxqpSNnBrhcvz1GcwKlXJXAl4GAWvzod6U0NqQvC2vcPA3m+OSoUK7YTH3J+GrCJW+FLBm
wfsWbUxIcdsydbkUm+nyidx/BMYBT+bLETT9ZlIS8rvXUEvw+3suGr5u+kBAmAUEMuGqqafwz3Or
MA0lWrcEOjHajVhTjxsrS8wP0h0I4csP0WDW/x+0r77jUg2MNoeasiAl0uNVV3xsPNz9HtxEsq2V
asPinFYLX1f5SDbDwnQi4JRJm2+b7kMIgT+YcOUNS/ikUXzTiV3juhbIQ7Oo6hJ7sZx/U3WxSbUc
bFTjvhy8Slph8CSzAb4VwQfbQfDqNz2nC85SRgfcoh2+qavO4K3V9THWU93GGYtXi6sOzBgkf89M
K0lpeORzmZpyLz3wM7/aUVsp/HYaVSs2BBAK70E3vtg8/Y0IWxdJEFs5uw1UD8opwKbKkDA7DPUb
ugIo8m4HYq33Q52JSePonUSODrz/d7C6MYFdOxvHSNoFJTcfWkGmQwTwB55aPJWP8zUc6S85PvP8
TSjxvJeff1s5oRMrrScqx/VRx6n/B4h5+zjOUXsnLJxi9OjNkxdDncSlMmbu4HUfE1vM0fA24xeZ
Un+qqVXlN6yHRlEfjR/BkLzfVeEU/qT4/F6byCQAl+mXbbjKJnddpauzlfev2O3dgS8t7oRWBS64
5hlmxrFhSbI+CPBQm6ajO71V7+WzwMlgr8nHuc3v7JkmReXgWyzCxIQCIsD0HDqyGFCF41yoc4GQ
BSF+3nxy+0CNuihbPO82DwDUUDm8OR4jDNLZebZIblDTwMMR+w27IXnJzi01pdsfkz7ruXe7xGdb
CCLBvP/nrlVvURnmhnJfaSGU5Wo5RiGH0G+M3swZAnp1VfgCSa3U6MlvAFsk1EGEr3UJJpceqUAw
WhVBgfFl7qOOx50CTLsVPtVoGvdhSbYseAxJzFV40vSrIs1OG6jlVoMwrnlDPGVnDw0xF4spl6Jp
E5rVgPvLmXYOA8sAtg5ZBwhPRpbl/vhrK5jd+RF1QUvK/ns0GicQ2YHvcz2jTLgRkqIwMXkN8C40
wOSEFKYPXOX68+dhgbJLypKGmga/X2S1GjwqH8Hxvyx0LyOzLc8HFXblPD5n/BnFQEJ27Epfhjbr
wi/3mnN8ja2rBWOTcB3xB/phnpGaeVzR0+102bchHbzmKErG614nWvL6P0MqPPqZ2f+oa9Q27L+e
Wy1/9s75m0OBw+Cjag6yNvRlsnwA2vjN5So4ybtN6nZGB8dI8BQVkoAJHKIsTYv46g9vjPL8ywD/
4KAPcZv0F7baFeUMD6pKL84xhAZngcLc72tq+rOq8EsOcdlg3plOtxdmIbeTCrEHz7GBNDlQLxMQ
iQk8Xexe8lFqbK7+9i6yMKlCus+stKo48NhGaqZ/aAwdq9I2dK8zHRXMIhRPxXeYdPEY1hFD3tM9
Y5pN3HlTjL/cs6j0h2L43midPgrjrS6PO5yKivT6R78UK+94OyLNnbvpYKWAIMHVbAx0HW7Lt6SP
e3o2dAGD0k/XO/c5/fNkVku7MS/7dmnfnp/ROWCqlTf2ftmJILTb5gDF/3q+pPu/kh/T2KGHDJ2D
nw7RA0lDj26vqiiUIrv46K0IHEmx793mp6FiFruBVtsGAWRXUXEy1Yx/GTVCRZBpvF8htnN+dDjm
TxYfnBPGwtV60BwR20Rr/Sv3jHu1xkVDgBZiaSU4KQZV3mbGfrFrhVwBWm34lcEnV9ZiOe+tUjA8
3T5u1kol3KVffugHtSeE3hkxQXIAc0WVXYUub8egMJRroCrQ7+7vKdmzBpr5Pmi5yumGZYLNXyyR
s45J+Sz6sJmBGyzxHCvwd+KUlzAuEn6a180QClgR6+rwYhQNnSQ3kcy/znQtPvmGb8z9t8xooh/9
+0bhDKGjt0heG9u3BmyKc9Uw4Bp5bmlcLMBB+dSzYGUvmMiQmixp25WA2AsZGIA9/67ch8WF4MM2
2R8O8igzb7X0yYXieAOwuI92Hprx0BK3JSONo5Trj1OaywBHVocSirEo/5nK/dw2KXyj8/AShYjd
V9AhSP0ia5QyvmZDGVLGpnT/KkH6AsuNBjdITdCo6g5DGaOiMGcIN2TAh2RD6kahVKu2uSwfFbCj
8ICRBzZq0dGDelPt8pMGX2IU8LzlS66RV1lGhs4Wb5o8WAYYEVUwMjf/+tHVp6EYRMjAyfOjGjzI
vkni5VIRNGLcSKl0PWF4E1scJs7ZzFKXPLdlsiwu4bkmafxjhSXc5chk2b+KOxQto97wsaqrgctq
AM8ApPl/coJ3kOwaPiUpGpHEDRXe7lFEYjIXjZc60LNL1oj1nyhANRytQrH3JXFA+byIq+e6ADqt
Eh6D0Ka++vIUUmU2O4FaxBqN7ub9h6sokD8az7WMTBcOumO9MwPadCT5vCmpeT4pXnySkUMcZ3KY
OKWWifS0DOfIQmi6ew6RWFL1i9mOERYZBfsSuDyM/84SmtnFlf0lZb3qiobHSFAL6Q4vz2JSelD5
GmIek/AzSC0kG6wb1XOc4lOJ6HW9ykN5zrb8DBv9PsWiNobmXOwYtXoaDSuKa9rLATT5Rp1lOlzt
xXIZZzlcon1/F2PERkhZAyyhsktvdXO9f+f1Tv8EYRd4CJGaXm7acioPrUJSwCHY8EXcK1a4hG58
VSZZfqQyh0NPOu1MPI/KvYOyP72NUbU72q/5TqSG019pLivpTNOrn23rZcYJ93YlejeOnLjPTgdI
ArpFTkNvgrl4G3pLvqrES0PTBQYPB3Cqoon0hTf9kyvPtWGUypNMTjsYMpxy94HjnpQwiQiyOF82
G3z7//Q6HDboWExuROXdYWKNLaJuDqS0KiHBxULqVNCE2IRHkNmU2sfa5dpfLoMFWglccOqb4u7X
w/qRQEYe4me+objn6pUiiPB707QzIH/jOMZeFD/Ydo5RK6kqdTTM4TG8xYUtWHY7w1hgrBwCmyi7
fopuqcW8LyBbIGz7wihgpmaeXuh1EMpwTl9Pi2sw4AJ1CJiHxUd76T+thhhQDIgiwWSw47cqNuF3
VW/73z08V4C0V7l9gGbo8Js7KEMS+Zc7L4Zqgol6ockLEF6ZxYfUDY9WI0t+G9zaUd4p0xU/py8j
jNL34wSBfU/7ViIrHLh7uf9fWa0V5A0H0ljGdknFwxFIEnLvpCyZFNLZ7CBVjk6TXHTz9JMBv171
PqjV8u42PKPRbTbp9UOdBjAql9mZwPWmUAEBEJYoDvUdHdD0ig0GK5X5jOstZLLKMYOCg0U3y+fz
OLMConASlA5EveGnS0kVdHOzjN7qIpB1QRvcujoEYjgkkNppqaHxLQcNU6WCBiNscXt/rlQnKOcE
P0PqweDXAXE8VEwD4LgnCtWen6h809CjMQ0jhzqshciwjUQQj9qEmW3tVW0skqA9OfH/h3a6k1mm
M4c05No/BRoDejsdzJo+eBlTfO1bQsvtecgp8sGI0FZstb1LmMcwkasuLTFusKSySqjM36W5dBX8
X8Wgft7axRsXnlJ7yng9cAvtFnfOKr9V0Dg837DodNsOp9WnASFAWxZVAMZwbKkFIw4W2D9pu57n
fCh/nkmFlwUHzBuNb9AqaLb3SRzOHfuInnWcbZr9E9EvaC9YadZOTvw0vsujOttICy7YrMMINhht
MOFdVQOrpn/Jm1nXxinwDmlYP7I1Xm0NZxfPHyc/2Bw/iq7JL8oW9fU29XdOFCBv5HR6Q1JDD7Bn
WOHg5mhbURbUM7CotckOoqICm+ttKgBno6Ii4wiLeuURFGopB5NRm8UGdda2kwE+TumBP0Nx1tdN
GuoGVLCxPSW2tFxX6ZPS18l0CnMs89ltj7SJVKx8kn8yTv5GQP8gvqH0vI0+1n1R5A93fGW29FYA
OWn1SuoJD2xwwHBuvSPptwvMzFgvUvT1lESUVGmz/RgkvTCL3G6w4UcWDT4MlMy0pOWDKl2KOTuv
yFQmmx90VRFFuC9UjT1WN7ReNKKgIpgD8cTglcQ9doD2zyBIHWsdHUg/98fnZvZ2+8e9hSpVJ6lz
TD2tAFHLgMWQlXIbhwseOiPM3KDmzTICrJu1V7LFDXgLNCmE3Y/fmRoumC+27RTjMv2nDny6I5bi
YE6ly30yKtwsFqmXvnmCt5E/kgqDW64lSk4rIz5MkWQ5L2bNmNUXIkvLp7Ku+aLK1qSmLmN8Pgyl
GlBYLem7WrqdaP4VO0Eo0SxmJHBlmzlnqZMsigK9sZIWcBT1KzTHHcNbOVwxAb6sPIbOBTClGmO+
QucH8enldJHrM7Ihcg7GXf0PfFdwELkX9CinzWLf7J/lQJ5z0mZKcc0fCVJvmYidSNSQwXIydW0M
S9tSZ49RN6Byzdx4HwZPgjv62HZ6pKdroMz263n9OAVcfOZlhfqk5NCqcEPcOnk1Yuoyn6Q3ig7E
jljRqqcxwSqrKqijA/17Fj89GaqbP8QPKJVrRWQces8lRmc5d8Dj3f+Q4haPZg+eiNLaC50v9tao
V7E4hEXjiX9OU+8/LLAiiC7ojCzNzHZ6Uc/830d7RQkezSmOPismCLq5QjI/KUqdxmERz3XWCEUD
GgxslDNT80cVRZMGxdz/ZvDmusZoZghaGsCSz0M7bc8n7OwfB04kbbiMpX7zCDg8v6XXuR7EswdN
IbzmiR70kaFGdOIGtrGc70AWsf3HN0dVLb6fdnj2Xua1imSzGksQMZY0No8wH2lvzMpGbiowLX0l
BheVRH2m3GbuZrsgoMTJ3oWD2zG9bfJlWvj8AChK8pqpGl2B1TcYJiDUL0oxMmGkEHq0vDT4jqht
a3v2yXm8tc9UatrAUvSZNdcciDI782GWTkhmar2ND/TpY9MDECH4bg7h3vN3/igOEYpo2a5kO4A/
joWq+Z97e2c5UXEqcDFAwGgRGtzO+cB72R/838fl8IQHlb/KC8BmxCAv0wZzqBQaW7K+0WzUcy69
oNF+CmJt8Klp670v5Gk+qNgHnIJ3aXNay0GZ0TA47OhdbPHX7OD8gtg6nPxIQWG5r3WcGo5EAznH
b1siz6e2t9YJf5+L+euks8WtKVBOk7VcV/ZBb9/+yKGFayFZzjJ81szAdeqtYF4LJ4IynCxSXn28
VKk6m5CTsWSD8RWNOtCbs5jveqQ8uTv9lCoWt2gC//DwPI8CKt9WNjHGSqOluZFM3iv9H5z72ku4
QeVyixUFvFEoWUiR8wnHmekcRl4GmE2SwxFnk7QUAwk/Atl9vfsxqudcNyRlJLtmYgOEjaLfSQdG
RwUXRTiSGXCOWMmMLetcjBOTExa9kfOnrQ7mlYfrO2Yw/5KhUDGiLo7Cgktn7PVQQ94pIok4otwo
9nSDcq2yxt798Wgv1z/5qsLonj8opEM5cDTHvJI26q36iCN4oVW4MJcrBuqMuIdDjPSqlYs5Fg+A
0qhgxVc+L/zyhBx1j8dhRwyp9DW5bcM+DBatSB2yrgLt850zIQ4ngJ8mxTB85G+qjTs1e/DtNkdm
TxEdFNfZnbk6cQg/sSqJOVD1J6xLyfe1dgZUAb1PvYN3X52cHf0lrFmdwE4lAu7Ys4m54sl4w5Nf
6arLyBMU3GkbOHl8sOA8Evt51Ma5SPZE2+vk8fZXizGazVlEzqI/GXHuYKacaquUHY6wudEO1eaF
9gjXISZtKScHLqev16cXUVG57ufv1br4TVPcgZOPEYSc6XFQO9SRXbsSgYFZ6nOrH9mHR+6X4Zrt
wNNtN7rXZs1INB17fYHdkacoOnFZbxvHBIME5GYXGC9epsZQ6LtqJurYxKRaMvdCDCB/VyoaDpPh
CscjYyb5XYm0TMRikYLqu75OxdYYGiGXCF1WEYEeN/E4+c7PVCLzEWbfMF6oaBUxX/sM82tJPJoq
qQnyzWaMz7V6kAvkn1KPNj2+xMNs69QGrtSC4b9bINjjfW56lDdrkXRUPQ6hy1sNoJ28/zLbOcGU
r98lNibBCLvw48892DIJYlmD/co0gUwIWFBQaTnS/RBW5Q2qjNsBS4jXH+Fr476QcRYob30SFBHK
g1lu9QKC5tLRisNKj+inklq3DsNa1SMWMImW0q4gifmeYGr6le81wK9IUZ+txQA9XtfEwrbthyya
vT+e2358KKu8waeg/XHcr6Qx+xWR5MOZBVvb9z+PrY246H2LMI7mC+hWARY58CI1oika7aGyFRck
FDow0yE+w/kn7BrW8Jw2ZdR7pRSu+SiYnk/WldPdSPHwzeAhYS5xEoReFOMWpcyn6LkPtoheaxHU
s8KR67083BageJYAzfYnbUHl5vrIKUirjfEG98KtcJlAkpYwECP+EZLvmoSgTR6QebpZgwEjJ7C0
2YJv1//oe7QDCiBLImccdvTSx9AIp2AD5RnASd3J11AE6NG7lJZwnsqj8hd8b3fj0MixsHqZDw6b
NuXn5Ny2uwx8+QjfHsg7vDBDqEQQ4rFWG6CAsG8oHNcF/EtgDV10mHL1IrnOufQ3mAFBhZviRiRL
E7DEu0j09P2KSTNpptna1PFIH8h5YYVxSYVethneqWc2kmp+Q1cICav40p1FjJRJyuLAuNMC3Lsg
JdJ7XRo3g/DkD4LolOnTPOZqMS+SB2SpurC69sUgJyM6t87oQd57mfSlPEIbOq6o22etLg1maQ7C
U1nMnkHqlz4GJFYkBt/rzCXKjPcX5QRfzeEal6tg0t+5JhtiiRmFFk9ku70Q0/jShLEJklHx+7ht
AvHzxZLNWkHIEnXxfsBKuIRAPjVDcoD3NiBhOIeq08XKUa/b4Mewr3vah7JzP6AuOoCGsXVCV+ok
xcCXGAKqJto8KsxTK19oZvEmF/7YV8bOY0XC2mBS40MyVTxkMLWwJBExbFqFmvWjhEfYBEgVRwmd
Nn43cLxbLgl/quhGsfxIIxMyQfa5UQJRwe3Z/UHbCfZIMECwI5HT4qsl6eCJz2MWnGOJM4AIbbOu
cYDaH12TriExi+svyaiBHUpVVNBSwZn6sEGskvgDlrWESQl2gKLQ2EHdT8rfEE/PcaBnlFZNOn7G
HvOAh9MeOCC6wdXlSk/t5QmnBPGAk76VfN+ttSs4b0Ht4Tq1EEmg4yP27z+FBRM99tr8kJn6d8UB
qXChyNUfEwvF1vxrgf3smxVJQ2N2ctePwsa6ml1hL7ku0AcbqF+yNKJK+VvNCh/tfuLhTrkwQ2a9
HFpLUW/9tEhgiX0sEwtaWoW+vzmvI4qOwQykVtWNx+UwoAukxj2NAyx9OGqhSyT6IZSOux9vszBv
0JUyiqngOkn1GaVgkHJ2YU/ImfGy3ICvsVcefHocHU2nXKEyr/RiD19RUcxPemZwTRf5kwfxum/c
HV0LgQ8ReEAFhI7YzciDqgVEgwQkTV7ZfnHrCMQ5GVMqITBIZlcb78uFSq1uZgOfAKHaZT1DbhXx
kEy5QqBfKMG2EpgEtc69jE2/HsRKrNE4oJFRsx9ENxO4V0p65mKHcMSm1kIJKu/12sTEglE/VP1Q
eSz7jLY2UAsskIyxHk8vu24OE7yJH86XCQtp+jCxGsRhcdaH9H9LcLPTew6u47DwS3gPMyUNWURY
OG65frMPkBYn8qjrrl6FjvBa4XA47TZUBNfez7X5gpnQ3ia509p/+vTzBfCPGDL8wun/H4BZhpvY
Vj2guyvbiQkZMqLTeHfUEsVm4qAM3RHV374sLeNI+5j/v0Ybk9iHnAXKDHOR6nQXToyENU7kIR5d
tPMttFADloGI9QFLcobfbMOKyoy+wkyFkKnP3blg6dLBivHRlFkqKIQj3t4kZG4d6kpLCnAYc3OG
8ibqd93vhwh/MPgQbPTsSi0wpQCSkA+i70lcV6TN0f2asBiAo/sbqPh+eK8kQFpbVrOv7LNtwufS
l0LgNhJtzDhHDGyOMTHN1JF6zEDNPI1FFZPONieihnssU/BQao3zEMbxlIy6LeA95Ndt2NKSYC89
JZLM/jjCORhRmRVlUs6lYz7W6BFyZ2jV6tCuh4wxVqi1FbBfwKeZSlF7yiCgh93dKhASWeYhEjrs
6wQAt2mTclss6VaYDd8gczQIk05Xuw+ATGW1pvqhlINUrstnvVCRaBRg24wryii/58U0MEYioAzs
75eYBosLdZULx27aIbjSJY1JWcmppQO9ZwNOsqjh7Sq7kY1mTmDgtHn4OtsN7W3mlfrtZ0m/aGqs
mU89CQ74fnPyVUEJNDtqzU3mEx5y9thSHZghh7zVLBczExPB/yu/fjAn38itztHZz3/ruvtWrusV
FwA5vqCfT/eYck/LODbfOvr8v8bYwHlkiRAoFzcOV6QgVB335yz/IDvI+V0WEoN3Yc5RquKV+gfE
aG4byAlMzcbALztxj6R5QDRBeR9yJnXd3glUZ8QC6hE9K0BIMBQLTm2qWjavxvVcqKkHGRHHUiH5
+lNaBrIcjXAKO5rItvS/nWtS0+XkXOBxSw60b9gV1IpI6qNvWi3PTBw4KmwHEQaFJv/YPugQO7I5
QSWjgt7BAFnewqgHBSLdrkTC0WQ+ol07C5JwBjiQEP6RPW5otaIHKQQbiCTIUGIu7qx72bd9bXqn
DNEdl28/iLhBzs4LwAWXzgfJ3WDi7FZlFcSXOcXqDF2abcLt4Jg1S7dwtb4tfROqE62NsQKWds5S
+ClckS8rczftciTf2E7DiBbeMboq5iUQtgGiAe37FyqjrIEbDl3iwH79FKdRZS2lQgGPn2Zfg9HI
aM1hIaVfP8j2o2fsYWWEZmXnThxP4Kb63semUVYbkQKkX8nUmNZGOx1RUV7vCyHjQHPs7mTdktu+
ukyp++CdpikDYmSX+DJNFNypP6p0JSvPbPs148WCxpHsHW+uIXQBpBILJOhwe73yeqwDdySMHpz9
hYXj8ngSWYvWpAG9YoTX0n7CPfQmfEI42ykNeNvcfNLIbsUrwzzGL3hCFuGXel5vKi+dpkKnDBsK
vQtdhTBHwYAOXro/eVUS19h74w+QKR9mKwxJeOlgwotRSKZKmxV7c5rL5NN7s9EtB9NkM+7enS4Y
Z+QKOuAf7qLlSH9DI0E5XBiBfUWKznvzGu/Mkm6SP95SuhY7kqCdj1UOo8dJInfZLV3jtmU7TUH3
j5SUB8+egDRFtEMsAgU+5EuvFttCEcB4RMV8XjqnvkDAUNxWh1loP0iU8pfNKydM/u+h9WPWC3mX
SWzZ5VvyjO/TBy/2EjPwxJ1wspOntPmjYWhtYQTy88NX1lnTp9/YsOGnKfXNJc+rf4OAoaJVxhiQ
RsN3UmXqocMOeDkVomzkRncm7k3+s9fD3486aJlSR0gyJC1AAHkntCsssLxojzGp8rFxKJdYrpQw
S0UhEq2BqWwXno0bJuD8VUBFZh0rhn8UAB/f6p3g6s+2mVg121QyLezhmKMtpKbrYGJcJfsfyOEq
KD193MnJWPycKETi10i3pdDkn2f2LaYB8JckD1xK9+rqwycFFzeJPadD7s2RB9d2iR4NepNPpeN0
GFbsotBGLBLk4dovbvEZ0URsZAkRAiKCQu9Rh0yuh8GyVyl7WlSVjT3X3qpENWJNWyvOOtZyjl6J
ruIyZbu3ZDMTqUUAYhoYSNzJ6ui/JkGdV8flaQ5YK/ILtnMpO/eBzKRIs/WdUY1fDsoUpdVbNOPw
OnrB95Y3TXx4+FNu1Mo2rV2bah8Vd0ye33KT3hEj5hxs0rEoPRTB9sjobdWbT8sfOW7N63k4TFvY
ajg2BnlNb4AotYi+pc5+M+leiaVHJUS0+V52GNRPnJdo+q67LjGSztUc4ALZLLgYWEegzJuMifKe
AzKM1waOixQY9KDdZp01wC43yl4bj2AzQjgb04W3ohyzGlv9A1cqlb4Q6bVcg3fh8sa4ePN9a3NF
rCC0fIy3/3X/IW1476HWsN49a1YyROeoov3Ofx//+LkO5FfHci5MoBiEDouekVdqCtojsfZn+gG3
IKmrvnlj3YdPi1g+zCKNYmfMf3UFOqqIBkMQRzsEmIf4AvIQgYi192FI+hDt7s3HnkmwagZfyAwd
ux1dNnOyzzNd/R4dsJj49796bkf3dVJKPYDHNAcnIxTOQMPQr8F42xaDCxrljfS+VwTBOCdYDl8B
eCdcOyRApblmPzEphM0OjKjGOth5/Qw6w9GzcdiosBwtV6mptsfpjznEYFG45V42U+V4db6ICc+7
9n73ZADYIMkeQ94Qlo4KqeWk8dBsmNPowra7FX2aBt1mXfrDzmSjA8oDMR1V2MtFXlbI5FYQiXT+
4J4PbZNhFEUsPGrBpCBJBiqSrpOZ69DFrog39MtECCg8GFXxdF3/YWmWYs/dzduKq4+RmSyB2Um+
Bca2PtuKGqp7EVU4nwePeYR0yNtNiuPZLO9KSevWoKKgccXBjIjG5L2LbT5FmDcADR90/gtPR+PJ
DVTkKIzp0cEctBD4ej73/BLENk77ZK7FtClzqqFR4m6ML/isD5k2rtIPQ5AjFPHKRw2JMxoxQXy3
inU+GXAjmzP39c3tqH8tNRhKjxmt4LE+fMceEtKgLrMHX3oml7XuKxuxFZ0TBN29eBsnlySfV1oM
Q1ddLogTUml/ETlDb86cs0FvCqA3N3mIPFNc3sZ9WaUuuxYvKasPqiEQ2K2HWz6Xs8fOsaRiiLxy
PHz0Y78jw5ohhmAcmutSx7aSIDICmmGkoea5482o/cfOak5Uh+kMNaZ4AapxXK6HAHozUKoWD2qt
daZKj/CdZOc++DxPE5000ux+mBNburiXyk4xAEDXE4C/MMGZq/esBsBGO83P4A/t3Pjy8a0EM75D
jgrKyVlTpydYYXlNOK2F11F5vbcEsCE8AndxIE//fuZB+Ff8WiJsn2IiWlaByoGxS8czbivped/I
xUMOVwposbldTkWy5JyUKxOatD28Zm+0bMdxqqAz6SfMgLMyjwF7fN3kyJjgMsudSQpRmYO/3mOy
QwYX9XwIRHHCC4M7hhVFWFUTPLc9pkTK3T5sR6RW15fQEctFkZEQQaaCfO+GPnssDH/hmDCQWGUy
ZsrHX2hFa1ZA/KEvNTDkmE1YBL48guDcl6hOeql6rmaY27XCVTcQ8g+KFpMGqbNzYO1eo5DCev8/
ePjVrTnh1YT4ji6xrFTVxV/glMOEOsD2pvjjDshBCf9TEU98GULrOG4YU5bvK71O9rpsYGyJtKPx
bCUozKbVIovFCApK0bZ2Im94TQGxOA7zMILIhYPwGUZiI/REKdFrlNEbzvJvZoAQFKLcB3EoFN53
UNIGTD8Yn3fret5acUnd1MSLhvwTcdfOwS4a8J4qWPo7SZajwk17FHJT7bO/OVgqJDX8fK3T0MQh
drkZfGWzJpRe2J36wMfO1Yo1l2v1y684yxuKGgLdvil4X8okUdoKxqeam9W1q8Wzgiv9aKhzQeYk
zHxofNfqwNntTQdbJkvDvEV8etnEHCur4AYnEQU3zfbhZ0o4eZWU3SUou4pHmIIRZ0pxj56jTl3a
aBdVe9ToPAlzW15HWxCXZUdBL1jByJxj7+aQZufQGdja079ooVgB2iEa2rg5vQVrilXjWBQk4HZS
ZPS5Fho7fC9BQEVt0ejfhs6PLTx4bmVjzYTYMtTD5x5jeECT2rbWJcKXakfd6VHLCVYp412uv2Yx
j14zGSsstboW+LOm9ubolt/zrrsQTTGahK8ZajhTc95lA8Rd6N1yxg5huCuqii3dLhuQlzU/3yv7
39ndqfcET3pH+P659MAhXpX9Hf6m9t2vsf6wxMIhmK4VBw/5nOfhlw9/zH/6Fhy+/Y5FsC58AU57
GFA4/eLqOEtZdYgjJ5YneMuAkOl59mxRrC/xIczjlHWK2DXGzbK8HLctlFEG1FQCTxnyefjjguub
LuOFI30wwGIhm4dLJlSGQ+Yx9FvlNqNm41tLbLK6/7+7BdTdCnKJ56mMTvIvIt+WS/Llv76vs9Hn
y59q1vivqPvlRhdKHpXRs/9TOnoHZfalAqpSVlLbLEFaVbTaOFJidr/KlbaGGRuzxoeR+4GUvLer
3p4rgA1UJVKOVKLJ98V2IqSXopRGP73BKk4SDaAmJg+rqA99GY3+7X8vQBlOQew1bF8GitLBtCiK
3ZNGVwBbzdsdBEPHKQ3kYGpVmycsz9UQ68eh2bSWH2xgImoqd0SK57FeXLBqENrl27BEhH510C4l
1kY1caBO69KeKZF0qqkHf4tJp0nIGFHMeSNa2NotL1gMTW3ck7EG0dTAR19RLlAlc/btBSsDezCY
RYbiJyC4HGk9bP2U34RFPChp8UIZrgCEYkbP2BQA1qEhIEMv1pE10irnyN9aMx7GZCLz2kmkCHeW
Iyj295uRmUpxHbys4XCR4wrjItbfmIUMXmv8ak6tFEhn7bzr+g0msLx7Op4S99nY+952iLfyd3zp
sU3WcrhzR6pD9uk5CMVWSlU4sRJOrSLTaE0WS1Nw0UxqEMfTbDIZaFPStKsyp9070AcSSpL9Og+e
C16LoPuTFueH9J8OPch9XE44qdQlJsZbdOiZ58T7Hup+zxnFTZY+vKXonBY6A2OwqiniIBzDi/tz
h1D54ApyX82s7/rGucgA+qUbg1XQz4v8aNro6kRfsxym4Ffw9TeQKuVcEF2GSTtOnnNLvcWHTDBQ
W+K2EVooJFb7HEDTL3yaGlcBCKt3LOhZPkRGMWf0y8RU6xpmfAgIcWMCinLGT802WBTe/nluGnLh
gjiU4p5wbxVylLxxc0zTnol7ReIHs3S5xUlOvolAzYhrhwrGGbh/wTCVvlvHNPyUEDvEBUUtSc6Q
WubwiOpazxCj76wOOgVsr6b3nCsiUHnT66vCiCQMK8qSaDOokeQAh4on+lU5eaFaeKMDjZPboXZ5
8z+VI3O0Itn4tG0048tnygX7l6pstxxStxhV4oCkaeUbsb7qsV8/AmRW9Alzkw57ienW1tCBeXC+
rgQ03VkSgJT6uffLr1ROA1W3FOU3nS23+hXU2zM+LUpukrD0e8jAVYE1h4nkegnjeugFqueiaE3T
3LoUQIXJEXHi0ggqWqE8/x387+Y94hlLAH9c9g/cPG+kUE5mlv1RPzjDph+SWY/cEaw3ybp1MLbp
+torTY06h0vPW3HQju0TzpN/zQXftFjT8lR8aLfhbt2irbTwrtX1ZBjTtPcMfmIPTZ6TruRBGHEv
CvGkxSUkHUiYWMAjyO4tNpBMm7HQfOcVP5Exv5gV7M0zEK15vQPH1zlCgfg+bZ2PGVUmxoD8BPVV
aKBf6la15GM2Vss+qt2K1xMMOiaOA92d5zZPQN5gbaHcptmQEXHPcpAhU2fvtSgY3Tqm7LfYYxMh
tKKsxLpIpbvC7IZ/hw/+BcqD6LgydyFUvcVXz4mz55qteDgby9XIK0S5FN31sZNrh2VK58H6BPSg
vna+sg5vt7s7/HqHjK3ykodN+/z3edxVoWhWfoF6H5BplTLcBskxhh6QJ/glkX21Jefwb23WICZ/
vb0n29CIo8y2ohRrQpW25s/qgUbFWGDuikbsYDGgRl9n5f/IUlYJavO577p2oZGCHcksX2Mw060c
PLy1J9NXkc76yPmHkzb4p44qRu9oeEOWYThndB5IGQOd9pUoSFj9BMvPmL1ipujMfUpkiqQLXvzP
kbQ9Y+gxK/26a924vvKUr07nWAFZrLodkLf7IN0Etz9jU2u/IuMskbc7nk8/7ks/DNKFae4L7XXD
IIf8Bl/JLDN3Jyfw4ohzuI5cJ3mMHEBA1oG1JYu+3SA46WFSjM8ldUgWvs9ad3RpXK9ZMpDqMcFR
awugXihGFLhlnIBDW38M5KKzsL2sadXpImZfQCpfKMS+uK14deNhrs3ME6ZsErr+7v3Ifmm0TJWH
2T61KFsn7DI63tmhLgs7ibo8FF4cZjP1OhbQRqyI36lSh1NocsRdK5PtR5c9SNZaHetDz3aMMV7R
A7q/ePFr3BJH7lM70V+Avjpvsky9s8tJxLW0elcvv5BBTQtmvarLyW5+L71HEqlTgX/zdWzfvVdD
yAYaq29lXQw4r862tL8n6l3DOpk3IXyEN1teRfptd1sGxxPeo102HokkkazSj1Y/oveqZ00Do+dj
jOrae6HwjzEFukUtVfhUfDvud3JNlC/NN3axjTcUjGGlwES3LVKbutGhb5Xxd9G7WT6le8iJQbmX
izbHJFjBYMp+iE2nVqe+ys6+P7CHOxW7tTF8Dekb851a5ZupH8kAeeE6iRuxZm2iWARAd8Ek4fLp
SmGL9T4nzhP7av3TrQKMnz84RDcjjtbtxcE0s2JnCtme/efy66qe9IL4I4gC6/Df9tXW5MpDxhaD
c5HkhLxhXhAhhzTSPG4h8MJMZ7T+qMy8YtVg1jqeZqmA1mL4PoppoDb9twow3kS00MQ12jTV+6Gr
+ydBRNvNUVp8yMl4OwECNr922RA7OGifzU4yQEiZ+q7XG3MWjvxyQU/HiSRNE3oDWxxozTUtP/nX
X1bDCttyXuHxSqh88F/TQRoifvmdbUjiM7A/XQAL+v5WAj8OxjDdcLoIOhzgPILxFvogi67EhrRr
ukacp4jW5CcmE6KhD4AUN3IP0U/n4zrSqwislR2Mr4iUpZsgp+c4EAZ63wsNe4s3XhgL978DcFHt
1yCpFzhiPAsDHmPDVvNVgakMJ/BqFBPu7tQP4Obwz9x5eEb+L1IBaXlPFXIDedX7kfnAzWF9RuYa
CgQHBk6Nh/P3lK1y64ZAzEmOdr63Q1o+BxIQDHgdjW8q0CkUnSiRReXVJJ+FtQWZ1zhn5q3h7JGH
XC0UxxOGlA6DciV23Vro3+NkTV+cA10z3ujr6Uj3Fth0hO1tycnU1cbBTEQ+9jzWE+GE+KC0/0Ud
cENPeEXAkDlZfx1vhpkRpKaINIldo3RhZUL5e/txgT3RZg46JVckwbcWPNrKLUfXhyI5dA7aJJ49
WKeGcNfkunl8P3vyhKnNxUVC+rlRZIigPl6P2cWr0Syt/7GK+A/IeCr1yYUkeXOMD+sQrew2kzOz
WwkwcBM2vVXjQo9n/hPQs8AaySH3IKwJsPr4czLZF0syc5UYXYcUf6mcv+waxiYltrxLXxL05BNl
y+FJRK5mpFe8W4Ifo1aUcJCOu59GA+kkXD+17DKcgEALhb/k9LM3j2NWKjiDxlm8DtQiMk2HbQHC
kmgJ8CC/hipUTJGeSL/2S0Ojx1gUlxL5lA+ZlizV8d5CqZKQHRvQu8CmTsRvwq8itA/0AbgGGiuj
vHmRVHPDpvrdjnuIusP/wQWYnKChtyPv/sfA0p5D1hEVBv41w6wKF/AS7235VglTAljU7QRDWBp5
kUFLOlDLKlVjcLKQ7El9A1aOhze8HnYp/BDbELhOq98nnMrOM7kiuYUPeqE4skhGspi4+L6VX71y
Ht5NnYA0jAS4rsnFX2CLGu63ORmYBOVg9aCfgmO7h9hldPXwK+ZUnDxrxnpM9ldBFlxXgx8UzPOB
JuxtHhCtbMeHcTRqCwcnEe8pkQE6ZQoE7RlQgfKpluZ7Ch7rs2usAqeEfNvFM29gmt/Rk83hqtyp
rC+DZ6ZMEtU0d1WXBWkAdKvsjowmKD+Bs1320EaEmb5DoYwEIGXKjUNxm8kxTo0FTK60MHydavU6
b9OmM/1SROSLeJjJRx7Ri8h8upyqOaQf9w0RV/pK36FutyqAojGnfp24hYOgfoH4tEHc3/l2IdXh
i5vKXKGIUGFllQidTICegqnzT/VzB3jsp20vzVwR77zSKmScvR1ibLH6fgkLwKhR/Glv9MoGWJiD
E8lyk8yUXP/AiSHoeTo5vn5p6HyiyEq6tHPaN49M36l9NlLPOdV4ksw/KmxGtPM0TRi8/2U+3N+m
K3g2HPwX3/ZhwL1vpV9nTsM9jTc/wP5IpsTVTA3cs1DLsXojr/+hQQ7csOK4zYideI5G57oZ4n0a
YGIMfTmZR6cW7ML/I7k0YN2HRlXm8LuxvDeYM+6OOb+PZbp/o+B6cn6Qn/03fDgnATEXXprP7Uir
wB7S8q1K/81mmNqaum78rP9q6suvqlwEwwDGl2Z2Q4DJjEchbjbqe4fZhCvuFlvgoFGPMrfDs0qP
J46IZb8YFBLYm3/iF0UAj2xadtsU3EPLGlZgj+zpmEle/n0Pk3HVTg2Yxg69b++BjAqontUZzyXl
cgNjdT3xUvU4B7LU7InbooAnipGDxLeCki4r1UQ5wTJ/FfVggUPyi9zCXI1tuDbO1rjSrXx9KeLk
5duNAKfVY0pJ5saJrSIWSuXbuhGrFP/4H9+qCcuBvHGbbH75FV+0ErsV8D+4BxpHYRtfvzqBrqRy
tIw98xrn7gqYBn69vbJCWofXJKl9EEvGNT6XoYQcTUTKMNoUYlQje5+fdznsHiWMHtpn+sT9lvSV
0uvB+ieAecqU7PptxEpHRjFziLSmPm5imxluMAoxnLG/U+pkX5jGWHg/4UCSJrIfT19kxgD2auiA
sjGXV9zQTZ299U6WcDsInpF2WHyjc/H+8SwogM7ojJeKx+kkQoOoFr3yr9FVMFCaXBz1tt5+9Zuf
Fu/2jxoWErTKmb6CfjodMGSlNKILUm2u4p9MoPm0QLsq7UVpTaMiWmvdBj01Ra1b0yJa6akzHdKr
IUztrnLe+bURTJN6DlnSTrAtnuhoVmQnzIL8Z0Is0FTLC+hIoxJN5z8679id1rDS3ADEzbpTWb4m
vqzL9Tlaxce8DjnUXCsF51T3HWLLNtCNY6FH3JjNAFyLPIUKDhbPNnYVHY+nLc/QqWWYtYWrHHvR
TGrqKCGGG4whJRwRcessalesQX6utUU1E+foHoM57Nxz1sfDvD/PbM3exyowcvpay7+W/J3UYG4j
cSjSILQJQkAOv5gvhSU4CShsdtNKd0/gGyDW9ZhWD2sbRvk0fzIpAUE9rN+rZe4oyG2+WnyNtisA
NAJlVwtN/tLdmQJp0vr0P6s1TVp4Zv6B+0oF+gl/yi853XLBltc3oClw6zw6EgfHg+uAJSZl33S4
0MvqHv/tEH7DX4vx3GxA+cIXalixADCiOMW9po2Dwr7YfPpw7R57HUhphgn5i2jaCbvVkU9hjszt
YtxOBdvYc8Ibrtb6NmuKaUYpIaWLuKDSmqqUqsgL6D3KWMwapHvWy7U7d3wN/mg2VG/SZIm0ftal
ptTA+sntiTTX5mUfl857Wj/CEIUAgfKjjOAY3+hEJ8ucQR3GtwQaqtuVDqP1bh5kQo3TfxihPept
XRLxpuYzcA7VQcebNPqHYaNC31oK1B1j8E8aBZFcAK/HuTTHAcvMVw0/K+7AKrr/Bo0ApLXFZPYH
ZG2wT4CF0jqtX6hi2wI5d5K30hEogQTWPiqpLdwNUQ/RfK56GDgME3bvGtycudiYpWhfFOfyCAja
2IKMmJfnW8Qsb32SfvJjkDTxxdQfJSZ2b9qgDd3Bd9SF/knTNEH2ndhIhGw8KbUYBs610+v9IAiP
nbisRL7rVx1H2aUgDD6ygb/aY5eqBDB7d+Dtaz2GDN3uvr4pliCSJE+6d6KN95KvJm8LAjC4e1Iq
C7jQ6C9h23ZiukKgt+rqLGFMGlaxKzgpUVhN5FXfSR4AlmZ0BmWI3SM5t1pgEGiKtUA1FT8SX94p
f+Qb5vmjcdSt44tzPY/aJFfR8Uwg/YW+wtwfoZDeEpG+appBcIGfzVj6a0IYuZseebmV4qBRPjzL
79ZJt4ZwUYld5XOu04lljfPfBkmc7UbSo/pfwFDTPKPgtCaVN2gbbU+hb2ESrGnGuCc3VkrP8RPu
gnwysExjhQxaUhnK3byKjNmLwuoqcWvSc7w19VfdUDBuqdnGrDcHkNIl4M+ROl4J3MBswtm1SIzZ
GhCtSf91yvuipvIqbuGUey1i75V4o5SoMOTlssNOGDSjXQSnu6l/IduPK3ui7p41n3TFtTJlSVy8
slH/VxLmglIHaiPyEJKqjpray8nyRzZ+HJuF0pZL8h0UCIjiMnlzREJUtXReVe+8Wa/CCPK/ngeN
fM7GiGFVe7RRZvmTjioHRUiRBLBooto5pUsnxrIuD5j3Xa4cmG6aurmd6efQyBH7/LQJMbie2ZXC
lhCeKRqmfs6SwG0qUUDApqxPLZoqWCqGcyx7U52OIAotb988DkeDfiPYlmkHOsRqiXPmJ9tpj7UH
8DJW+gWJycLUXndS8xGx+8+eyTRauYo1VpNtqWTjuAZjW0cB7wRFv0L8bLdv96eJoadJdw1QEPXV
pWEqm7a50k7z0BDYztGnT3uqFnlItU3Xw5MPPd0/Vci7D+jdYCr71Wb36WpiBfFQ0yItPdh0BXOy
MYrC2+T8Uqh3R8XnE+EEUeyBYk9ey5rkCzzx6C6aremWpBbebr86nqBixMtDhRTRXEuHEjqkP7Rw
c9A85wUq/MrvimUkGKljZzyDsl55XGrQqHii93UC9ksAmh98ldwBnc5AFlcql2w++R0Pplgplkr6
3XuUZEOPxCudgc/3Xwa6PnwERXgVN9yePJkKFvfACJ9jXonMB3ktLsPH/vXOqsCEIpXIE6i5fRCe
hPM9GgY6NSLFw3/t0CZ3PyrfEQskQefctgq6BJszBJrEY98AXLKHely91o45ygr+GGfKfvmWM/qs
a5nUJA46eRbUTFO340bZV1ipjVZGndEyHJxMR9UtRzWYNg3fqS+8HB87lJbdZxVVHs30lBnomm17
OQOEee7rTHeNrFpSNcBkXfDlDvW2mGcB0OAilXol25Kxw32/gfp9ZHGQA4+AgtTN7wdMwwe+CIkE
aJBnK0/ihoBMuLKVi7O7p5//3/0clM2oGMyu7Vb5/O1MZdGHp0P/78TACH9CGPWsKQ4HRp07CMLX
x2F54DPj/YWZlFCaokUUiF5FvqiHXfH57b8HRSedZafJ77srn7xnGBgth9bm6e/ojGCkFRvUw/WB
Md7NusacxeO+mPY0tDasmKBsxKHGoMAat8v8HoxqoCnbx28HlUkQ8tZ4F1MBQTnHqOA76uNJ15Ft
fK7C+wcMCScHynfgwo/v6hghz0g533SINsad8QVSSAO/d0/bcr8dLBM6QKhfy7wr2kkNlyWfSrUu
NgN6w4/ggw6l3nJvnD1cleuSRqa6siOsKFV37Y41oq9gLCT1psupqP5sdkP8LoB95E/Pw1MRSMyp
GcjC76b2fAZRGP3wbyVX6rCREwW5N1TnK419uRp5baGhyf3HyLvMvE/MP/ks1OukWI49eRZpwAhh
muobDPGOaDWC/M1GB49jdFThks/fqo5AmdkRgvboZGP8PcLyQgd+m+SrBJN/OUfSQOKS0wThwc2T
xheXlRUr7jv5zoOGMvodkkWB5havIDDZd8WMVr3xtKx+yDj1eE06pihQ21nsJFXlVUCziGFVgW+L
09l6Fx8wl7vBe0twPfiKRD4qAf8i9AUjGedqM0oXuqsddz+heJpuh0XswOlLLu/L3fPykMJl2vGB
SxJDmaFWF1ScG9mvddYh3nCOriI4QLKR13u5ckwD3zuLX07/txtLm+BfpG/XCa67QsBZjBnZsWQv
lSwen888Za0pRnuTI9bYx8Af78An9lxKhP3iXwZJmY7EiNj/cHaYfnSBlKa7nBxOYde1M+Eu1nDe
pRbCwEjRAjq6298q/o143wjAyzwemL3WZpXJUpz6LSImcOGCPuJsao6pxCEDCvcvu732m7Er04Mp
UtiGrkl7AeEQnc877aFj/fzpcO/UfK44Zp9jNiFBN2kUparLGrWv4J5FTsfv+xj1NYLOB7F4OBFm
wsQxTC7/kT+3YXFlJJvrVhtS0mh8XzNFILxTCaWIk3M95msLzd0kCqyoaifO0PBTY2perO2GDzCy
7osMImzOQyzcThDG2a0nECqkF/sqzDRnu5iU7vvhCLvikrg0yjKr7pe4eAeXgAkm44wmufbKnV/Q
19qhVOubHFThBR2pKUy/K8DXDaiLTpOeb8zHOU7gWSf0G+KtVX6mdBEopwwGsp9DxT+U8s2HS92b
q74wUAemCSFHkYhgn+b/Rbokd++fr3lgugssfwGN1LU1euWavXFUcG3W5pSXdfOxIOPkOd4MT5Ws
HfMWD1dkd4sJznIrNVDnejnnEh/jm8pPsH/oAma8nGcev91d1dOrlW7VzC8nKsHS+hBoEPJEUmy/
k3gJIkT7mQYFpXCbRHDEa2O6DBG4Rlz+tfSRYEuLCdvLVn42tGftLyDR4SnuzNeL7CTku7GBsd7Y
UB1ywQx4Llnf5KLoH0peLz7LMKRsI/Hc5BAFAxCxrnuMGmS6k36CMBBs56J9XPkHv60D4kWC8LCe
0bYrywAtG4Afqwjsl5FO6nWYQkG08lbB9wavwQT1me9C8bwa7x3LSxu2h3w3Fsu3XEiG78Uy4VGW
KHitvj8jt3oyn/gVRteU/ceK11pSEiptQdw+1KA4GADZWe7WjPKwYtGYIZaijAMFmuFlWstCgnLc
0Dy0hGVtVIEsJaYs2Cu/MEsxDLjqDNFPMLkyn2gJkpa+cOGhvsx/SOMxTd0I3PkHBi9WwDhYkOA+
hvLmvJn2vJL/nDhpSc8cZpdHHGb2TlaY/KuY/esszCegKo0YLmI78RuMOiEJy/3BMa2jn+XXQ3sn
K0j/7fL+OrARgrzwHDEczjO4VCm1qX5Ub1NI3o6+rfS2DsevuZU3t74OGWcmFbYG1NEDDs3xAaCn
3PISYMAPbzjHz7Ugcr9nDxZnhLM5NBuIWuqYDlWb751Bgu/WK4Pk9oFmIqs1DuDo/jnlvI7XixkL
pz/8iF1v7jBnpV40ODOhJdRc/uzQpykk2YxRM5cnQJpxDreiOUq05IkMvGKFTeVgUV3CCVkY3RPr
mGYEFEe3Mpi4V1k2aiD1gaSdaCiAY0udyRkICr3bFYqYulM/Q8dasEzNNz6gmkUxd1iiascc4eOO
Coybhd+8ePQflZ23j33havHfwM1EPIirV3tApmMwpDTyGD2o8HLzLLRtCfeBA8pqZVuAVft4+DRw
g4JRnSJ9tcc0R2shnmOaDAKHD2fKdSlvchZGiaJ+AgAckEi7jWXIjkxkft3Bl5es7+vBe+k1v9gT
1jgyTliQO7csQ7btaXFRoKvGOz3ekPD6Wk+0cr7xF38HfjyS0xohaKRdgAnbBnkkuuwcz+sPTwk+
t3eAn94uQDuZ8Mu3ODckGOIZi0CHW7tr+/y5nPYIzhUJglrwf9TlNfniZs+GmeswBYvcLDzNdPgF
HJsRzl+kgWYydgWAJ4dakMM564BqrwkTGPZp/ls+i0kJPsu3Gvx4X3Ns0Esb7Z+LTjF70MQcRzqs
i+pGOLG1YKzrB14jiqeY7fCKgc9lJKlixATinADaNcDj8bsZYm+D9GY+SSJ8y5d/e8nt5g0NecEi
B68zkw0ct3pSEYKMgb4oSHFMc2C745EfuhC3MYgXE6veMOzekx+WNapZcCQioFjguD3NG7n7RqZg
E07YFnUY/KpRhwN4C3e3cs6A3vQctMpm1ixLnSUimuX5kWPTMgYMFfYniMhb1szgGoZ7zZZWS3hD
7qS/Mq3TEf5gX8KDHpqsUh+bkvflv303X85ts56PloYH4IU4QZ3vGj73C4Ea3YB+y3ULZ0NBJ1FL
Fxwus/ofU73+S01p3yEeV89vsdWjQvH3wIBg94UoEu4vNjDNksctLp2D8OWd0hUFwHFPZGe24osv
vGO5zMDXRmFdSns6OwqvFhMM8lxJ+JDREbsgLdZiB81xcxdDd8sSZHkLkhzhujJ2a+jmKKn3bIMU
hRTZcBZ0topb/nAvYppqGW692eYBvma3on7hpyA3qBmcE4n7JBYA8lAaA+pgn3ptzirZ0eBM8FJT
MiZHyVwNeIbhbI4KXl/DgtW5OM+6h310vd+kQJ8w3An2MZGCl0zWqvP1mKgvQdZQs9CDsWSIynWf
JqBD4jeOkhAvT9wQ9ta1IPxsyMpvNKQI8gSgSr1lVkuvFO9rzOdI9+01PTls3QF+tvm0mvEcgGb7
5c5LchGILX/X1/0ztBEvccfDK5IWxScskIcP9rivBJ5PsaQuSgOzBQoEmzY4P+RslNaJ3MQ0m/Dp
3/ZAhptKr+wrHqD055SwTfN1XkmToKPzZUY2aEt119VwuTCmv/FD15TmWC7LQdIBGqN/bSqalPNz
BjDDDIAczmO5EjHeld/8FTvpdpwdkscG2R6xa967GINu1mvz+yvZVQBNaSsAC/f8vXdECa++eEXV
Mp/tWX8/VOtiGCK6lljPcTo700UP442vWpABCChGmbBadibm9vlRiVg+0GHRGHjSRhrXP0jUOBd7
wxObnRXIN4BQgSNvmOEzsaekP92ySOr+niZ7ky+12vXvf5fmi8vHvKXf5rYsYzZHzxVb70IRdF2m
7BAe5yzdTHoPLUPn3iQRBQVu9AH00sFVmlRvGVAK7zauoxgYyrlRAkuMcQRePabWvF+mft5UluM8
d9kHrii+mGKn+bYndoQClm22pRSWBt4XGK3zbba9eh4YwBFKuu1a1iJgg910O26QK9MivFafwbAc
KK/i8vnb8deLiU4s1LmkZymGpRb5jbWhQsohTPlV2VoH4BkUUl8z7Ou/F3ycl2RLoICcwATZz0qk
ZPmydMpOmEtCxbuqmqiSAjBC3MSxXQye3KJU3PV1UEnKopOH7I59ctDu+gedlE45/qLETnoRdQ4L
9ML30Qi/UxR55MPSqW30PtHVS9UDLp1ZgAs60hSPkGRsrn22kGlibPFh/dagt2ucCiX19/gRzAwM
QZsoKYgzTo70n3jggSc9Y7n/kLbl+SPx9jpKbgG9r148PCOVgmgyAMCQvjBrMYIP4EcniDO0oGOj
/sMT3dgsoSwVCcYyXr65ZkMfe5kHI6sWSmyIQoggN5EC+8jdfCIPKrOk8oMV1Qdrv6K32/QivUtf
7/eFOKPrhKgnY/nGLndu9XjIpQ7Uc0GuGt7x7/tOVe3N31+4qmwIt/l6yZb8d3SJ4lu3+xEv5g83
5Crr3vuepJ9F4WUIT4QqAiHekTh23Yssl6CiQhrFK8hgWfUNmynn2qKIYx2ZeB36TJd1PjbAqABr
jZBAjSoPq81MR3Wr4Bo/g6GXw/f45a7wmvYKck7WkccJ8/Em0qFnWilN2l96wSeLe8y6PR3qiMr9
E50QCl7C0gZO+mF00ZYLqT8V6ib091/QomBKfwfPAWv05Rt3M7ayaQTQIwSZgdwQapVrDm7VojI1
R0W743ULec8va/bdwbGZcUemWmbC8q05nCybRPFaK1TuWgUP8YgUo5Rdc87oNOniLeiQ1NRwibl4
45uti6Nou3vGoQWXYGBzD9+Iqf2QooP1h5SRSK993KiUJqs90mRi/VsNBXd185DXch5QeLxnQojV
/qaQ4gNz2vCu23SfBucXxcZksji6qVp6SIm10NBD1FOa1frGQq0Y/4GyMQLv8sFLnC8hINEP0dmO
ecmSoG0zUZMn8q7bHxgPdsxDq5YAh5rvRjoAIrUu0di8Mdb14xCSXJMHH9VRPToeWEclkU733vBA
kq1in90+r/cVUmLp1SZCQW//DcpbTGuHLiZqwOwrvtWU/iIfqE/4JME1XTS9jmum7We/lZ5YGAdk
KBPTLvU8LHV2Jx1TmVgB9pRWKa42RyoBat3VHJjUqJXPaEKezbo86aTN9AgeuUPAiZqwqepMFMGI
jLmYvKfcv9mK5kq1mOVx5bTA8lhF5mwXQzfHoC5RrHcZtu468lBaHnp2/FNY6Y/V5BBWAJCJ/MVt
zJPC7bxQMm+qvSBN1QrAkYvdgl+Dy3+QWtY00Rf9lOF3wxQxXz5I3H2OOYSRdh+0vN/QXTgda7dJ
b8vekLzu/zhB9W7jkx1toKz51OpvJ4p/eQjpgLiszNwxjRmCE+adOWPgu3rwZt6vWyTwNRIlBCo7
lzKn8nB9cOKbeohPO5Z8nUs1bhXrkjLlOxFTFKGh+rdQ7xFNvTDxtWN4SuM7J7ld1MnEhIuVrxs5
dzuj5GQg8mAwfkj/aJESCzajA+6O9UWzg0ngJC09/IegkkfZnfGSFvy5/6BWlBnRyswIFKyn3Non
r2VFClL3MOJgpgcj1iZdaxIBGiR8rbg1z0MoARkz/ITDcqAA7HN0+3G7dEwpNmC8musUetNRnf+U
ySiGxi5RT8u7KqTTQ8J0/BSutGFrlf6Fy9GGoFhglqAd2YJ8RdTsywRms4qdGmK5Zv43v8SNnDjM
WCPh6vtX5VQ9UYxu/M80a4lT5fgTqA3GYTR9XQu7I2q0pQy3is4ttPz5Vdsm/oEP/ifHnqe3mxyb
YzkJg8UCtVyDcNHMDsd5gUsfBbKUnGcbVP1L5xH+ib2cVHNUluBV7KTHgmSp/nShGboAofBJlnAJ
afCnWu7FoV1WB211zfMeHjpQeDzqq18dkQ8xru+i6ioZ4xDGPkL8pMiS7Jkkltq+9o2mUY5yoCNZ
MIb7ThI3QDTACcoFV58MzVMWxpxea9jPMAj9WPnak6aEFl1B/wvbAveEFT7xse0vFd5Maz3G7WyT
xthBvqNU/YeX0/ZycS9QoYVc3sCU/RYknAYTNbNWhiN3KZzP1uqYrgATcvuna5oaXd05JaISNdTN
jojTabMw9bbO40++avBg95+ahd+UDglD1lDax4R9IhszSH7JqUZmhtgi34janU++urHmFugXIuYM
fhNi69Ytsn5u3x+kfBioMn88cmDulZ1BzliKXQ+z3dqWR6DsnqpSBbLtj7ScxW7KrZdiaXpiywpE
+aCRfT65nd9icwOxjSMGxCrG+50gW4OKlvNSFrm1fCYLt4tiyO/JeVtrJEkLaDPKibemaBDjccU1
zVdLc2CkQhQe/mjcN9ISU9ResBQ9PnoUfITL269fGLq308sQ0mxu1wE1PH5+y4FwPacQz4HkUGfM
OSj8+JW8mUvAhtANuyHJrlWUO9OHh6iCOFeJqL2+fIkASE5ovXLjU8uMUBhCLDLD7YT5pixgkbij
u0DHJeY5hqQ/krUSqssVxthXP6rhAEe+96p5B6kGXlmCRYTZnQjyXMydZz4Ys+1jUqGNT8uytu0/
nslwO8aBPd1et5Xtx2CsgzXjMM7EQmhVwiUn86M5GmCH3j1NdFEb8DYb6ZhbmwjR9XZtwYigqSu7
QF4L9yJyAVLAPqlcw0EYoSb9+HtUh29c5tfwjkVqKl5DnEaJb0h8HdK8Sr91zepYi+fkZOM00SDd
L6bLExh4Kn9TF7CaFVUKlcS//cwmqomYsMZDCpADpLvqFUWHSO+0xuxDKlC+dJdG81a2A17arj2E
Pd2Anp1ILDXsdaRsm1ob6tc5Ks+udKL7ztpnts6HFJY1qOQFOt7Miqgmb68D0zaYXXT4EM4eZC5g
7dWb6+HyefLIoLVvWmQefIHVx55et3ylbLfdN9u7DjYbb45oEOHm6Z0Ag9mXDDoYmREtgEQJQoAl
uJ4LZGOi0EtwfheWbEk5frxUOYJ4P2RjVjY0N+1qXEj72l4gVMGTe/FdExLnS9OT1qEo5FpO0dqx
dKMXHic/RQyp5xgYCfh/w33Xm4BBOUKpHeYlz1ZxDdI3jmheRFDHAK3f4X1gZ9G88UCyHbqRCZcH
YqrNUMSS2DJTkeVe3C0RiyvCHHCKolLrX4pOf8C8c+Xzfsja0l53FTcqbSudj7Lo+U56WCDq5Bd2
0PkgYg0fCK9O0bv7PjrTtvSLqiblo1an9DWl/DhxeYmSXv80CJTs1yGSSKeTdVwTUihx09tuMlCg
Nivw9800+BpdzqzLy+PNoIYHzZr7scGDU9r6ymy9uWR2YtN85CxaG/OdZ7M17uqp5FJgd4nTc4Pa
YxE/gnBKzxhpP3voHjXgaLBEacmUpxW5S82VgpfGQfygzr5II3WfAkz7OYJbuDDAPEy+knzzGmBU
ZUKFAOPMH9c9ChP/A1lfert999CUmkc8gZgfDBY8tyxkFln8GU1/0gyGF9sYx5g5XYUfn8xvEzRJ
thvbB4hEZzPjqlNPQH4T7e86+yulM1IWknUJy84a7dQ4+yN3T+dyH5WVaX95gKldLktx7MLnBzwY
i199C1exBAILyFbc9qNFY++YUJ0s7J64B+eDw8r7I+H6DeQO8zG1Sm5U3RnDlnwqsn6EEpPGdlD2
hc9Ep3lTv/n5UzvFsNBTmwICOA3GakKRH+8NAr5EYFZgFjeTqMeDZDtwTg64LTcNnhlOQ657JYNG
r2VEILIN70MNTiWOSYjyU37m/m0Bhk3xXf5wEMZz/Vbark/l4GN83+Qs+w64EnROotd0I/FMO/T+
YaD3PDpRh85wY8gpiEYdjCcA5br4LLKMKEhzk86ojletwTeIQpnSbY+I5Ctgnx82GDweGC7Vn4rl
pI/AVkaCELHUB7rMqODdHTDL585LGDmYOOj+MoqeQjlTPJqfCsmMFJtqyrUSJR7sjFbfVc2FQAVW
osTQFVpoZfxO59NbYWeHtNtVRp2lwPZ8OOkZxzSBsPcYymUrL7jfIga5DRkkF8UWJyfJwacurAdX
mMLXAkqjVZ5es469AbXIV9Eo0pMV6KzDoynu9zkfQykkz+lZUUcWKTKubjf7ngtVvWnBr1wVCNhn
hADuWwRiydnIYVsluG6aUQpwT/H90jL8e3faUAywYIdJ+3bVROmxsntEj0VLSQzKD01rO2FP3KVC
VaPgJ0YW1eSwA+X3lx8xT9MgRKQz4po1+d2+fR852Uwf4v+E7KVOAK3loDgFyNm15qm/xDyyp+68
18G6ERy3Ec2J8ukSZ+LONjq7J0UItWTA+7nNUdGWQHK7pL7Mzk1Divdse0qhKcQMlQ7swQSOoxVh
HHwSc4kdgQG7b4ZUjwRptJW4n++oAikCtWwyyzBG+xv7JW95t3dCsPJ+0tFF44ogI5+drG2xUcwi
Au9NpCHovnszGYPBEfF2gvWy3tiG57He1VmXYC8aFhSEnJNMb+kkivo0aP0vpbd/wlFetZL/IyHA
6ATSUhFANsF6GorM1wel7jDWZBaTXfqEmK7h1aYil7BwRVyb2x570r4yuWvDh2GEKGeymcW+gm2S
mWwALeFYN+l4zzbuVEwD1aGybEbKSwRmOBR8XxVHDSuH2RJwlo0ZqBp017fBG6VRlGFz88dhvsKn
km4ylbjebXQ1bMi9DgVfDLb51R4otocY//g/QeujdLvFVM/m0UaR9BNuF6rLqTbzHjR7kGtPHGZY
/LwMfktE9dHF6JslRlRI/TG1w1r2/gxI9vNeF4aL7lqcDEKYvS9QOVL2vv89LLL7j1oVbQb0EgMb
nSQzgrxfk5U+eYMpvAQB4Uwug7XCgF7FG7SEBZ9qdWbUKsuZgJtghrKaw90RkSnbdahrPAASDzxn
WjnCzm7sSP9mI44AJ07GoP/mJ9D3L6kCDL9N3anhT32rv3ojTZkF905TmEVWdcNWt/Vf7xp8N/LD
II4BQ/8bc3adjJl+HIrER0KJKESScl2GSkypkU3+Q7nh4cBk4xzaq3Mo/CTyyfx77M5XPUfZc5bc
fNP7HDioAG/bZP3jz6qKwHmmmiyEEQdt3qEgejzBdlGfYOIrtK5dzlgGuZusJ8Sx13H85KJWLRjp
T4qJiyfb27V9guHa7+ffRRnlMrVyleHeoZDgn7Iwi8ntMbXrTA1GMpmxXD43UD9DqUE/O3bLX60U
TAXzzfJ5BN9bbxX4LOt3AMDcBvTSuEGw362xeT8CWW51Ic0h5oLDlt3IHFkd1YhOZXUOKrHXN8Nh
2UW/h7Pk7WFaqRVgitfZq9c6tBTmPuSYYPHyN2yGYxM3D8746tP7UOmEKHroH8kGunrpFSFEF4ov
Mc9CjS/iY9TAvuwxyoJySfSbMmLWvWVgqCT/KHXotoJNUxRT2iJsFAUOzlOGwQmWJaPLHKg8S03A
iB/d7NbnRBlmKOX8iMO+LxtuLSYdSwiOAohgIMkbpaOnOFX2MHrt3mz7BaNzSa+niNALultglmEt
Xl7a0FiLXNAQ8lJUfQV9dwNCLEW8SIxg/rg6cShnEBIIR4QMQeQZzOI9Mfq3kqmd6ppKNIbPJpv/
Po20YGcuUbFPG+QNUgxvAbso3yIlFC3j9zOB0TWLleOz4ZVKYTeqPHSHTzXC8ykbIwWPJIe7ZftQ
+wYwWaG1TAl3bK/4KjveoAv2LSLJbQOd8V9scw1jElRb25NEB9Mm4/b/y5a3fLuZVjaFSjvNiC4E
lDYs9j9l6Vl14yDswDGgJ0wOhEOQh6aNQZbpYic4YmHnDRosnrE9FajBycOdZJHBcyAedkAQEre0
OCQQLrHLf47UvJ/YJIFUAQ42/3KxQeQsNUPCv2OPyRVu94DppAPyYRYPMG5Zl1avoYph2YQIaNq6
yLoLZfbO86yCCmeyLfcRMAxp5QXGPLuPNvVDQXQFrOq/239avU3ZZwaobfwrpZctHCHhn53yKJk6
aeNHJDBF6HSEHOhyUgnVGwdnKfP88H357Sc9CkYGGCD1cObspcSSs2iy/wAGjwETGe8nATvKOOJV
UFVSiKyy7lY/wOI0iMavCS4jPlEMtPKW+Cco6UJOeVnA08GlsQwi5PgcjdwSk48lXE4JMKZaPnTB
5pbKZpXbHL6xWCYQ1PHzWkwrWAjynsil2sY46fH1XWvtqelwBXwg5+OjJnqxdsk5M8MNEtw3j7pd
I6DAZeMLPXPdU6jguKwN5bLsiWZGTXVSz1s7auj/jIQNUVF3xwiz/ciQa0KeyZv3g5mcKR/Rxaym
jcyQ0ao8m+HRzA6/oRAXFwaDcZQmEUcinIVAmnr0CO6RPnD9FBexQFn0XAlWppTniFqQf7hXM5AY
KcbrVeCVo5Qr2BPkD1EuiW2+Fp7uwHqCqjBxooTzDyPnyFT2H9TvV+RXpW2Yd4F+5MV6aTXY0/W0
yzmvnHA5Ao/FUPIQTnATMIdWQJK9ZtBBB4bf4VyNQncYQYtNqg4YAjIJQtoeh/cBIZ0yVT38QBzz
siUsqAqaWfcDHSM9ulDmCTboySdKPMUm+hrp4CO7RgiSbwnzn43dpSf1Q4eMChmSnOGDWip+tUN3
vcr1h1wZBcnilL1TMCFzTApXlnuu+1ZCFpcAdq1iYK9rBb2wauE+7n/YFqSyr2xWJ4H7rvkx428D
G0GMxQptp2BZzzywvj+jgZfHbQ4mUFnU3UrNMK3rXurDuAkPfb4N3OfatClg/7j2FrgEeLTiJLzY
P9fGw4pps7cMfDuNte8UOMDGwArEkH0wEfaONe1/cULDDMR9eIR67PtE/vzFDdlvObd6kWpd/MwR
7cck2MtYLjrtt3yT65+26H7/1EwF2xULADcZDiPyZhEgTMUgQyU72u+mi3Ijog1a2cs4pE7UXpdW
7hEK9mqXONoMKPFL9gusX+emiXwtXvbVWKfnCpLLl+PjG9qpSex0QjHWj1g57uWeXhVVcwJ5dl36
8A40BRiCy1bok6lxQFr8N7y7VRRPzqEXDM91M4H1t/E9Ti9Ic5uywWiZXym3krLpvR60IvH29ZrZ
ZAx2VHMGsFXVh+VIWnPDMn/J50meHd4srUogQZ21W4I15AURthcChPV1ZCA9pPWkMj9W3Av8FnGE
4Dc5Rhx0/qaS7LrGogP8i2GZvvneYvJyJBiCFv8e/gbcf9XjRvRfhQWxdtrkAwPOk4XGMa7yzIgb
jsnnRJTQ6rlJMyk0TuxL2JEFGJ4tfTJSyf4c1DmCnWSgE8QvkQOorGNqz99TBrrvz6iq8J53c9bM
f1Fbmc7WsaOydRWdeZFR1uYhoc0epZggoNeSB/d5o2MyE2St7LTIZDE1PSBONkKzEKKIHzT0zZwz
kXrAMPKhi3v3Oy3TROuZKhz3WiP8BP9yVH7iootW26/8whQ7AcTWqsv1TyO4/mjCCsLJXK82rCGZ
oqWdK/5u2tf1wPOxtV7bI8Vhqt9Jme9AFH6YbzMgmpBgfy7AV0wtj/lc89mU1z4/g64hxsc0LX7M
AesVLffScCdC5BRmQkFYPKmQORmE6RksuSxu8FTMzgcpzmOutCJpkuPARWYtpq4bplW3RuHXEHxV
zz4VK8/3/LJalDRI/vgRHSfzEPfctjfx2+CoO9Bp13LhZAZcUUtpsU6zY4B00dS47nnmd2ttTWyu
ZYCfLFo86Q2qgeZFo6tA4vVru047oWQRQec1jYAxavSSQjqIXAcR6RoFIZgMlWbx4zR+bp1/fAie
475olGPEHf49vpzClNd8YElUzF/DiX0+cYww3kOEq5bUZNPW8oybVahtVYU2nbfQB97xyOhPvlmZ
xbWaCCoOTDk18hIBArKhEJNnOcd0f+/HUsy+Z+6yzxq/DivOwZcQhqKEWLvfjLPzdPYNAcBTbaoM
JFCsUopnko4/K4UnaB2COvyir+C2E2lQbR8KU39QhXuP82vKFTxhLMdjePH4l9rjG52oZZ2bbb4a
nzJVhP2ffDhk0qHUkuCB5XDWQM3MG57qYlTscj2dsS28e6tYVeRFjRbDnLyvp1a9foagqUXEXdFU
B+hKiKAJRYaUgaXq8bWSd14y4V1NaV/7dVJBrY6VDzggGQV6xMR4ruwB99QgJ9J2Sd06CImrM73j
1baTlcWD1puIGGl1opjkc8Dzk0UrZ17g0yD1P20F8w6GII/4ZSNTqLDzx9SzoYKHyl3I4EyDljZ6
8IcscWnVyDWVwwilWr0d15NkqeHseZ471+XMRp4ACfdaOw6D4CiRdSS1kycTC4ss6f4HiAPBccQC
Ho9D3BkFOKQfQzZVzxHp/6kPjLTlVu9n0fxt0NcalekhU7Tz4E6l0wBwP1njlbl2YOB+SiDs+Pg7
VI6pWFgcE8gkUpNA0NeWTt0sBU8wbzka+2HwRS0hgc/BK76nd6tXh5k72Fe4+o+HWq9TBSVs3YNw
mcwoEK53UTgs6P9JEG1FR4TkrXiJ91uys7O9iVM4K2a0RfJ+zVGqbq2rIU+fI0UzBHLgszl0ZfKd
TzPls+dE65PfNzOBCyrL1jAY9yPdrW8POng1431IpA/IwrCSsLcwPPlmOg+THeHKXfKjQa1Q+g5/
3vVTIMRdtS8k7c3WGCqA9fhQf7iAwGRDOXuS3rNwEco++1dl22/PMF8+zBFidg+gPdbfHsEa3y96
Cqv31Zd6xNDnw45fPgTpEiQ8ZXRfw+vnFo8o8s099CitC+ccdk7cgaox5MEF7JgINoisveP8SxA4
pjS/2mJuhkMLiUXDikjmPqv3L7zHILVBCL+omclhoNdFoAsSDiY9W4RMDtwXa1Z/FNpM6vo/hhbe
TpFvYu+70VYMfkR4abbG1Xa8/nReJkMzQb7OcHSk4f2REjy54cRs1025AHk2gw8MrGsCcYFMIjL+
AAVUNaDqKyzY+EjIVdwAmrOK1XrVwURtHdpubp2GWBqPD9WarTykv3rA2/GNbjhautzFEW53FA/E
CBIhJyMUwN13Xkb91oDpvnFABvFFSftKpoWXQZZCWHpxetKdD5jWxfpWHFkosZKDJDWtPoAuk9H0
Kd0OdmvGBJIjzLLoV/uKCoVGiGRoP0n/dCjy9TO3QjRyx0BpE/pCJYJwZO/AZvdNopZFL3iQ5u8K
lMEhvoPPFCl6OBz2GvZCzqt570iCIMIpXo03dFVmt+7buZ/2IsS/A6GzuFUuuId1yony4/QnzqtK
VYi0C3QxgmK/C3YNKism7NjwKpDfFICA7FFk8s3OIRFNfoh79rbpcNumAqEVxtvQI3oRV3iImSEe
8UrVWay5+iF+X49ygU1spbkDWt/jqvVi+ZXC793x05I3NGKLm0RM/c8zUz87eB+2PQGHAkaaylPZ
VD7fKG1Cy5kqiIbxab1MW9eIVjslAqTqIXGk8jjx77Nr2mzz1Q0EUNxR54qQqucqaVlszAm1w47q
OMqh2dpr8U+5i+kgGzzNXwdu0dxffX9ZhKP2m2cOIY47LSzZf4qw/xUBUPbR7LKC6S75eYPt1hLb
04Iof7DtPV0ZwLGzn1NLgwzR8OcOni5IAUkj7CedjdubK0j48vazPkGGN9wBIlayh4ue4fzNbH/X
LW1wydkoONs8tmfwQO6/3+e0GerocJSvow5Hx2XKEn9tFKX1b8kHxJRWsTX2TpzfzNaFVVGiPJOb
n85oGhRuuSoZ8Ab2MrHSXmFoLjX2yD+DMNSDX8LSeXJpw3SmhwR1IOwx2ipPO7qeeyznic+PA1Lz
XdfUV0YpeLkP0rxVBIIl6Eoo9GtVAXLddEzFwcFAOK3JAXLdDiWGpdKjaXHqzs/9a8HdiqGq/ZhE
/TVkdK6LBsqDqqxhejxaDURtkhZl0ZTJiHnWFB++Jrkbmm+sc5SkKX7/3kgigz1lAapV8zGabU9D
bEjbJ1AkKqLOtbnkKZ++jqvXBCTl3wAn9U+gLYqQkZhFbJySHHY+vNTQScGjOK88sO2yjg99M0h5
az8tv7bjMXbxoJA5qqzKs6Al9H3NUwmzD7gTc4sGWgjx3hY0hRnx/b4TInvvRe4ZVv1UbhE0mRIv
JWFJYUdQXW2u1KboL4TO24m4EsNx4qgyaSvDv4i1vfN13ZEd/KWjNc+DCZV0lLbNXhAjejGXn1fB
51t6BA1rXZmET3NZcn23suGdY78jiaU5y97Fa+p9OoCURxvVZU91lcWoopM6q/mueqOvjHWwbCVi
p+8irCJWK7IdgG0LtwZPIoKLcs5i6zzjt8WUeaFNRSGeDg+UHasCUtAX2696kze9ERtsoQGL89Mk
cDig5aYc2y6LcLJwqTMMgpHdlwa+69S5F5PjZQcSH2/CCyKp+e1TtYsFilzP/MxFsggnvsvzMOq2
UaltdxjJNWyh3fZ953l2qY+AUCAVywQaZXcKdHuGHL5imvPGXOtyfrUBA1irvjMlvOqz2NzWeg/j
I40XAXwSGn1+rY6Pz4PXcNhEQzo86imJF1U8hB7zTVbh7Nrhtae/qKvziVIer7R3vaWbCSMhf0jx
8m3bfccL+2b3UrYaUd99JqRvzV8xwtME5EBgf8Gs20LGCd9CheAccqopF1KqRPAEFbFMe1WS3EjY
xGEJ+NzWGrf+vi9AcPfPoMawiHXCFdM1Mec9mEtDDXVWigecKTOGrsHwqJmOcNwXvMqy0nlE7lSh
aslpDHqseWN3vaqziEyLaTHMlQjkzFITh5YKyabQb8obA21bq56ouxXq3FSu8pDbj3t5JGJgpz2l
rxzQ6m3Q3Tc2QAuzu1MOHhdCCC1IjFA4W74iLBGv4RlG4JAVTmW0dUuB+uhB3wmAoxhUPqNpWVqu
I6yqXPDiFDkSRjA30Go9OLDKW19wjDwlwfT89tOuRKJ5fGL6tueg1kdtT+mmV49AL5LNeyiIZPYe
O2WzsEa4EopxZC9/yQcaZYZ9a+feoFK0ed6vg3IZ1SyQx5KTgMdL9T/5WSW1yUTy+I3KbJ+f3/9u
si+ySb8R5s5GhxA/Gd1C7bFArH4qvBO1VFByFuwbSqoWP9L5Z+lZGkCaoQFS327zvBIDOB0EkQT4
ZOT3o7GJVChPjLZEdP+DzGBK9yYLAmVlPgTQgT8eWGNwU+RjlM6O9B2Bx+ub8cRf5izKWX9O4Or+
j1oJTOkCFEimi86s3J2Vn6nuy+fH0UAPB9RNOpppkVmFqaDzvHQrY38CZhUi7oMT9Ksd4E/OsYos
TCwVAK2k7k6To6mtCurTk1MCERVDG1JZ0+PnqR+e7eDFUv65Q4hsdeRZnLGg6lBM+ujT3FmLMlOr
BspF2QOOKN+d+/JD4Yp6xqeEMsXb4WCnFcYTOPueOPwyhVFjxoSAbl7VeKql0wqHbFkr6xm2qwZz
UeiwT6kDNC/TVrsmuRZFW5khjgdWOht5RbHNes+AFWaAlsp8uYSGM8EtUlYCF/wiVhvO8Mry7LGy
OBH58hevVj2vrQ0r28q/yZN7QvrH4dC9iGV/V8Tf5QA25asT1H7a698W4Fd4sesnQnNDI3KIc4mZ
8pVtJWiNxbZ9ouT+5mAqqnYpXgFl1fu4gYe+kU7EMLFFzN1WYsh9R8X8C4n3VBl06gXqbOOvTWTh
OFO9rLFL+Gzy4GJJgBuTUHKVyrWlgqUv1lb3rLySHsFINS75KUvYIM3GNr1RSOn8NCJ2bXYZr6m5
7JNjv35E334jIkYWb/EQ1zuKRqnrEKI+J1CHcIDx839wMJppImtc8ZKFLs5KfegsSI0qBx40f1vK
u/2jE4xFx9E9QwXdi/1KB5aOJoi8ksn+V6/MrUTtNOjZ3HfuzNokNaCcFA9RPP0XDdLj/hlDxmhH
OHN59ke8RZ1N66IhO5rpv4x94GxoMDXqT0+5+X28ZXMtElovya90/Vm1QWZ0MlZbiWIXCQ/dbJyX
NwiOcWIu0xMFlaGI5fguJzVcs8wOAyCuc8wvkfkhzNXtr1/0JRKEAef1oybQjoE/QlNZ8tZXSxwj
yC1R9I4KV7egvuo0iIG7GRJu4qm7aH+O0nSINwmBrzwhuf2bdXMgeXDM3O4ut4BHv2cqla1yMOHU
mh/jrjDxDH7LBT5laXsgLSlykhFInMQnBszqmpvfWezGuAL1Oujgpe6qXYFXMpPdSbmXjZe3eTlJ
6c3KPKxq1ip/ExE4t2G+YctNk5RKrIOLBkcsal8mLAE3Qjsgbyt0WCFDGU3APsOHU1QLlySodKGz
A9AJRR9pi9cVO4qQr6JCySMEIxtuP3Y15GN4dPphcVdY84aT1lG+VwL2vhkODbczO3eWC0glqKcP
UPaxLP+tgzY7t8Yo6eI5QBBUc9YzyAU2r1ZL74waH0fJQnaLZSQeJF4V65Jo9bm3+MreyYBfrG6q
cE5Vrgr9WRT2qoPjCg1IW/U+JOdy/AafRzp0Qz2UR3W013dkJ9LO+yeMWG2uUrUA5blpqovzzF0C
ls7QETKiSbGjvv0uBO00WGMumIKVR0eQZCmD4AkAUQVjAxKmJREseYO+QXbWz62P49y0MaCBPX6A
hwm8RCPhz4axDRKZuRNk3uxiKyHDG5BeVlVP3dEcn/T441zQpS7e4vPLXP/pN98i37tAyP6bpICH
fqMufCYuTeiCXT8m7pETAo0zPYU0hi1je3StuUH8LFdGlGJ+AezZ7relGTpsfdGEt0dxlZsVWh0P
tLUTQnzX/cyVfvuz1JQYnpO/355SfRB8UD0CjHsV+kSqw5V0QWWLnGXmbnTI8zd+JV98Vd2vzryK
QLWUDRYkWg9OYVBcj3GXLht0VYcMd+Kw7fuogi4RY2/nDc7riIO5SlHWVmsIESqo2XSTa2G6ynOD
GBb/WC36bWVQnfiCkPkW04QymfVpD0Ki1t+M1cFt1wmnJ1+NetwEl1cyUGRAoyGpZD+fd+i48uIi
l0rp61HeanrgMv52ql9sn5YuimxW47Ria66zl232+QHb0HE7n0HwtTStool8rSfRzV51Z+FAc2EM
Ico69tcA9F0InJ2vS9gsLSHabfAs6GVkmgpMiIVNOsafAakXzMc5OeObeeL1UiPPXTTd6ClhFULK
ZcTAqhIxXKIrZz90duxOvHElIS52Mzdi3lr6g5glJnogBuf/rfY0lMow3LDErMBut+0WGrDcwE1/
H4LAg5WW4i3NxajLKKqRaR3BPxTBnlyIOvUN0NfA6Cuuh8Hpz1ry3Q3ySzqb5IhDYLafQvgRTsaP
I+rl6PTDuiUVw1zPtZ4gHkBp1efjjphcH4h3AZca2o2+H2giocYiMoXdPrp0M/XjVaUM0xM8Boc2
VNIIwreGmIjPaZRFdrexlWCyEjmUf7fAHzyrShn/6SsyzL399kyEEc8iBcNt6l01n8EIRkyiIAj6
O/rptgXu/8+sMcyuGGLzKtEYnCfKo7J3iTiiZY3FGO9nlZ6pophW17JBTNYu6vaD02ttCk0EB56Y
Yg4pUs0eOUR69d84ND+JRKlpKJQXJYuN3a9kRqGOj109p2WQLcnyinhUqHDy7n9MckPtOaF6hiin
zyhII1VvMX2H6jD5Tafln55M6e1X1P75GHUleb5nVH0axWeFyeaycKHa5MLKOrQsk1oseKHK1k4x
1xA3BWAqZS8lLNFhXJUQpzQlaQbXlsehteSqLMtR/15GOcY/WapvstXYDvn5VpIOxvZDn7do0uY/
dzD0YgW1Pjpea6e+dzTT9mV7LluKtj20awPG99vSJMPqRDgisz2XEdooyTIuyRzqYDCNDJqSl72h
vV67vCOZFdEWnFFHKJ8Oz37TsCrscuGJWH8YZUBHKxt5BvAyfUmt5EgK1hOHhQk3W6kJtDRHzODy
5KcaNPms9pBFcYjs4y86II/POfpJVKGZOQ1LMWYIvHWUYalnmXDuuy3VeC8bJOvrhBAX79ACKBIZ
unRclZ8s+anjq/YhyGre4NrWEgPlY1vZUtxJbeDBagmDoBv55ngElmdCrXhytO4PYOqiD8AI76Yo
Ds25phTjG6FJds7oimL1qRbUq41rR/IuJWtzhpI690bY3W+seZXo17MSptFR7xi9pKh6NJOX//2a
Psi6Cc/3sy5BfyIjHFgYgDc5Wji4zUmBs0PE8V/pMXG7Lev1mBSChsV1/RvkmYGOdHwtRObogsjU
qkTHFRUOXX3hZQshzDXE6I97E6mkjusfXqzF2S/gMUnL7+nuLctTqDtdm/7hJ5Rdes7XjpkK5rs+
uihx9Q2NiqHtqpGZnq9VT65Yqsj7czIUM2gMYE2+1GrL3x35o4oOpmxgu0qQlyDoetl3/ypec+OW
Z0tSw53ayR/RhHgNa8BKNzAla9jrljslPD/27H9TETSkPkHR9I4htlpVlNi32F5qrGUhlaMLLhsZ
EPAFVghB2pivL7bsdKvdZyylADWi8L2VPwmBk5ixzeBbCedjoYDAdslXnNXSAdASmZBNO9lEdO6R
PP7pFXtDn81mc7WiDBn/S6Eq5hOPLm9WYVhOJWYofq9y94ntFXtCXJNzUi3zGeM72SC8kAWrzw67
s1zWrB3kuReWV/AwBwT1oKexaQRmCujhHLsViZjhuhflZjvIM/MSb+38Mf2Ht1LbSJwHNjWdwk51
hHLBAeuTEWL+Z/deCHz//HMca07p/XSzmCnByIo3o+zP0pXN8ofDTjf44wYY888641BkuAYyS1zW
LYJ/qRO5hq3zz8Aj1HqCxxPMjkQucRqwwuo624zRM7NIba+KTFXzlwCi4i7JJvRhW+w2+BnKKb0l
yVUVXdy6gWKG9DOBv7noPfirQgq4jCgt3bpCFIp89HRllEC6Ks5NjRkzgZLMWxDGFqBibmnS14it
mpzH8nC+EHfaxMWXsVNUk0VdWtUnopbQnWsi+6l2Y9Gsh2LCFOHIEn9f7MRVyCwvgkPBtlr++Xll
pMQBjsatN1qZwlJLpLtwqTxKp8q2jO3DESK1meTYd58AfL8EDxGtMTJM79ya67FI6vx6CS0GcdQm
YqnM6JrK/cGir0P+pnnwd12jlNDArdNDY4mEOWen8P1HG8LBGt2Y7zzGdK+AcSsZYUCen0GEX+aq
IxfWmfIRSj2aJuOWiPX4DF3B2naE93sYm+zVc9XkpwHASINILJMQeGIGDo0IQhgx1tuwJCFgdDgS
iZhaCbYUY1WKRA4erqNcAsDj9+oWmJ2pd/J/wOPG4ZmnvkR5TwTU3xU2ojjVnonwzzTgnqweKCHe
JiTQgJxzl1qCCCfH6c6het3UfjrdHBJ2r5oohN23/az5xrMREP+4MOrq81QrhP8sCoh+LXt/bwaX
guzOZcnSN7Np2ur3bHYun90qstzSj5RMauUEvOuigfx/HSqqBwfl6YBbJMJjplsGB9Yui/ZBEpYs
wlKE1ORJIqp7325GojMX+ZgoWK2szybaw3xr6g7V3wHr7GM9KQ+/s8MFH/4OtPd3uB48exBKp8UR
tHgNNQ0SDkkP24cFt9cGMYYSqMNkQt2uGhL50POlcursJb6JNBTlBM3m9h8KL5R7ZrAg/mWEZL1t
zMsgyuA+fdj3QiC693dJ24UA4jFVk3IPDEsyLDh2LsYQzY8s3N1QyD80gZOw+XTfVLVJqEv73/i+
ZlB1YeK3iexVzyT5XVlnCc7bOJJBD08Y9dLxyomrLL7QvE/UUt8jjc2N5oEaz0dIR6jzsospeYqF
D2sw+ryeIt9j+8daMJfV3OZZ+cBt/m1daFyY+5YWYML/bB7STP179fLg7PXHdib0C545PRBKWEaY
wRNWbBH31dEifK/GTuph0h4DUKooNpYNnFD7c1cB3bqmX06ZlECgY4SYzhYHCteOp99dUrBuUc9t
eyQS2K1aROB8SinBNyiy984keaiM6oZxuiomrgX15+4LSEXnPe/hOR/LopOP+FBCQUu14/x52BIE
F6i/vy6aaV5sCnG9be9pBAOu1ADTxK60MvMViNY2L6HSD3RSjhLUZbfQFjJPIcZmN7ZHPOrVvL2w
ujJd3k7CdQau4YQSqY4l95iqu2QIyMdzxlV7h1OC08vCLYRqZsYY0aNkL8yA84N7qQOea5k0JNE/
bAzUH1/FiETxstzUNN0chl9fobiIQvLBZPtG7++pP7YokY+MfwWkEBFYCWsYhqjpzdC4xwisiq34
gs/7IkcmHXTvbkx6eQGOsvvJhHc+1CQx7lrD+U9nPCVl5ELVz09in85hjKA7p0bDEXphQgl/6iaD
ay87nvurceizTv7NGROTa4IG50tXsz1nw/kNi0PmEU5SQmRal3qdm73lD1+bVZROYfSGh7fNuPjr
1k5sh8tA7vBJ8sYKKGrtwI2cSm3or9GwrrL1/qZZZuW7FdLg1fRXN0owsIaUR/xa7ncCcdqt1A6l
gUdoa24Np3wbZIUUjmVX/FVblfyVaVTRWoViR7exdbcCwuABcbWMpn/8UgkK8hBvSm1JMBZP2ii0
9Ms0bmwAkJ3Fh4TNd2wPs9+c4eCpGxL+0147U1Yrc/PbfMlb+0gudwk4GfarHBzGXRyoy+fHQyU9
JzDHK3mGfPL5+hQ8OpPSJirq4ZaDFZKoVobPFkugJEp6dBBgxc0kpQguW1hkAOq8oFH8UdCtx+Hm
KLAp1r3HHxqABzgQHomQvlUmzh4ujXp7PLiMwYn+L4UDC4reDQkpshg4x8BjaDhsLeeg+C7FkQRs
ZbQ7qqneHxaQZocpSTmURudjJDXIFJLu3bKwAuWI82Z3KmrNYJ864CODlK3O66V42o4Oqd131ZaH
XY1ptrwXqiJ3CeG70kcvoO7lTxmx9RuP3QJAwgjYs2Qu4Ct/HOGU+fbERNlgRjwKHp+h6CPJpsiG
1GJfxDgKojgx/N6z6tVaHHU7xQYHRrS930zGAnmXecCQitKe9dvbEDo7EqULWwgwYzg+1hwRcC/0
sSr/GlIv88LR6wrDXgzdoOkIgS1CY4L9TuxEn8+EtKgoJWU5Gu++Jg1Mqic6fnDrotljH+3txB+X
9L6hFBA9PNp/eoQvhC1yuLzNOD7ihpfdZiUcU7Nxe3CHZbYxv4W3TLkDRuq8WyftN8pBlJmFKTQZ
sjzt/7JR0mva/obHxOI1W3xbef86GjcqewKGfh1h9x9nh9TjTNXj2KrQ7ucsGu3akAfKjwO7MH2W
4icKeWa2Q33EJfCF2woOqxTMm9Cdd9MJMfswv3nfhosJWqrwKEttFdBF+J5ppVqxQs7NaRBnP7i4
itjNeVNawUKIxiPvriVBkme+iN72gRSX0HK41OqJBYOwfFKD0Y7SK+cp0xX9g5n+iaH8xkTseVpG
lGPMMwWiQI6860vO7/nigNE6gb2o/ZSRkWQvZmrTx5SbAUZWJI59QAbd+LU+SmNRus+X8N84VUpU
i/MW/tVt219mp5pOiYvnfI0Nr5HjDyCxlp9hKR+qo3KlW3rIYe49QeUSHCGcTbpxeyJ2VpBZlqp9
5vV5ta1jWhnWmOS7FmcbV+gr/rGlM5PyGjpVCSEDv546P14nDaOeKkSTcqCiqW+YjUfc6kWxSTiN
HSk7GPQCkQ1n8TyZPq9KL9rfoytf6dKV8hng2/On74apwVHr3sAaZBCzQlurNl/GsLp6Nfp1QJho
J8SIqW4W2774dVDZE4cZTPrQQ1VCKqQNdfVyaZXbPfUllrgvCYm3CpjzNW5SqhV72iOvBvGyEa4a
YITSFzmcOumMRAfTuQTbScjP8VMb0EH5knRMzhijYzbI80VcOEB46AGqQHuF6Xf1DsYhrdSBBO9z
pq3e45UvdDTGA6NHcwJ75H4JmZ4/ZaZaU4rYNKS0Zdf61EnrVau2wE1zQuS8QS34M3TqynszYe+i
zjtBLmfnxiUKB5QP/thpfbsHbxV3PTSAiLcDvO33e28py05DNNWwdCZ4KDSS8yrtwsikolF/GMod
vyfA8xJ2BYGpOkesbu5q3ccPak8Z8jhpwMpRds3OA7655eLmTnsftrU43zpNeGEPuNnN6jf6IhaD
sgwefq13TIHjgPFd5LMXpXDTrQ3gDfNtkm+7Z9ObZBVrKL+4psxcSuU1VH0AAn8CiqJ6m95mu1TV
dI/jmIUtx8V7HvWhp3T0VfGA3jK3pf1Kb5vKR8eC0oYVqEoGre9m2klDb42SBnsfGl9v6cFQ4F3N
4b7scNEatXNFmLnnyCNfR05A1E5uybOa9fiiz2Gl05VbTUabIze2Pxds2SmQjzqiSGOTuQNpdtKH
E7F+pxSW/3u37osN54J6RUwaBD9s4fR4IAPy0oET8/+qjYG3DS1VBk6bNTE9Y3PWTu3AIZF5uAVA
BoANQGc8wzknthf10a7hAewIZGPHTUabs9B1blowhscYodpOyN2CEzBHtAj4OFGnFpU1Ulh2hA3f
Wq5X4njtQCNrfHM40QXrXZUWeJx79y+7H7MAERI5RjZgqFMEktaAg/qv5OGHu8Ay0uxKuJeqhysw
UDREhWneyTLTj16SX0EBJUKjvpL4mQEiy8uscLf5LsDqcj+Zwgyr3V+HOBVgkvh6PTO966m1wVdD
mFfoleBzyRvef3vWMGKQEqZxgAcQshVVTkgBbggcHns8oFNIvhUbmWbDoFjgp7Chr3Lv50LqZwLr
pmw2wGwajGvN4w2V9UHQUjUcfAnMjahIYqQi4ch24zidVjVG1xqZhVBMB7Mg/1CvVyx8VI2Bj89L
a30kZsenhdGsGRLZPXiapAmwrTPLfLY+4VynTrp5o3GUrw+YY6tgPAh8mnnDU76FKU72O1ZMNSEJ
JUi0sqWaPBaAVvl4UC+/iEj2vFtGEmzWf4ZDDBQhHQOzS4HXzbnOE3WFEoGsJ0HxTn38dSxSlWao
D+tlalpXPTrkQNX1ArZnYEcR1klEguTZOqrF1ig0wlf0Ju8eOc+Ukv28VyrfFVDv6yNiqHDmHNZb
pXm/aN0RIbvgcvYdVSuXkDatAcwa9Y0Ik2hN77dpyogm6cE1+PhJndYeER0+PLL/inN+MF56GHEP
gYJhesjF3GlPJixkiKGU2J/uYS72XssXrJFqSdIy/gL3oY4hKkaMeHg8fl7hZ2RBAinwozx5PuId
dmuNzVwGBLRt16gftRMegbiJ1m/VERzA03ldvOuLl/Y9Xr19fqiyKykX9JDkZ4L4aTNqGk7bezXf
qp4ltM3atl+cBcibMX6cwz7G+WpVJO0W2vXbGacnbKbdEiiDEXKAJSSBHBsuBHbArfwuqHHOTKQa
2sPh17LqSRiCFZ7V1thNKgJTdtGihYmZNQHTSRseOGrc9aDVloHJAn/w4CmjhS6ZeSdRVzVFSPyN
WKtko4ozQIXneUQFEuwbDau06d5Q41WalCsqqnvKwtkewlrw0FKeq4Uwl1nD6+HjkpdDLuu/WJeX
1UV1qLq2mO7acwEQl7rzPOWFFKLhgbFRbuOPDmxWSIE2gj37We+PQUz92NLIApxpxjOLOPwKHWqa
0cw4DD1xri0rO6x6I0DOifRSGfNYS3bMjsctQugf/45WF3RdwqkkP8fs/5e89mCbxRF6rqhc938M
XdX7os1DEH+pY5vmT5NsyA6hd337sOgfRu76W5rcpfRrlAUOG89LPNdKcEgopnJyX+dUvJ26FmuS
/G7SjVCow4P3NAvYRBBmKZosJcbGXUbeVqZXYbXy2BHXyeBCKZXVObpVo6XspV7s1sDkkgawT+GH
sMN628B7f2z12Aj8NieHUWCDR4MGoV9Kp+YXS8RoMsp8xacl3ptxu2yXFO4jkL06/uoERWcXOV+O
jLXmSNT2YmxRarIfuCB228ih7sW4sXmYB6I+ID5brRaAvAKrHMsWyFFhP7QV030Ccp2ZSkesiD1F
+ezgWWbYHQ2FrAQPt9/K10jjmdOvA2Mbu8CeglWISTJiZnVC4I3IzPxxN76mauaNaXZ4Hm/vFkbb
nRMkaxa1Gauf63a2g46EKo+UeC+xNrsqxqztvp9gcFrjWM1/Mb+N9Y4nk3cTIljnsyZ8F+BRpxNq
or88NMBthg+MywyAAbtnz4QeVP6wK7BOSPFPfmgZyU4WPfHSxf9Z4yAtSht0m/pVcJxK2Xd+2tXp
5uO2CuLcK+gEYxzmsvWqOGkRNB/f8FxeUhCdnqGB0ojh5R0UykDpzIYuAb6R903SnidZ3mUdVr6g
hLKbkyClt4LaJbqPbHnuIUcbsWiojX6ioeJ7Du3HZg9O/kyTaLsKpLVq6hXOAcpbeEgI79VwdjOe
mndAhrSUbsYq7EANeZHQDgjWya0tHgylNlx4vU+6KLmoXeZVJczP4/+mcplFUfI0a0PStsqanVal
1TUFV33kz7VuIIUYgKJUvLCVzb4PiQ0sxB+zdPiwT42NzV0aNanmTcV+m+3KU/HZdJmV9aO2MFJ5
xQG1HiGRV0sLsxCjCESkg5V7R7Qrj3GuCQuM8NYReGFHXE2rVxlqzhH/NqzuRSj6UFaMZWgf0IpC
mWrvULCQ6e5mj78ySq7E7omWbGBx+J9s7QcOImZEULLoen4HC/O9UzYEFnFbEPsJsdhIexU+EGGd
LQyCMdiux52Jcuo9BSOeNraxmCcMKVcdRbJRGueFjCLeH2dkYZuasuH7mhVNV+xBBybml3jpoYrK
93w0ZkaavjtK6632Uy95ZdmhZIf4KwqQAmLs+dL45M/+NHB/2ZuwBe5yU8BfxMigcwMSn7GxAQU/
2fNcpjVPg55De/klh88FXPUMw0WlmxL7VrIrEyDbbtehN2kR+gJxu33DZjpy8/EvmmHQs0ZTExu7
dFTKMnhIvbNY4UEoKNTC+6llI3d78nXMnJLyOC/Jd5XrXVSMUvJkhsiJ9fDZYyRYaGwL7OeS/5gv
V0z5CwT0WaUty3BhO1G9lIHjs5HDr4W8vByPBvDvDs2EjYdQRlWYK3jUA+9AHx2nMGdzHcyj+Yyp
nQiTCc5Uo8uveTi5HH0p21McctNm10ZjbM+YEVPTzx40q+LDRuTbFyIiRbVmryWxppxsT7GttfMa
g3WycUneEDyzJsFkxQbe3kbcHAqTb/12LoJ9ioqtybbrnqWVFjsj/NhCBNQr5lCMiw9bxGT8Mz4S
9BEUMZvKndMtjkmaJ+YHu3BcYBkU7aGwhNYYMlVSDaInlngUGrj4E3htyj/9dfeQRWwnHHek4m5e
jDaLz7cJF9XZgGDPpM6UckMZTsWTwNWWfv2Kky57Pv1gUjoCFZUFUIvvb5TLIBb/yJ73Ug6yQBMp
PiPzczzkSI+Jsk0499F3yLJTIi4pUQRbcYr1oV/CCR53jrFqkhhVwuBtY7UjbkTF8+kaPGATqmJv
pWSv29WgfFvc5ZbLBhwiV5+CWrLnmUzGcWbiqG214Ja+zdJGV+hwS1FtlJS5h/e5VmpZvXsdsrFX
OOdDw6GDc0QwcvU0hLv0p/4CbQTpgSmspCKJtJjuAG4T12I3yC6Tgmcfqgfsr0JgTqmYKRug7Y2f
FAHxItXJMLiC+146XNNNmJ66cmyyviFtp1SDoMZ3rzf8KrfLdjdvWjhHNmXhdru26hW3q9ocNbuj
I9dq4MROFfFIoQEGs9yJIwt2N8pcotwcbx1+ivH6Qvqf4OAnFlp2mw6BLs/3l/mkjgEVk2XilrSi
LFacPs28QmM2lcZCYTAXrIt5ox09VKGs5XRZTkBWs2z2+bC5XhWz31Wi4VE2hG88ajECGMLo/C5e
qcbuBgKwMqtOESLovALcGWN9TY8s0z5Dnj0/dkaIa8WBHrcFdb/KB+cdHj0Lh0BkA0hNmHoIjMBi
iWG17xRGrmujVV+64ZurM7nkGRB2GvK54JofQ7J9Mq+Ht39KuH5QA0qiNzrTQU/WeZOdE+Plf/jr
7sMyYiFVLrwlTgi7EpUzSmv6gDaXcGo02gnBM0Yw3YwIi40iu/MSGNn0B8Gk76+DIzWfdwJxje6o
jR0zmO5FqYIWDQgL9Mzsj4Vn86+IBpeZzE4rnNtfteZ0NAsJEy0xExHG0pMkoEPUxCIE+J7uZ1Qo
6oU3AaetTsNXF2urN+CW4AU3zOQlcW95GrmGQS/00m0B9FRdnjZNyB7/dh6Ia5Bpw+l11Tp7eB10
1Xva//QmNKK+I9VgoyLaMGho3nT6Cg45OQ03ORut9ZZutuP2Pu6ZCgq47WGtrEo5AB6KulnoABst
ZkfAacS9HywKYTQNVQfomS7rQfrwIONPDAkZ7ufVU5sRF1ZBZEZfx0EQUAKJmDc6xnsYl5gGbN3v
JHUDhz6Ow/D7aOAh1AOSi3BWmL1Z3K1HhfcaUHtzmJ6TtjU1x824KSO/SN6xuSZ+034b/DuBkFWq
FL+QwhuHm3jhwqEVJWABqt/+YX+FMEjpfRfKlJXJ37cvx5oTqq5UMYNX+dHOs8lqhz/lUJcXTC2T
cTu7IwARbCYqc3r6jRRKrd7uXmKUtho9DXNmn3fBmiqsVok/efvX/PWdSIjB4biDnLrPfq9ztQ0G
791pUipMYWv8JKGj1srd5RwJI8V9u9a7HygzgQ7aML2nq+WKalHTVdWNESOyTMa0NV4cdvwDVljB
+97uJAkrBJuqJldXb8mEP/pjHdlPB3Bjgq7PNhcBIdFurzivbX/SvIG8kfgC9l0Suuqu1Y4EAw+0
DhguAk//nukL9SCvsCiJZuXzaK6WFIQOFiOzXXdd5YFLzEYgSzjYIKogFtz4kEZc9tGi7ylohBnb
GjroMyWpUzsaPF0w4+PY9xePdiMc1a9dExvFZWhk8euMEqujB6Ment+KTRRO1N+897Q9RpDqkWyc
O8x4+CifqkExW4ZahBDt33bRZotahhzKj3fvuu10ecR/ZnLPJacOKf7v/uax24WrEpu0ZM4XYlAb
cg2fT4FhktIKe2wkFvuYDvXsOdyHsRLr+tuojFHaZmxVidhPWiepzkciPUT5SRG0qwDcKRINF8jk
/5ZvoJ9tuRgtO4FR/Y0DfeqkBpPfUKTeuUqzo3Cm8TvsWMM7LLsOHYd5e6BqgxmPvPU1LbNMoA8x
FeEurFk+JtwGiIpOnVmpNHoEXJFgCkFfGXBu4Hxn0L6tAJCmP25DmKV5D0IjrL4eC3rPuqhfxDd8
nsh4IVfW+OHnHY/ywcuUuGsAaUBGtdsqMP3jNXLz7/pVJ2qnAHeMuAKMKQJLda26x3ec90+CEUD6
PhkgJ5TsL4PQbnLZ6e3dkxFKv/8z1EQ+nbdlxkq/O43jI2nVOoUzh2MP8HvEFq+X9RurZxemSuGc
yNzX9KBWdPQLlAYEA6dJgtI0jQqLHzFJDnf0SvkUtICoB9qbPRKGLYfvRqCbzToc0QjAIkoUGswI
MN0o47l7IFvxcZL3TMek5qXg5fnfgStxToMoDT/MQxkxgfpkPcdPyODP3slDZDgPSWIng8Iw1/hP
RtnOcsnLRkWoDbkzOWxNO8n9EdVMisG/50NfJm+vLj52rtdOkXSxyCzmcSyY3wJeKDGjDu08vwIn
h8HcEJelqA+WuXHCfDZsUA2lGYdMREYJnFJ0BdfW/Ab6Yg72RIiqmzUvsILEzE3m3fuGB41DRkZ6
vGznb0z0maOHv4qTzTSuS8lq1By68eZ2s7gGD+ez5VxzSFRaZTqzh5Yk1/zqegi1qPBWOGa0+9K9
v9J5+1CvzUL8MwzBibl9rk0tm+Wzmxb4xNRd6z5dZuW/U/2QWMi+715qO1GaGDvpRvWiQ/Ui/OMj
2zy8F+8XTlLhsaYuVh7hqqa6rprn+VYLCWo2opYaekdfcth3fLP53gijqGfdcKMZ5riUwnN5igkE
j8V2L8mEdN6p6hmcmtHr9ToM7tqWWfT9I9sxlXobfoa93rxfyU5phUwzysestBKNW2yLk5MpJvFb
Rc3tLTPDIvAlOn1j5Map/NFTrZxSYsTG+Rdeiu6lYHvtp9eJeTSeZf3WzzHcR/eE4ozqsFts/N5X
Hp0R+V9nKcyEnC1nD0+aonOg9KnSy9v16nP8Rr11Umk7PYAc/7OBmnlB18A2H34Crklw65gw4GL8
Q5yXVEM2lP76TyhkFNBra/91czPMx9EmUzEbhXXu2mVgTZGYouUajxKf52r8tfdi6NipPBBZIPtl
YFr2iq4XXEsDye6ZuCU0VtCidwzQWIZvV3bDVsiDT6LpEy/0CQMR+QS9H3rhdEJs53PdNmk6L9F7
4CSSP5ko5M6PbeXMBbmZK7qYolVcLFHDMHUpxL1tt9L8O2GLigdphUZ+BM7vZhx1ulRngWvQVwu0
3vYOiAWX0M9K103Ov2ZjOlwATWfk0YdOKZtaIO0XTT0QTMp264NsJi3BF+VWRrnjOVwVSbAYsVP+
tYwLvH4oSnARkR+537FaBsokDl5suFCl06cYdD9gL0Id4b82ApLOrs70g6lOYT1PE8FoIjuMtK2F
K322+FQcqLWXSQi0n7UDGeGQJNOKvPhAhHlTm5jBESbkg8RMaR7kzsQbG4nXroOV4s6Jr7T9jiqp
pVDwzPKwVYLUWIulEk1wkfGwaOZZPjoC0Y+L4oLUx+vcwyAVwuRdYZF85cHc6KKL8HoQCi9R67vv
9gCiH3AivH5s+pl3DwK9XchxV1YgwE6VUPZbaC/3uWIQ5ReM5ilXlC/jO/RmilUTZMz3kL6Y0RJV
zafGr3HxDLtGxev/tROGHsm7jFlvLI8XSJ+vG8+cWmL5vICBOUMguQ1HelntsbSGqvqvo/94MW6O
taBNvQKMqFX7QSNHOuLXU9i+J9d0XIYxWs07vTMwql+OEL/Qm1mBIgIt930qedwYlbXOFQQYuGyl
WB6TnIZvLDwUqN/6EX0ebRwSvGCdwbV2jCRTti1a1iY+NQ/ISr1oVAqO4qnCB5JHtYUJlR4Zuziz
WqTFQjETuWaFiQZ9CI96jyN32uytyPRHoBV/ISK/9jnJ6jV6HU1lLcMhjinJub/yr4kOk9RZ+E2W
UW7gYDU5mzrnehAQfnjvY2mkZdY5W011GGWkABmqsoTbqVqTPcmFULbe2GtHOHRtoBhgDQsawg3+
9ZWKAxGsz5Z8OD85m4h/oyDPV76vYLn8qb92PsbHklFppLyHJTr2z8JiD+sC1hec+RBaZrkyWmb9
J9sekIb3LXNqrcM6y9VMsKnxQFCpR3M1J1Kf1SnirM9bm2BkFKTLq18o6qPHRlfOxLl+TOVXc393
7+HXBqCEkEtqFGmgt0c0iPeX4ByzDya1ya/5VqtaEWY+cLFT6BKj9Yu0T1N6vIxdxpxKoAdy12pm
GdlIQq7H/x3Z3KC1dhJpXhDoMKpkdGsbL8whKY2VcN4eKgSTiwXf9caEuuoDJGP7LGUu71d0OX0X
jLFEN3r1dMF0uD/wk71gLmmcTZLPvn3GZ35t4LBl6V02rjyAviowAgjq47z1H8TmvPBgQ5GdYbI+
NZNeOX2lZeKmPEx0fZVR6LTj0By+jN6X+pMygAJJcTLeEXH3hBo6gm176+X/9r9ZcjWMp7f9hnj9
IYrHQ5SNJvmR+bepMAK5cXUFyrS8y5dRH+EwTaisZyXfCXuafF2TEuseSMz2xV7Af3HgiYeM36qg
qsGWaRm70WtlH9WZZapuBQ9XrRJmymvv+AXwr2KvnoTnww+1hicC7ixQH1/ElLkq1O/FoDssbp5n
Djht/tIqHNmZi6ebj/YSpjeu3mQel1DND0cvgCF3CrluCntFfUFQGCmmmY5v4aakf7zPJHZy+LvC
5DnumenZP6PhtC2rNKmvel2KBbgV4R0JYKsXwUKC3CDFbz+CKJBuHApqiXtlfXf4pWitO5Z9CsEE
D6zSt04zSdzipCONROBOi7p/+NZlp943FopAxkmBl/9J0fnD9aN8kEIAfdBCdhc+/3SGbMQUrXu4
kr9WD1c+nrSf2sHkVVdxtAxhWhP7yGSWCwKlGDL/v6Awmy8opZwORegteOqMSfd7ccR4ZcFp4ifc
5B5DBomRMwQEAmwNJHgGUYTw3h4Zeh942+1dEkA+VRMEtam57a+6JciNdYZ6wEeYt23CsQLDbLoN
mr5TJgdJk3ZmsISgpHM6ZEX6ATlbnrY8bBDIoUoMRTh5AS6Nrm56tSLayEduhQQfz5pg4Ls44cL/
4y2dNJZtYfAYaMxabfyKbmBaXR+xebdD0g8nRuZp4PSAOtOWU8EkIT7vC8wUkp+N4rsCI6rzrXTn
CFsA8P6AkoMh5S+t9rEGVcX8ga02xCLHP9oDnIKN15hBltrmiPzmsmcw2b1hf4lGWYjqByPjWlmD
VIB2MvrlLvigw/gwmBAhVm2oER2bp2LkRmy/ZsyL1oPVmkhubui/Vc6aPCQqEF2VFQBbwMgks8Md
g7Tq8kIa/Q5IkOK00RGNtPHGIjP9/sfnkFLdZ80je6/bAOy0LtqZww2e26jv+3VcUJkzKUhjneG0
ifrOy6Ji7R1ym6uqOt88zCT78bx9J/dtloO0yCUaLMDlQw9SHZINfhF1Bsopf+k7PoKTVl5/J0i7
Uh/6+tMkq1yn0EYkwFTT3MFfqRe0Y0mQMU24lCiYMiJrhaPaOFIWw81BoV/TAx6e1ju11StfY7QK
AaezySfd7HScVP2FltPfnweAT0C+vWZ8CnGlb7CgBqDfAUZ1MVHGaVAO/1R7CcAzzfLMss3qA1Z3
/XdqRVgFs2r4i/l8VD3Q2DGwq6oQJQnGGMx35OiioZUsiS+PvFo2/A7NhW/013K6MhMr/crT68zg
2yZyT+bacIQTWEbkY2YZavCJAsddlXLUqL+vuSTH7xe/hbjYKV+Mywx8CfYhRxLkq2NZEg6LNgcI
UxVA1yPcOJ/A6v6kc5zWVPV1oTKdinxzhL/+9oi2Tr5q91Cjl9ZJFR5Dp0o9g5/SUOyjrVczaXsz
sqP5yBrHx8nkpDcphfhy7M5y8+apJFhyjEPtdsEz3XgYFBKKATEVsXdr6VYFDYKHJaY+xcIssQgW
VAnJ6g6SU22Ss6sTtIirhVdfrvcf3w+W0Xu/Y9g9DeLeZeHym/Lh123q0HzSzqUj3hj35wYFa87H
CL9Ns9UfIRil82loHWprtXZq8A/uqHe52I4nvuATSToZX3gjJzzBsN/4EAsGAUm8XmWI6NmrCjs/
u7BFF3eGkcKrLWBYuMjRIkkEfIOpcEezesFNZ0JN7+J36IhwPNd2UBPb/sWkusEa49WUS90FwJKa
zqnXnCCrlUWaN/m7T4SqRxNXzjT+cJ6GvIvU8XCskEApGk9sGL6TzblHdBF8rme+vz1oCERaxHF9
5zZ/D+OXnc6tSgpqBDEWRlbRR7oGTPDdgc68nOxjmTpWUaLN2d2S2hpZ7r9mPxvzATzlCIawj0CB
kB6f4pIkR40lK+lBIkeIBZZdDzfJtHvlT3/0M03u4mJ0uK+XY3klZx/UNWk1p4N+dMOj2+r+oTT+
maxT/1/S+lBelAc+tAyW2yK/Y3kvjmNv0/R6CZG9SysN7w5yRsXuo8OP2n+s19zl71u38SYv7rwP
dmIOWcArNzQhSnZc4BHiE8yPhnca6r+XTxc3VeFUjQFghhyIyIpbPYE/VPf233iEs3Zm15EMg7yu
MGYdUdCETLQOb9ytEgNeKIq4i5RG6RkTXog6jQAWcnF/r95S3RmbA+GwMX7bRuBhHf91fmLd4G6p
4hpTNvMtB9FkxTD2bA+eFR8R++8XMf16JjEEBbbTTuyej/1VcvaYkG1QYiuWMqAQU+8ja0pc9M+d
jrgcGWMK0wu7MOQa9R7J8A0kIIpZplQie9jeYnTu2BfYSLPawBWZWjqsGUXsMONjjAD1UrIa0G6V
8xZAyUnFNnjPbNUTWxslkhqG1cO2Ly99j90alDxFTcehfpaecNRtqH3sOHAdZOfv2BRiWeUN6HPM
a5fsZUP1FivF5PcLRVvo4pr+aa41ZMTjsYxpcsVvcIYdMcHhrFN+8i8XyN2Oq7817QqsB0oPpuNf
udWsLBv5jqgL4iCtXLuRYwx5prAmSbD2E5mhnY0So1zmsWPBtsT17S7FvVlTZ+YSBv9h9LuXOzEf
vPPjsLmlPUr7PvqRnOXPvz5ps6NEoUCLpzANP5sAXITjNfkm4hBAtg2uHEDN4360GQ1Kq/linZ5q
OHUPves0LAMj+DwCYRd15cum6mtXfLTxaUmdXZ+BphWhST8nFzDsKeRKDnOa2iDvApK+SuT4NI+A
3Sh9+t3hxTvG0tLJdqY5eXdBWWQk22Z0f9tal9Tnz5sbLGxg98ZPYaSCtOG/rsRst6I842U67uMK
x7ML7iiKGIRTFMzaL6YttYkSvAvP4JKdmxT1hVDUYCXNkyANzHOWIdQlZNClfeeO+tYu8tn/QVSu
zZ5AdqZ7lIBXHBFtgXl5O+VllVv76Ra+y0QrxSZbZY+AlODt4E1bD3Q9Fl2OI4nNMaa7pd/+1piU
3ibHBaeYLCwkpnJ+b4GFEZZJM+kMnFVJm/1Yz1u1gK6R4CYPDcBket7mX7MVCFVw2CUl+t8Vyw/V
T8rlFoLo3bc9HGetk6Wb0z4F7ioH8gyKLblpT8Kzti1Onk2cRrDvuP/7a+pZLuQVO2F6tCwilXtV
e+OD3aHfUD1RBJ2pJdGCHfNSCZ1Ibt+3O5OBlk0KWcMVJIav7P7/bLS2j+5ETrC6bvB9RYJjs7Sr
6REY/dzzCP62dSeEZ9Y5DRwJ3Z/iQdJZQ3QfFITuqDnU1zT6BUO72KIDogCQV+Y1WBr8y7gpp/Lj
3ndn+wcS+G8ehqT6POkYSFALv1ka4hE9ZYegXbE5Gwq9Uw3A8I5UI+QmM7YkaPUCMwqeyIUL+9rX
XRT39BehjcTUOLIaajQzZ/R60spem5InVRyh2woqAXm0xdBIb6SL5ARM9XyCNrWj4DWYYl6bBP00
F9+Gvx8EYXkbobbDKFH2CHmOSqAwu7vHdmXiAfqO3XH/T3ErhXlAoRxLi1gJIigQBabHgRX86XpO
6QGISZDzOGke/6V6w5HMRjvztKfZWQq0g4JCGSha8cykjNO/Z52xu3GFmivcu1D+KLwHpBu/xEaL
Y7WEk+OU2sZNxKgnoTVwG6uevwb99gn5Slnr9o+aB9XcFyiPD0vF2cHHEWTggO+ZhWfYACdztlTI
JI3cHPghUwDbvNltrx18UhDvmgpdRyeGuoXwxyCE8QKq6NEcvdFiNp3hCM+WZy+ibB/CIbX9eQd+
IbprEPyHqGk69n0CVEVLyajmXma4vK9oJulLb8fYcd5UqghPy9gRRjFC3U2mYf05SKCChUKoOUTI
mX76IfZNtO2vtmAINxF8bWxNVo6RkvSdVGfGWSkUlwN/vF3Rmq7WzKXboR9UvD/yu+o5muWi3xG1
HLyiwYvJ9M0yUdOaeffF1blvBdw1mBaqUBFKLxUW07EMaIqL4OqKNigPABuZt28GEiDZ3l6rPJ5A
yY8FIn4Nt5+05pmwjeLNauuI54vRl+U2k8h3dUU9wWDNFFB83fSHRyCkac6mFvSD9pSPvMP9ZRQq
y4IziCerd1HU2Rz5KIF0SpEV1aev4uTLYOl0D28GxrJP5JTmPkclrbXlmc41VzY/BrJcjboA47xq
JIfkhtQAPoQhX04znhSp5xG23DycozRmy1YtmD/E8rJWUUrLwSaPbCecFRcLJtKjaxI6H950NfmS
hNS7UT9dvrP9qc3EWHBxrhn4xcCPz2wVRFCnJ0VaMfcZOeuq2RXrVSenG+HT8fPAIQjtXLCEv2TM
+alUTDW3NoRV97Gpi8YqTLtxWaYZvpMMdW50YTjxajB79y69U2XpBqUyME4kqYgPRNHyBROM4PiJ
8zzYqVdIbRRBFZeI64bl1TAKTFDtSbL6KUwvSBCqt3qmMetM0xK7+ExPWJQhKJdUpipgtx0tuyi+
IshJ5NXeWQsaVx7hLnkWJ3N0xQZDPTXqUdoX7uoRMPksAZlgrt+Bv77JXpB2KYjTCe7VoQmdJoff
IZhxHxdsdkbVGQaVDnJ67Es+4OOlF6kFBQ/cMyg1fN+mjzEaC5rtLDt91fWXh9lw8XrDr8gkGQmL
1okyhQZTjNq/PR7eHfEAxF3F44v2+fXYrG8DJLa0Py0y+tLltRFEbtsGdIYRbp6looBFB4K4LfOe
w6JAntUhG83kgVCSHvP5XkyGnw1VFwFYpZm7zSVoxw9CI1yHLyMOUtX5yZCD5OYqbSI101auavY1
vwfYbz+h6MZ+N3pQKLOeo+pO83E3enFGgCe6sHcaYL7b21NHwneioWBzLkztrmNihm5XQO2mFwiz
Bij03UyDXh0R/1XLwyTMt8xmmcQ+BZ//wDZiZCF0c8HD1HJGOLXpiV5Ey3F9TNvtj/bGVk+AkEs/
qbZt2OgBGPCuEs2XEeLAcDoKgBZWbEkKF8pshdOlw6OYhU/PL14Xz89ygY7D3EZI43WHdAYP8SDn
/Zc5Mm/g4/2eCVDYBOrfJpovOiu94G3BHszwWfErPFauNOEja8kepbt3NKPwb9gwQ6yMuptnuDVx
M1JQaC+dyfxdR2KyFdOmDWDHhKyW4AIHWCy30WeYwFwh92xEuaYQ7T5bTvgipyNfll70Eey+7qcE
baJdNdstI4bF6ZERiVPQdAVV9zib/MWAEQSWK769JHaW4sdUnKd+zLGEWVhDxPOTdrPOXHs4QqnH
iompGA/77YfIqNwEXgAEZYQMi06+uVmCSJkQ1aIY9Myd48dPNv0QU3cJjDXDX4PiY0iXmaFY8qJT
kaBLc0Mq7ECnEf3NdiwUudYZQXXrNDSksLU5v9XdzFnDsH7iZVt2jh3QhjzlFtP+um42pu9eJeUJ
d6Na7gGJ6b2ICMOtV6CGbcjX8vXgqaQG7xbwcPpp0CGoOVNhICfClO/+PGp92FXDA6tcYk4WXfUq
9y4F/4c9Qv+ykTn3vaIuT8HLR37e45vLCPt8921ht0d50bKx1+W2qiyPbyiOOJ4KCR+3xyfP4DrC
dxQEQyCMsPOrJj9WVbv5BxGO3zt+cCaUdk6Sj+ek94FDditHy4Ey08WfjjLEfQ64QAMaaETa1dmu
/laP5uK37pFKi0n4a6ePQrlxzvEDQRqDUJktTtoBdGkl1xNIQ+9CS8jNjSDZZSYGjlefb5PMNd8a
j0YG8zp5OFOeRKKH2HRsRmvGocPjnhjppwAd+DBY5Y0/1hoFk4vHZNAPJBMcN2to06K9b8ujnkgY
UM+BVUvuP9wbCBpvSm/5J5y5ivWWBr0dxj7Is45UarynNO5PmzJtkHlt9iLH4ESkaksrRz9OafhU
yYEeDCVFxyUEwmiqZfys9haRlcnWI4/LafCaEJ1FmOlNS7KKcBJ82Lx7JCFT2TZxf76GuRC4c9YK
0AGZWfeBFMfGOyzoi32u1dEyTwm2cgXpaVYJsMlR8HdcfiWC6jiG1EFitaKJxAIc+uCnwtyLa9g3
mlmdwMoFdpy9cwTUGwT0zdk5Kx73pvuWrFmJi/hApAP/vT57hh7pmC27cXFGG0jEztIcYSPkK3Ob
JDDZIUw+u8e77D4QfDq5EOa3hHnsafpYJWO7+bn+dODAH14ZlySwtid7QdhSYqamKooUD/wIPChB
3lxMAOOIvLCKFddcbhxYO9AiM9faOqD/9bDG9SUA97GSD2/UB6UZ+cr75xZsq5pr8usGuuUtMLmq
ydumHhfmG8GsYyO2umskd31hHGvdDV5MJeauAXhTPsWqa561Y3sTb12Hdecv/aTOVxlbS7WMBOye
iIdVhMpcMvmVda+T4sEWovXxgA054nTF9d+fAR09VMuhdeuEcf7kwaW106n0DrHnnVBfaXh5YCNU
/eNmbB/DOWFcZxrAf/MFmox8VMyw4kOBbU3SPnvMRkqjBC+S7meV1KHApASHSB/kVm9wmvLIXiHu
tiAkjBZqLTVwVHXCwOWFsWlY93MjWrdCfKq3CI69qDFs38gn/VflsgiHvlIU1JrSoZDZP9AMP+Z/
5d4YrP4eOVK067sZO3Xf1te7Ndb7QagxK7/NaTgb/pWEuSZrqEKiPSmNnGiKy50V1IAyhMj1OPfE
OAWEfi+3FstneWhBXwq1t5cSbEVELLTEV+zhBIJe4kvBp8K2+i0ticipS+v+yNZGITeOEz9uaADX
UpJByVoE1fAGUTiUi1dgnRyZI+/GC9y8hbmTp5WKKWdcB9nGr6L0FogQEuwI03BVHGuGy7bJ2yT8
3Jrd+u2E7+TWW16Pio2TG8BKO/LCGRWiOuQe/ebez1ojahyJbJhDD8tHh57JtNL5p9wSIoKCx9g+
lTlYNWoMRn+pizMiuiYYUqoi71LxO1V8KyEORJeOtjqVRUwOB2jw5LJ9Oj19b4M564TuFuAuzd2h
ARaA0s98/dMYX8A/E+3U6RfGTuYcrIi5xd9drsY5w6+82P+yO/vceGE26BeBqAaslWjgD4Maf27d
3YrCqSZMmio0UFXs8YoTCYIWlPehFzY/JDs9CFfDcqjsaWYvsGPPNo/TY4n1E0OjSJTdlzRrn8DT
LXZOuGV7Y1VRslyXQDo8qcD3oimWBoHWxGj8p0fAv6ubQpSx9Kl00CsOMpg+Vm95q3vdlzKtIRJ7
QBjZsEHquCSvv+vPI3Tuxb073vFFr4T+Zig17rZZWPbd2VmaEhhExuqOLW3JdPnXd9Mekw13DQso
/tfdtP0eHXMLrvJVHzMzf1ZiIKj7Un7YMaPIbc2rtdleH2MTXS+NzIEsGLu+dhbaDpg2FGgEyrqP
ReR0isE+iCs5bqQJkh6O9IR0hhLpA8Kle5MUHFpNSTAStBK9Q0xPGgFeF3m6X5exkaCmfzP8o9lH
Rww+llTuPdJRFcijcnTpn7LiA9aFquz99mLjm+NPFy0+12cX4cGPhrXSg3ePd4jBK6rCrG7QCUcc
xVeeuW2wHKL5VEDOhYrYOYa8YX5Wo9oOhblJUxJRe8MLS+w/aG7jJ2jkesxH76XrvPZ6ovF4ze8n
xnkUbV8Eo6CmgNkocLwkMrfM4S6ZQGaF5ZAQtWLjHdQSAbSb8OAgoEBN1ERWVI/hUsQeEAl/9YQ9
ymwQM35B4Yds5C6ohw1qxcTjBhjJ75t83JuDpNRxzqKpAa33S7ux6nn8LtPR2eHpLpewLQmx6MM/
wBfu2/fUEPd04I/OjTyELvuvC1G5A4mS5chCuWTLT4jgF0s2+UHh2RPMZuGRf1UggO9zdkP2HD5m
cGW4pMBpj8n0RfXhh9YjRIUNxNFjjbm6E9lIlF0jR0OT8sme/noiuYopeXSR230auwwDAqoU6pF6
uAT3WdjwyEw/MLzszI60AhVmjEkHfG8Yo5PNm7L+Zm0kAVL6YbB6dKJKKhBZz2cAao23Q4w4sWkz
aVjevNs69OD1i4TvgJ9YrXASgfrc2rx2gmeruq6NYcfSH18x/FmycvEY3mryqGjLUpZHdfnFNcKF
O1rkgpxJ4ZYzmJDUmU5amhDoq4KkHtcCRMyLwXTuTA23f/6oJ4s1ygKEFogm0OjT7AmJwE0btOj1
lcdxupymV4lwhzOe9tkdjtVeEzIt+m2nuXq3A66C4MkXOwMwgGh9GpbeWUAu5vkJEG1h1yXIuQF6
0cDFKU5i7eysMmPfVUBoKeZHSGimjLLoQoT6E2i18aMKx9d4SZdtyAtNDH2RsSFriA50GP4z8gT9
o+6qlAOVGsqQHAdjWtPwjidUv0hWrVLY8IZCBYBUH0ELhJO9SNRi0Uc2Ykd/BU8RkheVIYHi2/EI
HfMhFUHZoa3gTDqSJAGNVIb9tBgr8t49shiOH+mn9N+4hv71l+FQhlrk6gFEhP03FhoWkdr/bClK
fRAjbxZHPoAoHaIPT0Wnv4ROvBCwIKKb1gpjKt/hPMl5hOfwghI6i4JstYcVc+4W05pMTrgBD7V8
JnAf8csGnncoQY086kNQdYJE1MsFu69IVO69dyp0VRjOIvOp+Q4Hvz6n1hUn2ZNPBKik3TRae00t
NLMjaJNX9cjwuYGOiiD34L8uDpC0ShmbLXGrbIVdCPxpmdSrCGbPQ60M81U4u5+0BIXJsUL8P3p7
Pub3u5hSxitmtMyY8aZxAxwo46kYrXhXRWokT+3PgtgXDED6IB3dg4mQ36UrWKH0ohuRy6E7slr8
wIo08OKBT78q1Y36wgcBmx3gZQOJmgSBPhoaKHOLGeDq5Y7I7XCivXpXfqgMiqmt/P9JH2Hahe+l
EY6NhmcwVIS5crDflitdnt/hHimAGyWOWOAu+x7gvkuLhWnwchT6VLxqSLX0zzVWu6FrygxgDcoI
t2arqpUAp3rcCYYWW9qqFzRI4SMYsGbcG5Ve67yhIe4oO5gm33OBytPsS9bkOcLrUgaSmMa3zYm+
L1DzN3rMFuX/6DM47I27jx5vyMcosccS8dW44qCt32Be0fOuL3FyFsbbkBY6JKyDhPDEe12Wi7oX
daJEDmtIOC0elcmnz2pFGGsd23NQBcen2OOKdXDX3vzDEQCe5suUbuW6AmwLEjQJJaszQ3tQ91sq
03EV5t5PTkgi5jJkEodpTqmk6hZh1uooHM1OQD+jgKfAs1RSWLuiH2kI2SvKkQb2IViE4mPkTGQr
eVZeyfv2k6V8iKd2V/Vxog+V1Ba9K90X+mVNXLudIiikTFeJguZxVj6b/PC+Peeeh/zwDo0hGa0l
Pd/OtvCEq/Lt9TAxzFC98OA9xQwB2kXotNCREEJEAKIhadH+PRzg1CIXL0cBlxycigAQMTmhItOt
koRnwtq64BM5Fl/lLK3GKM/PEvQACUPfpN6Kd57B82iwKAKol/uFxVW+FxmvT2iVjgqFgroLFqNJ
oG86ZSfOGbnr0K9Ib3wd9VHTTuQwtqaPlkJxyY5kiOzbI3GBVsSQdbKKYGjB1Pj2ob378Bz3gxR3
dSwEaSd/Fn3lig0opGhkzwBVlNY+g15WKw971HCGVszkBfq4xljPlslbH3HL1Oe8B0MGNlJCfAfj
gDRmRfEMuoMPBFHhNcOq9EfaPaLay2EnQWdC8vHbU0alTsZTKf4rNYBSY1deBDjr/9RLsvYnmptW
A9zYxxyhRAKBvEiQOIDuNN62dggrEuqx6kJ3nXNdVL+1UcwPpW+IgmeMdKCVBsxzt2gWL9rqh7cx
k8ziuWKrz1j0AoM87fO+nxoiX/BGFla4YkbmoIq2Wk4hAi/VNinz86qa4fu3VXu0vv337qlvSKAl
1U/hHL+lqCU+CsJqLlO3w7qTzegYjKYHUkYT6I4Po+zNbQeSRYTjXWDaR24mnp74qdU9ao85JFOS
PWGz+C2lGjdPK6mRPIibrF0qxPeu9fvkHr9uBvSGOh8dB9FEshdUsRMMIk9SeXvvTgfdZrKxl8y6
nwnTl8CCfBbnYCbGOoia71SPVZsoXGjxjL93l9Pa0hfbHAOukgbH6T6YLC6G9kUe29jRI8LSwRFA
x6kl534/wsCpisutsuTDggiXFwSoye8QJF5nZoV7gpPUuIfLWhToVsBTxk0/IPPaf/3FlCsRlPXO
KpLbnRE2WkH9uGAagyq0JO35zO4HmXWF9aq+uHoaNxzao5UNhoVtoEaqLQ9t7K/6TPsuqSynWXDW
bcuLB0iFBYgG79oMLJE/aN9zYvpkB/eGGeLzX9l4QA6DQ/M7kP9Nb0usn1fBMjki9mPaofcn2iLT
iT4eoCdC11hpsl+2nD/Ke6/qU+x01TETFHfiHOs65mtICRh7QOjpHHAXYYHDmv246lhaF0Jesa8H
wHGqCg52Jh0HfTUZe9jrSkPOP8clHVE7IiHsWaseuXgbPAAlCLJ9pdM6n6x89y+fv8C8JMTPunh9
kZfAn0C9Mjk1eFHlzz6dySGYZYmjrQJodJiE6CuI2aUz1xUBqla/lQYUOlWDeBXS26NowaZcuXAo
TqDLrQ6PBIP3uG8nuGawZQlyvozT9lqH+gO4fMHtjXKLhZAQHWdEbDjsX/t+F443ZteqzeCSA1ic
OzqapVDnBw+pi4YL3j/kasgmb59mXoW8lNNtfXnFOi33CVoVSwo9TZDblB8//aDoC9Zk8yzk1VSL
GPYrVtibMKIXxXGZWYTX96/4EPhEqj8Qd19gycAFY+1uWzyEloG5F45Sl2mMGFRI7EmmKtX5q3eC
QBHwvY9PFXQFJg4/LppJts3RbrS8smZ3kL8BPr1KjfKTtZBnVdaG/7dIgxuteS/GtbJZSL1kDFQP
GZmEAid7TyhQINFeCuJ9SxPWEyXfy32+V5ZesIpduTXPegfPUPr3v/DJqwqgQNXBzmr8nHGt68Ni
FOiiGJobe8MSpVAEQ/gnbnq50xRWcnbQGwy528Q1GoIb+aaZrBGJkD+WlGXziyRNmajDDLIAums2
1SYGuYj5rJIeTOhSoq23aURbPg1hBIwRX0lB1dNYKMUluLnJbyyS3khYqmE2LgEADsEg7OKWXpWr
KPhc4p1WMR7yQmHAzjmpoM+gq9Tgqm7xziIUZsusI/w8VMgU7UkjgTyJE7axg7vZ82TIMVChgQld
EqGtwqjXpz5LJXsKqAxuQRh23OzBsfQSWZ+jdgmC9VDmoRXP5nJUiHg7xSicjn1BoYpa3Ohy4gdj
+NaLLXI7GUqlLOQGDeB2M2qFS4WV2QoVLxIvPd7cQZlX+ugaSIbvP6YwAGY9m80A//sDcqzAdoyv
GsnHy2BR54zK5qV39LXfneRrMb7u6GCpt6kT5yTqWAFz7DW22bEaatejyFJQpnfVXdopsI0i0ZwY
Pt1Y01yTTW8xBIZondhZaufGbEOOtNxSOdCyvv6CTi5caSO6Nm9ifGojEGxvA9iIKezPSArPLvpP
gpssN5yxqVf4lME9K5UJAuIpW5K7sJhzyLPEQe9un/mnHolz0MQEmtzT5ew8NEfkSKNkkN6Otacc
Q+kdsu+kvttceY7aNaGBUARPI826PWSqPCfwR6tpvj3fgpAVh1UYx+OhI8unDJpoYUQhxQ7zIl+x
cv3hVjCozQpFeN7Ssh4xA5sjxz9mjy0cRaczI8QADuhWnn9bG3b+QF9n1JeydCIqkIegNQLcRirR
nKluU9wWN7yWuHbG1YC658fjtSZJqasLVjKVS1JwG1tznHdQY2hgiXs2/Ps8GsIIuQN8xO6RIQFK
kAorlnJilV2GP0M3yFgxrTwYOLEmbrYatoVthkU2rvRg8NAID0qC0fVCFkf9yrJy8yQNFRupFAVm
SV83dPF0Vk/v6SX+uTrDX9xY5VmsHjeBbZtuhrVsCGYVFdIkewEixwlo6GGa2IE0DgVRkwGsT1zg
oGPKbw8/7ujKBFgrOHq15KUlFFwDCMb/Xs2Ur1z7R8xHyi82WHHqmiEX89ikuXbRUmeKDXqo6vq0
l0thG1ffYCCiHUnTXoNYqvsQMJROdtZ4dXH0Ln14rUk6hlPJ2G38NPMUnGesZ62XhnMcuaUtQK1F
GSWRKEooAkl0ENa8yjVtzNL6NJ7GJzfyOX/u2QTRH5flFC08KGDsqYJA+B46wez/W9lLkcStU3xO
9oUQx1jzDpbr7dWNyMg4fUTFBDSod+5COPZ376KX8OD2MQgeNHubx+DAtgwcJ7IkTO6/fj/k2XV3
UUD2IXZ5CFaCB7BvQl6pI4Db7HzEBmROAruJF48m1yTq38u1Rs/IGanaaolKHbBN2nAjJiC/ALQn
w02GXFVrBnmXh3hKdo8WEMBQMPrZtdsVz56UztzxcDhqhQkHN0+aLCVNfQRihfeGws5pSfNxUEYV
bnQkxE72n87PhLyYXIAUHkrRTZ8d96SlBo7lkD9qjoW58hiX7vV3agW3EgZ60Bm9rx201gISbHGn
7vwEZk9UJQWHEr3mUoE1ujkOWvHi3TK116/nh110na8PgTuOX1n8gGY0IcSlYLheosJkdcpkwPW2
EmjSNDnnhY63TolZsvqcBbcpcEEAaJMcPFRa9Z3LCShtPXzp0KKbO/0II56HTKQxJL1iEWlNqPdN
1Bed+xqezJz3v+mqda0Vd0y5SCXJr5eN3vIuZbqnU+8kmqPpnGqVvAhjML0PFJQ9Z/TU5+4MBk5K
3iO/MJOreoX2XTsmSbA79OqPVZDd8WxyKGeprdA/i48qNcgAqJti7erU6UG1Bn8FNvX0og0RV2Sz
aKQXCtoNJzcb/A9hcs1avExlz6hUJnq2ZS2sOtE+pbl6n7y2sPtFUwy30CuQx93ItN4gjmjYp8qe
km8YTX6xE1HVpfwW4yTSQ+BhYKipJSQBOx1R/w8F99O0l8Kj10URlfLH4AfX8mAMKrHq8vDIyvFF
EUyhTpkUFb5VDpV/6BYOh0B5wc/M8Ay12j4p9Z2N6LmKpQbt/iiJof62jZwdLDsykRquSVA1jO3I
/lmcORHGQMs9G/7jK4O9UfMvaK91iDmP8FfoqVRRoq94oqRJ88e1aQcqkLMTzh6WonDaquwlndgy
xiV87w08lMLkeHYbgcPXl+TGzuhJenxNugZCkuyguxdI6v/6bcUG/dNczT0GDADNGTcJxnqLn0qq
6nqAIz5v8Vq9Xp9sjrwn3S7gOQxz9aKJRYxchqBxLOroltp2NEPsOIINz7XtbwPQZ2kPWWCBB/sD
l64WkG33Bc25j1sqruncrC7LZ7T6pOJnZCj/Yy6W1TuHYGtE7dmXx+6XuPBWUc79GACyi1wZl25W
KZi60aIkK1jkn6hNqRu4HCEG0sbmLV6aKg69zJts1NPWGWc983uKUaLKcukF1cVPV2JjaVoHiLxy
+3PE7zraOqsfd4/N+3ep6e2g4XGIy3O6e+P4UsFN0EhE3GNRXKXEOmv24uJqh/r9Lfrc7C4XPEMR
KiFLMvTh8cu5GXp+2lU4/9F9vTWXYa9AhBacqKQH0pO3a9KKEdT2WICW+ZQr4vpGjBHBVkXaaCSD
xKrnsCwxsqg9cMS+fwdbJXq+iatqGEPmMsv25F4jHOWLjEFBzgDlYvUdj0Fo83deaGz5KtUUiFJo
15v0GMOlB58q9n/cD1X8hhM4kxABhLmpL8irisRTFzOjF/7Cw15bXQ6fyQJ/Ti1vdjSj9F7X25yC
x3lRQTFbXYhEsbNV/nj9WRlT8R9w1VfiDMnikokdIOfXONZM2/65KgbiBMJhwHezFE/5avAvsdRe
ynLb8xaifJZ4QxsnTk/fu0Z+NYxRSfjXJlhoX5YAdHQuvDuCGxcjXGRRkcILmsi9cPPEFn6e2ugZ
kOFk3+BDqg2znTqR1f2TJBSlqDHhjeiUAaMlTFF5PD1YuRycp7b+xqkjwAWRgX0h4AhuzAS0UKMM
TnHroN4h6WofVZQCTRutdgH/79gTkMGKPwtOpcFsgOL8P52LUognSGj02lzg8TRwyRwEoWkVjE3r
cRLF/qRm5Ae+XBLBV7LXZOKLh+0jSp+/nwc4rvUv6KqFMKMvNXmv7DHComCSKAObcJvQvU3DBWcN
sBrmmHLU0DGs1oilmR2mJOkFXNE5vbl1M4AmL2+Pi58wJsQJbOVo6jIgyRHS2tewhrzK03WpxIDZ
fKT+XtBB2K13aqxqa54AFjLpxvLmjRxLztZdVJsA/TDvLHdKQtsKbiCXR+hp6lXghavW1FhjqhsS
+8WG9+SFEHuJ5Jn06KEKS8tVN7Wj1ElZKZ0y+rf+VHcOrfqJp6g9QZpo9Kn9OIChktCkCslJOl3G
ic0h1TXEsB3XQ/8cl0pPL4DaehY1oBytdnw0QK/rc/GUNL+Ap4zqTljIvjUXvSOn/VblRozPsUSd
Tai1arEcGEYB21LT4pCrGViHs13zROEeDqLbbK5Zx94zmHxsrOXzq474uwweo98Uf/uUCbvYJcw6
PDdL3d0QQIbUhVPhUmqGySl64Jmmzxd9J91fgKmf56A8pJY/yoRmJqf9Zr4wEqagoNNTVEebwEAv
D/2wqDwKZ/6vlXL0S5KOtXBk1a7peVs0YQwyxbMJMePMpGM12PSJ5J9aoIX/3IYbIAZ5RH8NApEE
LourVN9dH9I5lZgcyJVFSOmtivvcNUn1cYq/Y4wnPVrrvd/zKQwd7Li6dIrUpYEZImZGuDhMEHdH
0fogIWeRjcKTBHORCQbIkI/tY9cQCbqhWH8a9hBw0UjttZWoZ4UUb1OM9jKLNFhlIMGaCXyzKlfN
IkzlrqMbOkWn0DFyZm7R1ys2FPbEBgvQG9oPbaS3C9NR11Iap2GpMxaIhq8HafXALzcaoMZGv+L7
lqTlR3ErodimByC82QJVVlptYSuBboXOMwiRHTrMtFzhyP/m4iSP5GmnqSIjSnfXAm6PCueF3ui7
HKGir6GmVe+c0rh5F1Ej5yVfHfye7GeHqFK/Wta9m/uDA6sfSmKTCXKED50K86SBN9ix1V8V/sB/
sQWkfMUrdv4qcSwPSXXlQDpSFuaOTTogFwi/4slLDX6ZrDikFbKPUudE8T0iHouvexhLJ8079CZF
VeTugb2GeWrR5EC2JCmU/ZOIs1cF8z7G1RMK7ay3N7qs5r+QBe3Zrizz8/dAX6zf3vyevcWcaBHs
j48l4j7BlTJkdcr2Dy02UJrtaOL/pRPl1Ag6PHurALK+qBKU3aXOtNsC7khJjlJm2SFxgTDGrJRW
UNqA6vLtF5a2/Aw8Bslm5RQiNZxwEvmxW+xwF4nyLk7YEp8Q12Fp3juHEu/ZlNSBngD4Gh3lt9xN
nsTtVBrFfGlpSOU4qG8NuBJ5loaNHEt/MvnyiBR4/3xxCtZ/5fnTBq0+n197hxcChhqjVC0QnR9U
/c7beb7mBKDewiI/19uVeTTE/sMLYKk3CKgO7+V2mooauK51vRs++8VQTKL6Sg5U9xKD5+Jlesfj
PeoWWNt+G/rP/NEIA2GCjC7oGBLX3hFPe/zSmb7WBbV9aeVHlQC10p3pvEsTSbRbxvhAKxVtB24k
YlUloHjzjA7swmDdq68yoz4bUbP9cNSNVOo2fl/758dMf11wx5D8o1SDJcf83UbO9hrVWuw75wA5
++hzg3H9rQnIuD05qhQ/a73XvYiCPQMa7+VK7ApJdNVCye6mT/ckJLknm4Ed7bbCMTfqBDDgTbMl
Il+nCqf2NCQsTM/3n/7py8f4g5Qjg/3HqA79roFUKTf1L23c1lnSOggYiWHPgZSWiTY6tZ26d/TJ
ACGt2kdkAK4yg/s4aANC8ZOvAgYDv+YzE1wMc8JrNX2sw9x/YO8i35WIwlxydA1dDG1A5yKxHgoz
dS+IXuHYxhhWLunfsV1YPUHOQ2329dFM5TyBnHuaKITgpnyE7hXpUY+QefufDIsTbRsJzZuAFwn4
3damsoXxmhzmLND4n1+rd+sYAHYmxVp37uN9bjrZodWmgR6NUli/Rq5rSQTzM0lS0BQHcQ6Egumn
pTS5htx1Pu1Yd3n2mGoMnfvJq0dEdcWgOgwiH40yows2XXM8kvS71oqSAZLWR1r4YBLz+t5y9big
2lJy9ydkZRWoI/tcsSjjNqOvIDrQjCsMSwEeE597HSNGIHhxSnYg3JkU7f9C/wX+tJo1/5w1U4VR
GU9zBW/GkS5tQqHnIoaM295aTwuCMZibvY3wuCOxmS+jYtBRhLA0r9nKirfe+fcTO+Qn2pqbZVdG
VoDHIDxO/EONADoUlSMXmgMpsLOBNwIKqANfZvrwJu1woA2Nj4By7n4wa1l0R2acXF3v4BdBkCV8
wi9+c4qg8m/sVZqhSsLQxSSbPQQljHVG6/TPN2ErxpuBUWyjGAdysqbmTUi1qVB3ku8aUimNgwt+
mBEF5+nU8UDiFFgnblWqG0cMrAU2odBcwM/Ti7p4wL5jdmuSaH2g861PcrNHAVn+gIkrsRjXpaEs
SqF2rEVpgENdlFjFT7pNWop+r9wZ3T4fU/nYoBX4/wQnJqvrBHQaEX9ce1GiNKhROyqn/Ovv29f1
31RKohj3gCQ0dV6LLwddgRs/dB0z9YzsaNi+qrzUqwQKUqzVVxRz4CAREZ/RRXeeBI4T9Bs5K6SQ
oFUdM6kKl3WMF7RrW01Eb3lwuVrtGRQa+BNA80bRMzaIOVFmbAw7xOKjxbZmjUYK6dwbXhY5qxod
l7NrnKcevitOQhffO3YJWT5d3Lp7C1076T+mS7zB8Ng27MtlzAODH6GeWhoOdUcaHkvhnVAl0sLn
8l/wQRtBXdz4lMUxblAJ/tOr0920cZlbezMJzr3s7JkM70WGsbRhxdShFGp102/IX68wMVgVGKr6
kvWm4gS1XFDxp2pLNXBV4gve10Lif0Azuf6l8fGnia4cl1ftvZ0GuixxbWVSen4phkxrmNSUaH3Y
xmzmH5n/JXG/Tvg/bKLci/72kow7l6uWdEurs3yBRZBsfVF24GsBwtNY1bJcMp6tRgMKTTH8qeY9
zc9Xz30dToaCYYGoJwZxadPuARTzBS46CRxPclrMSCqfR/NdZQELA3ODOW7EIJqn2Hfww2PpnrKr
u/8ZBGrb0LqFu20NG8ibUQ9WFj6e0MeubokIzWORkJ/whxbGssSoqad4hhUXfkZDqBdQdEA+NoPm
/r2sTgRnteoANa+fEFKTgNTNMvisHI8NxwXgNJ8n61Xu5HSnzdMG/wEqO/Lq7blOXzNOF9V+oWXk
nxSDHfx16HuA5V4ezfGUtESGlwRGgNUYSgijMfNAXFU74c/MeklclE6LkGLe6I11ii0PkVUKvPhc
5KfhF7dRYBtF8Vfv6I0wue4rkvfli6+gehaPx8dxYRLtBZugNUcjvzgPSRkBNxOYqAJTQQUZdl8q
OPD8YmYn+dHPjCS07D7xVWG9At2qwv8osJjfw6dD5KtFZPS7W/4IV2hq6mNVRSJGPofcZ0sM0+pb
/Rm3omnq3TYVc2PBBUEZsU6zQypK7/Qn+jMCu6vnFWiS5TEIr59FygQZYIl37Yvp/U7OMFLzaxO1
WdZkL5nG/zOtVOYDpdmM7wy0aGeIZ2hZ5p3Fdyg6Kx0C915epHYWGH1CDf6I0FwftnYEmJMuRtHr
RHHbxyA3/IjTuizTxiaqFzli07QlleHL7G0IEDv/QIn3KVvK8CQRMCXzcIrtxyP4/cOd9h6OTYFv
3GbDiC/NFpOmyJ4qD+msY9fpy7IGHU/tsUhAb/xIxjfM7FZJqf19luyWRMXKILcU7wmJ9iKJydWX
O8NVDHFPDLHNF1SnsNrN5I/2B2+lK8flEg4NgHweBplE8dORAOrJyRgNDAg17vAPy/8n9JMFS+x/
HFIDxNu78Q+vxGskGjYn/uYxD4Y1pCDbPO9WIOqUAYEACIDyqnyPFwLunbxQW8I2ceuMtA/z3z/Q
ozsePM2sPGUL7tKrx0Kv436/MzzczKK3bQVKbGZVyvisy0NkpBFk3zCvj5HLwmNSZYdJrXZs9Ptr
sjppkI9jVO5NE9EWSwSatRQkRZWsdmI65RMj7reXBdft2rckIrM40axgh4VGkk5xZWtewFdCTXaZ
9udEsRdpbRPwol8WbBq9QhojIcadyQY9sfJk+CJaJ4NSMHLeVt/546jOuZWSXwfTlBWFMZw6VKh0
3W/GLz9E0POBpCvyY9u6tYiW8niXPRRDNqdfjBb+aoCoOaA5mJ6WtSoJJ2glpu3ydM2Y0Ux6Bqml
AOKF0qyIwR9nSKBsRB2rkxsD6yKNGgKtQE7b7ILiBcDSTp3NcdfNkiKynavXcPahqah6VqOLCZ5P
Wlda+cTtauEjk8mqnO5DJUf2qy+oC2wFmn5bMds6DWJSwfmTtgSj7KJv5eNReCa8Uvfo6/wFfqNP
J4YAInHthHxjb362w6926paHSfUJIYSQhAqnOhxr5MY4gsrWrKV7eT1mVX/n66Zvcqdg17vDcfdj
jEgPpVYxUTziPP3OSH7PzAjxJbx505Rbm2FEzQTJwbDwOAw+mD804SKVV3RJQFyuJGXZ2B6TvrqV
h2DqlenK46C8/Xfe628a3cjGKEgoILfyYL736AMEwMxvrSWKADAGYLHgLsMLPd2VgRrz+G2x+uPy
pT5f9G2RrPBjd0HOKlK49lm5VqaA4VjNF3eAgiOuwQD8SePrH6v4AdsRqfcbz0S0777cBnDjcsbY
5HVTE/hdYsm5J2bVYwhoDtOlo2AUcI32J9lEOt4UH9uUIxGbK3iCkukzvtQER6r1u6rB2TBPUHNn
wT3kKppINcJv+sFbqA4O5OfCuHFdWvNFbzWVDsZHncuYy6NWUzcCSbr4gXFNt2SO3uYzsjlxDpDG
rOD6DRc294w9b/JlS9zN3PQGOcCY1tWTBjVG10kl2LH3aWGqonc2aswDgu8iHUM0jvvX3Zklvs/p
JIvzeLMa8cp9Phu3fAlgZIJAF/IxbAsE8u1fUbhy39iUGqsBffrfwnOiRCGFyaZZ3Tqi9i8n0ESN
p4dbEuLcFkZCw5ySMyoQfHo6ljC6eRpoogsgAbn2215IphiCHSzOXOtQfM2PIRtxAKFBHBwr+0q9
jtr9Xf4lRJfmU7FpxtsTlYB7tvPM26Ve8Krau8m1UHb4Xw+h090AAG7lMIt9jRAp6hBVSnMzKTZC
RsAPNHjAJhEYzgj8QPFUu0nOHZM0mI0eUk5RiK8Ls4ARbtNUWPhyMNE0KkeRh936sUxkshEvqaSu
5+56fH+nr4r8ulSDL+DLASex3K4vgRAhZy3oUEsOjSPSA8Ilrn3L+OA8LNDO3kq7zmUPAtLQLWlb
7peKEa83b3IZYnkL+xOKcOF16ZPIvpPBG87jMm1V1PDNRwdg8jh8vvF2OrUqXteoRzLiNOXMLDuL
QAMBVObEDTiS80Uwga67atJ0zF+/1/tEMCNKE3wxLoFf5+pVujuaaU1T29nJ3MXQyLE99V5VYEig
iG+2GIvCR2b8vTWoCIzTuXOuWPSzAZMS2Wj8AvQ1Tc1EaZR7VPff9kO9DSva9/MzFBmb3UJZkRV5
6fy9rtDx0NFzRTYf+innvrX5B2/DPEyL1ArEl1yDGPmxYm/qJgqMro4AkkcviOz+P8FtGORol1nW
Z4keNxuxOHh3ttkzfRbH2AMWsWTI+7wTTuGM5SK05CgVX6115MaFkaIkLbasc6Qix6qR604ldgHn
3VAaGBlDG/qJOpPHIe1g+nzbe0EyDeu+Yw/oGJTmJFkZKLkOIHkh/3vkF3lONtwCqLSsP3iC3ggg
yQ7nb/kmoeFDNXfGKJlcII/TcVo9nHCd/FPSwF3sXGH0rknbADIR11XQieffomOZnyRerhiSJaJM
s44xLR3+Gxu9fTkNxqBc8M4jJ0ulep9lKar81DqngYlyRBUdgRKx9oNGjicTt7b78jORINH81jSp
U7R6YPwRHN044k0AZkCseUt7MttdHF0DVQ3CcYTKZpaATj0bH3ZqWmhYbrBt5Tg0TS/wRNsrRIjN
2roSpNTtqyuqrTMW3AxQcYHKFYizR2Dw30Fy7LWzf9GcNZm73hj2Y6GhWjtUUzJMQm6KtEuqPnh0
jTKVKzoh5JOKH7bzo2G6zoTKgwBM82L+rNhGD828QdWf4jEkM5/hyS4ERV3N3xsCNuhHBvgDLAPD
jC0YN1S8EjWPEcFKjQc/h/BpI0HZf1IsRTlDGI2fM8EWh20zxO+/FNNxTM5UGK8Lb7xSN6/QazKs
K7CcU90VIRk/0zkqT9et4McP4nJwez62JZ2b8nOfnvtZLWVSDf+i5S1LkjghSa+rfKIF/Nf/f1oQ
lujLYiUe05+P9R9cUNl3j/vpIcAFSkXSOCsEW/Hb5PswDDszVmKFOfUkhfxbyUY2yFC6h9x4hLol
23wWeEaJJ6zT704whjLq2BUbuW7xh7ePDJ+G+rTTNLk92uwNhaM7JEb8jB3g24qX2mt8qh6PJ+EU
bDymmzyIlmeAwlf42iFtpeCuc4cI3zNe/QHz08Fv9C2RrL+iQfpoyS8mJ8lamwRIymb2T2+03yI1
e1Sy4PbTJO5SmEiOBI/wsfNADAQUVWQivzdAuAmAzxHI9pdW2+kyQ4a3XFeCUEZNLaE6UTuA4MxZ
12l96VJvdX5tUF/GMetPHAjN/GYz2367vXEVGJRzh0fAXOATY6VlC71HHCbUsrg3iBROQDNfrMPZ
4r+d6ndDUO/lN5uwE0IFKrsoijH8uJ3a4jmFnHDAzncdrYO1IjOiLWoZJMyUDJGg7U7QcMEK4vdF
ezLeQOX214GgLyoYxYo3NRvMNCOK1iTz35Jjd0MvG/lA+N1plqC0hMSsAPv8NR1U0lgsGcZ3lB8w
SRCPnozBQTDCTAHP4cdcwKxaEzURwhobsRfV9LX7/bpRYMlWz47r0P//U9K5XJ8B7dEfuIVFcidb
VKGRq8IMqGE7upMb5icx5CjOyY89kj8iu32iaWY3/xevt3o76wKxDBxRA4Z4mFP53bpEeqbotbXg
6KxaRQ93ewO6g1ruaUa2Ng+QqpHz9DcXQuF/TJNbg+Y65F9rTB0eW2yLlbORJsiiMmnpWX6Ej2ov
4vppk7qI5XbyZ/216UcULTY8QWnhT/b+Kzz13zNHJAK+iZpi3O/Cx97auT8maetqhFwJauSSFRzv
sfvDWdzd22YOspXjU5PmYayG1ySYFPKx+b9aiB4YTYXAehqAyiGh8OigQ/HiH3c+Q4z5ww8vNjLH
sjQ29Y0sTsCbCdfjEUBdnV/fXEud0QvUKysMEsdg1wLFDnlaMZZlSaFH+qzP6VsJoRta9Ym4xEBi
PXQ02tUF/HuX2iD/YXRI/CtA/jqoIELupuWzMAQjqhrn/xf3FcO8U2C8pTKIVJtRT0c30cbnEuhb
A0fScq62mC+R6KviSJtbf/6BjgwPceCTmg3M3n2/3qnIuQYzaatcfgz446OikZPdMwQ37VfKxWJU
sovXlTBY+P9rFZ2sdrPjn49DAdnAzVV7cvVwz43wqLf8Ub6UeUYA2cn2rC6/5+EukEX/eSslvKk4
aRX4lTJMJngH09tYP4id2/3QO5+1WD2qWIeIqHH8Ws9MYS9Cn9aQfdwBdFbi1YOCVjBSq0pPSNXI
cWVq4dGOCOfXTbgWSjMbuBgxj6iEhfmLMpvzhySg95hIXKvrg747V56+cewP9oRs3XFFcVC1+kuA
FKWIDIT/93SFo9/Mpw+fx3WSNrL8ugvuZmdIqn1QCT/SRljl6m3BRmUBEHclEuucNN3ao+X4ul0m
fc1+sJ++kK3L8PGd9TaDsdIjdI4lfOwoTAQei6KNy0akAsWBylEEGV7WJfVfSxRc1CEz1rSGu/H6
XtOh3c3pyPubVYmfh6QhZGIZ70SW9xV/kZpUYUs/7APARbthNarW0WM+vnHkmHph2UZ/J8N/XSCB
i48xO0MjyszK/gMD0jpuPw16a/7ImZNt1mWo0GQTTFm5qY8G8tZYX3E19hCXPvzr59DoMZvJ8wjn
dO9McyIMtU5JzFrI35MCs6ZxY7t9pw9DVbRUonl+HDFsNYRvpFX4De0A5aQfknpJoFKAmp/2SCty
8egK1SlwExVEkSPUr7vzRFNH8LX4Otg8qj8oskUK6+uWC9UxTzP0IRU5UsQ9bVWBLTGfI/WoJYFH
XxYp3G7EtR9E2uZDPAu9aOPOo8GaTvMHm2ElKIBmU8ZCyYym31fZAYS+PAbxmo2efoGRUSf2LTS8
WKd7tg09igc+iznx2qk1IpRocB9Y1tnVmZ3LtRWIMaJMVEkudRuHzIeGoVE4DOP7bc6MwblgmLyY
cIoAMevFaIC25DhahRSXHcxlpUfhCyi/bCnTZKTAgOM9XL1EZX6RT4nSrg1uDHSqJncj4J7XMqEa
24JRUrpBS+NyQGODGumM0pZePeGsaooDf7EEjQfAT58g9dy/mTzGNz0TfutebeGh6039puDL5+eo
TKxEWRcIQyIZdsIx4s9O4m6mMxYexkPx8BRxCFB4RUGamnfOsTxhuUB1iVmPhJVJed+jBLrtwjc3
f1jvC7K3Sx91rKceZb5U+UNpd5C8shSbTe9LihaCA8kNZDzS7364BDrtueS2FKozZUh2T915wduD
oupiE8V6XULrjPjxRmbCOhzlVTJmOZOhMHoUoiTRxT9FU21fdbmcy2VPuq3FKrk6oqF7Nz4S/Gk6
6pn3oyWChsYVFVrEhjrIyk+5a7ossBnCouYOsPun+n4HeJ2oSHPSWUk2hS4QtwHvql8hgGsd8TxV
QJ34YssHlffTCrmNBIH17BYow6lBo36ngE1kZbLIAO57otdvTKzO+SVpdsZWColiUPWbcoF1NuNz
qx+jXhAGwOsj6KUD0t5GeLz8qnlZNKs+L7Y2sd/UCJQ8lAW+kRYBKDgw5GXSoFOJkbcOPDabpHmy
hAsmP6WLRmJTrx1l+EZ4tcBwQMqKcyutcz4Q190XVgKMU479Xd5pGQtLRcyjHeX++NPzKuzofTLx
9AVUNUIlTl1RjOl+6M+iyzmaROm276i0033xLeX6/OQiA6OWySfccOmC2TsOTq52UVWpgOB8xyW2
P9GdE8WFwXI2IBWz/QjbLz8lBEbfnZYQgpygiZ+XK/9+7dTmGUZobr1RlBtVfJrHQnB6tM7/kAa1
1Z+jGDc/+mpXdTEvSrIe4Youdq41DgX5lrtUGd/kOVG/KT1umUqDDQNlxOL0UNHuYl5fqqt6lyT1
jKjNjh/h58u2DKwUf0uYHdfGctwIa/2icn/rDBxM/wjy5lmPPBXQi6PdnovOA5FKdTPZvQTSAUQd
KUq2sVxsO+WNGkUExrWIz/KS4tr64ixFHxNz8RNZfZx3TBWfByMZ26ACDdu1UOEM3iW/UFhTEkbC
eWVVpnaUk4m3JQX0h9mFOiMP12ObpW+9bpiJi01t6V845Y3RxWFISvjpTCpyaXsbdJ/74CQB9tKW
yPCZp2hK//W57lgG24MgCrSxOboCQYN3Lcqc9NVSluGsHeDwfOlpuOlZLIIFXlvoks5bLwH6uI6H
qS0gqvfnmwcel4BG3qDIwIWskeR54la2IQZtDUDkfOaJh6tss3UHWhImuNDjyKPfs1ZyQ3swLKqy
pBcYuH5DensvSj04fHnqhD8wPGzFzoE5a5klV+0w6XAVbkE2ZlW0TQ3g8v46o1/KsullktSIocs5
tlaLBuGB0qvVyGal6XaF6QqMRHEudOQSqhHFExZBtUwRczGY72ay2ZB6BQMtPyRPYk26eHaPIN5/
5gqiRz4oKzGb0BexH17mw9ofJ6213kcAWMwapuOO1Zct2JorWwu+lsTvhPU+y/1jDN1s64tokRR3
4cbBufVBRkJp0ZXZYukHYkVWpOBU1N6SAMxlIBZxc1uHNgo/acrehD4YzVqEpYF3GJr/YnS0aO7p
Uf1Byx0ohi8hWI14bpWQFBTUWM8+CeZcRX04TP2HkG2BGuyBvrX5R6XDVRxqjF/YwQnLNOefnrmk
a1h2HjHrIDRHf6Sx4f7dFMn3Y1JsH5Bt6A0rVHnDgFnJIDhl7/vjouYIpRe+Sdpvq23q8SfWGLtu
iPntB7UjteebY5d44FIeNKbQ1XN/XKa7mdMVHV77rDaQFdY1GHAmsq5Dmc0VTvOt0q3AUmd9AM9Y
YriKa8evj6+dHqmuHNnfZOUGmri8zAAtaezIwEA4Md3fc3r/baz/1hz/tyLYd4cmOsWJhff0RjCk
4DuIu1hDBdXhzv/hYvSfdteEq3MW3HgviU8BELxL3Iw18lE1hi5L511KrBdLjN5okrhnxl+DBHhj
tL0sXdhyrz+jQinDhLLmesOl5eqd4PfD5bstlvRxSluOQt0CvGjdPWUfIZ2DoVgwTTHpi6k1kKEJ
9lk07Rs0MdfUdV/UcAGr8VczrgEyHa3heTr8fLOZkJvQnD9G8UWFfmAJYGsYTsYC40xnNZGRYFcR
7SvAjyy7q9B1Xp4d0vHJGwXQ104nLJAFOkpznDa/wH5TKJvLYmVpbPWFae5q26JLC+NxvgYehvpI
94gfJk6vbXVWQHNn9mk8t4jBNMiw5R/xMwh29DpTNiliNy1sXzXHk5qiIJNAuiurZ8EQmErsa3HT
pCd/IjECI87EpBQnfwksJYHNdwoIWG3RHo8MisoNgTH2ABnqRwFHkTpItNYta81A0aVlHJLeaQ1+
ufk5cjBWKq0NVAbd82wY4d7SL0PX3JdhBKMfrC3NF6IieMdhi2o0zWU5uafhHjCx0GDy6PrPYvfD
6qfFScGixIulVbGbgu861JM4AYX1PiwmcTr9a6p4sfiDZcvnRuhQncPPV6lEvrjzDqsE882lUZB6
gGu6kRgyz1dJo7RS8EpjIUNOcxVtxSoLjjU/WIAn/+wvmGq64w+daIagWoP2dXHpWxdIJhYZ0md9
/ktG2/+9+UOHnkBQloYPATX+tcGCmXcLKOlmvNsOqUs0GLEWmrRNKLDXH0tnV5wjrFm7zsktkPUp
/xhqkFTzfUcOOIw3Lw+2rrl9c4hn7sX1m/CA9mTU2J8tm7R1DfJ09KXpD08eRHLbCTUaWiWVck8X
iiMTa8aC36YykNNF73gTJsKVIVwypCuU4Hc1droIYjp8hzeXLwMbK0Pu1LmFrIEAmIteTvqHHhmi
lZaJgY51jO9iMdBgrc/qr/jqFlK0ITJo7HGKU6ZnNFIxFUYwCHaXf4pMoPmoOzq9K/3VmQuNEHPe
CxasiNJzcWhXJP8G2Z6MFP1gXYfFgPdNS/mltHTZLwqprZJJAxexq4J1kKwTcagfMoVFWzOMlbTO
l+HPR6o5VYQiImd+kRZ2uiS4X+Q/AxW93vq5D4r+E3NwNf6bx0BjzrZ4MSN/jqh/1vmEi0Zfsfxz
sCcEaRAgPeiVqQJB8j6Z32QXWj4yMnEojKIOgs+9YB4PSiA4mvWns8mC248EiIP3rvMdovn/WaKK
Xz32mRNIbYkz7z3hXd9nCF2Eo7KfdX6eJZqY081GGnli9+vTCa4fdbyJTqzmdTx8aJFNDWAzXIcH
R6KOz059zdoj9NQU+ECOSqeTaMTmoIgQpdOV6FRE7w9PYgsEh+4agwI9oE+mEJ9pudM1Yeq+hun7
dt1/Tcb3QsZ31F6K8rVKL3sES92NCosbAd4swjLwOBSOSFL2EQ8GjOTkH5CKXdW754jmteUvy/y4
84iKYmCgwmMiq0XkKW781yPx1ddHTBypoSduMlpWvO5GyjpPCVoLOyEPV7HGzBrERg65oXcfjGNJ
OocSUpLTKzkBsHbTbz5Mzv+fihqPvVgWJEOMjUz3khk+LtFbHQDvzWkjqDDcPZ2kDhnQbeQpTp2u
ug/YOEyoavVH2sqhfbRUjjcoMwW6KYr2h3HZ9j1JwLrbNvZB8f0ScGgFrcyox1I3wb3Qz6irpaEN
zKstnDomxU0M5N6rdooTe+dF+6yJoIldl6pu6O9RoXMoMCY8ODIWqMsbP47ceyzUXdoY7tHHjpoZ
tcJADm4wTjC0GPWLUgGo0jaj+dPMHZqvaCNKgs95ykDqDUVw6WAJjUu/7VQSovowzkyfDiT7yNMA
dmsZTj2IBb9kIQ+bPKaaeb/NWbPrlRZoFA+o+4N3Fr8+93HzZwqI10G+PI0lktBdVcNYUtlbDLrV
vw9W/RWQG6COocPcpZiduS0W7qUL0OrBi/89JIANn86ZxjPz1cN9zhEq1pbd/PAkF/Ad0GRZLhUN
t7v57M+l4jai2qGX4IWvoHK+XWOvPUI4jrVhN6tzrgBtzAcDu+Mka0Ako1VuTB6qbz57m5SU3B+T
HjvFTEzOsZLCZuvQM2DNQG9kLd+TXT+NMCXxRLj7w6I3q1I4INvcROLE+GmrRHd4Jb3pgzuYKzGH
PEJfZyE66RnYqZ99xF6vXtDpD24tFVf8vOTOjNvMxTbyvdGM5DjdtXQR3wj4HQOsIx3EI2hTS9QP
i025dQaxy2civeOhygzoA1V009ZLw9TvmcgWi9k36YX+WpIU3xzZGNPc9YQy/waqKlE750BuyKqC
AE3JGUd4RLxUBjQGxWG0fZf7XrXGEMsyGCa4tdhHUwhYSFbsH41s6by7h+ki+KozlGWC920iwcZZ
iKFXqbTPtWGVmJmC+eP0CckcOc7gHSRTteRTdj8AawUi2zOcPLGkgG5+RHEYPPbCKUTTB61NsjU1
mYeADb6SbXbo52p0KDw/6yxI2uDD7xbp7D7qbIzzBPsxXFms6fkKjyFyY0fGk7crz1Uv93h0GO8G
vhrBeZfinKsZgsPbLNDpl0nVlZVnxRkNkYQxYsLFYmKqvDZer0eh7Dk0GU2vcb3ALvJYzAuAEkdG
Yw9S8IbuSlSPY8ZgoH/qB/FdJWeSDZi61PUiRI2fj1cDDn4IPDeWeXm806u8hep/YO3jFqulTAKC
cT/aD8Z8adI3HspawaLqGvgWA/xaMst2RH5lTAxRNdR7VezBmN/oKE8bhYcJivNn89GGfBHRG4LO
RxggN/87T3bvDO/O+UjVGk+UL57FszbS7i5qpaObabahi91oiYxsvq1XzX/q+uWluMjl9/tZEk82
OjvYPQHLpOdedqh+5dPJlxivDa7o4GPtYioYHAmDnaviNTyUi8jnuDGA6UPyTV1kwDSJrTwKjTpB
P/t4TTjXoIsXUUPwJGI2Zl527BzLHcM6AsqCZkZFr3n0ZJvy7LRc+/9nkXzqgjKsS3PFvSarmQo2
7RgkeBJMNhl2dO4SxZ34YLxAmx6mXJOU7Muaxk7Y1b2Od1mzeBXpAur6eiuk+KrlWTqeHGdbithG
oSV9IGk7d5uBT89XtJl/zl85Z6uu25XC8Jl3odirGYYvB1nZssPJyDJIGFpatIcNTmHa9tXditj1
E+T4W1hD7OR5DseBP+LMn49IiR7ZB/bdbz59xPXJC/zEtTZ8Se5RLelELjR7jXjpGVYfsXQVHzk4
eJzo746D7zC1YBfxa643iq/m2BoHV34BokNDRlraZiGCgs/1QWCci3sgbpnT0GggNib9NcPSVNW1
3g7WPABmSd15amJdvi/D7OIFpEHHgZroAdooUp2CKK40XmIGGFWJpIo8786M36n1E+N8GsfheYye
1YjgzAV3q55OQdEM4GGgLAD4uaWyfTlJeUHTgtSOzKJEudOWdE6KT0JmW+LsAxii1ArKrxN6msyM
dU+xq7t34nn9O9gyt6i105g1lGkJ+LEqNqeoFHmg8FaE/aWb2m+HHq2MuX3pBXoD6oiMMj/zkXWv
VSJtfsZHPplYsK0Du8AzJipHuAive3g6EE6vu7VW5vy37zi11+7LY1RzdX3wGmCEG1pAl3UjKhuh
m9/+dLav5x+jOVclOh4y5GozLYiQ6zMR7+5O8CEVgBG4MrYjmoey3+nZ/NgolMT2pK6oXKDYGAb5
AiOhmhsuayepbKrlkCGn7INOzaaX0vMCSnbSMKv6MJi2tNW0dsSAe7KSP6z3Fu6y847W2vaKj8zC
VSg9zleaHOJ3M1iKDyP9O0sh5ji4vDOTxpIzaXdOv909YJhFjfBA7GTcPCMlnTzQ+pgqfIUqZTUj
BEBRdfu9s/VOU2PfA0tXKI1ThwlHkCfTCmw6NEJDpg0+5glH9HPvZypAXlom18h3r8fblXTNNyqa
3mPT3Ivdl4io8Ws7Xsz4ifOgBeeEciMclHJ/vaZxkGn9TALFoWaHE350wfPrNoRMpy8sBFGC01H7
Hmv/hX+yNQFoYu+/n+bFuozh/PnICu+8LxIQI5NBX092sboUHWM8CvaYhh0/8z2+Sw8AnMEoX5iC
iF+hc2B3WkCjuBFPGChICT667PRicMFBd0TLdi5VyXiZRf3DC45epP4ad37Ewt1rMbJbG3SfQnRA
/ng4x+TgFUPIjWrBtSJdEK4xhmgPbJlEel3SY+W/gfB44vVGCVvSJq4rrRyGopaAJvMtzxtUlBBP
SPk0RmxGhB59WTZo+/t5nxfXCqsiYHETTuUBm+XnM2go75bKvY3btj+Jstkh1Za2eP3z34PvazXW
l4kuB2Gt28rp3LCJni+voUV9smYdDrP3yK7g3neSA1ASvhZh3i775sCHN2zwGKsaaKhgtskehHEg
9JGMIUIl1Bdib35sf0LXdXzWMGXVPcXKsiBhLahtRjCBeqwBdpusJ9buLAtwqI3r+u4zL+wcMdV5
qTe7KYv7CoJ00L2ElmLlKgtfRhinQfqkS1+iukPsUMA2L5Q5pI10jVXWQQp1ywqzvaubxDOumnmS
7tnpN8A5Iu8efQ0uJyuAr2bmcmYAOGuaPnNwp181aAWBP3wipwwmsYS26VbFiOGXwPrmMLTF3GqC
SF2uYY9v1lRu0JZ2FQ8jXTYenJ/YG6biNLOJygoECjsObPekxBCdR3V3BFJJjKq79etjWzcK/OOp
Sms8NWZDqP8LBx0/oo0pNw8jhU8VlmhE8FMtLY7slsRN8bw82SX+E9uLQcFD0iWuKVRWM+Bzv6Mp
IZAbw9hTiCRSLsAXsCXDpM8mx4oM/4b31wgtnHen1UJfjllWtxNldp1UngXG+eTRA0Vl8bj4d6nD
jn1I45vAwJxBw9mVxR1N+lwZk3uVYm/wECaacbKbyc5bjlRorputJsL7JEMs7cS7XRef7Ag7i5fd
VFF6PiSy2IT1rg/CrALuImLzyjqMKKKuFjkdtkEH427AuGtz2D2igApM+NqDXli3ajA5UqF9kfp2
m5k5/5UrxqpI9hi8R7hzrj+HcxLqKiURQoZsvYewJMf+qW9ofi3wmlj9KtXiChZYhj6+zOCIrneO
t4bDjgaWJuZDWrbwWlZpbXtACQWnq4PJsM2/lgxBjg7v98Ny2r9zxKBzeILI4hB/b/IBn0wK6/DX
RP2qeSfa+cKO30r0V5gKdkB7jVQuz/1+aEC7RgaeKG6bunz7pddBzY5KL2WZSTjt+29pUTX0I81C
chdKlRTP+4FeCTOv3yoRQ4TI95YsyfirAhgnLTliTzKyCzyIEhtjOesPtUy2LZt3hf15gi3jZqMY
80JqcE4K59kn3OFWX2/sR6xKqYy49KYwZtlG1HxSAHA5DkfDK3jsPV5TA3EGAzvyp4eWoxb/wPTF
RnBF0hLIV39q5KMorW5i314jjA6KopoWaQMXEGW7IFb9MzlFa9hONJNkqV/OUoJXrr1VAJDvs50q
MaTtMR8aN6OfjG309xNWZfTMeu3qcINwUdjDV4F2A6Vdi0uFORdxESFHMf6JIKETTLxlJe0Rwe1F
jJ3HMqmCtopTR/e2ZyUmG27OS3I+ml+ptq3EgURYnpczVlvX+L10X6wRL8KGTF22aWw0Ob501LBb
pHUExDvACBByXBFx6SALULlE+q87NsHRzW/kNCKKvOudVZ5nQPTEgVZUyIZiSvu005TCzSRxhwtY
jLM8cl/2SzVPlMZuH4EysZpLFIAiar4nmh/YyMjlKERqlyxI7a9lK68IGHCmytmjztwTh7y8ci5x
Be5nsEdk74M2JJFL/CUJQEAa1j1ivxB4tiv07XFjgnL2FxdDQ7trWq4GHCQwZQelgQBRYgnNRA5r
1d8UfggDyS1B0HpLqNWe4F37m6QURtX3aBgbStWpkF4J3RSojrgFk31/NHroSo54IIYU3utZ7hFT
9cTmhj9E8AxtMYTPCc3yCX6BpvsmaiuO2G9GNb1IW4sbwqwPVE1XoRzqutB2IxaNIPKLJ2fpN6oj
56R2m/Vxmg77sjvcSKxVHRvgj55bE3R5iJCUiCM3VIL6fvsI/KJnWlztn3o9TPoVQPAehG6loyfr
i7h6F9p7GrMlDpA/eNIVY7x/hAJgTe5Ev5OjWOILUjv+DwjqaRVxG69l19SwLVarPb8v0BpurJ+Z
UDmbPKuvpZ0+O+VAHhroogjnS3bz1sVA1b1cTEsxfTbyOmMKw8TGIJVuhIp0LancGtiAYR/X+hyA
GXl9RGMPcOTuxgsnJPaaTpVfbJKxnotCihTa8g53u5PM478JifCgUJU3Ka53bs/+eEVKEOQAApO5
B5h9s3V5zGx2bTtSW9SK6IZtDUHeYTlIKvWseLqAriTJwFqS57+h/kFXqYJAFBNsc/n/qp8ZviCi
G9hzfkI9PbC3b7qlg+bZT9ZZVX2JJhUuMWqAoV4+uvQXBr5dmalOF8EuLfU1OmaBPfvm8ynJkSaS
ojw43rk2sasefWbDsK9PsRWn7wowpjbzgeYi5oJnFZT+CZSCaCqW6mhC7bQmLx190LeoRSvIExn0
J95Wq5papt7bjOqk8zY1qBINavfySndGHQ4rs91Vepnd0ZHMo2Gq17mt+tmalt2ogRqqFF1/W2mv
oesqbLVBuQ/VKCNzrTa8M96ADq10ZVJwzEZYTERENAGWduckv/tS3dmq8Lqb6LQygye93SFdEb5H
WHkrLIgEMbkmRyx8IxTNnpxW7FVIhYoGk/4MJufYWscQWvOjIuBD3gfogEaz+ZI2P2i1UsgKXafM
Z+wKgVur31Xb35LdabXqwOUzNwGg/ghJasLt0gEg0eFelcp3/nbdt5HGzruKrhA8jXu5C4cV4rsl
nD2uwcjdfGz+gSofINnq4TBoXjLHjd4rCpHeNUbm3ECmw/uEtteogdOeawetnm6skrzZxh8YsB0H
TNtpZ/bnZyfQulw6lxfaNLx0Oztco1PjhcQttzCSl4A6Xi25GhbevkplselDH9YtAu+I7wgLJrNm
y7g8LaLkzj4g1sWXDsp9jBtZVBZgvwXdhYlm2+ehGfM691Oc0GRr19p39Skn0qAH3u8sZVpLrcx0
U+6fnzWl0t0BGPchGqN0HxAFttroIjVOMTgrXShnPQSGliqId08dSt8opIve3YiKWG1R01wZ95vQ
mwoRD7+YEEkAw8LtkMo39ZkleRjYv3SEet07p28fOkq1JDZBdgzBnVXFMgRg2gNxHOZMnDd1deh5
NH0zBAmsoC0JGlnuWmBcpb9ZjZU7+uWahy5UC4hHd6jwQPgYaDk9HMA5ftPfqzagNAqzueiQm+C2
vb/gi/UtNvo31wvGI1cPM14Be4eEzOj51lQ2O+PBNHHBmrdS8pd1e68ug8x4tSq6Y8G2tzTrBL0e
XErnwQmB89nf9Vq8jBPUPWFSt9nt6O0rVrSw3nU6SCSH1MzmskNBeJ8SbavYCx6xJ06NixRmW6e3
qEYOeyqKuqchhZJOuSIqNVhnxQgWYXpZZZ8dQnQqrjtPndl7DpAto0rmeFDnKw7L0RvQYocOM+Ir
3h7FtvCPFVpvq4ujxTdqZ1IWhzOOEVFTGyI9f7IbK0BcFU+UlZODxC98drSD5bGfKUS2tA93DHNO
YJwdo9IOg4vDccR9GGi+1dmXUzOhOv+Au7+2zNCb6nPA8ydvxSa3qMvCY7jURCJpusxP/hDMzr4/
cXmKxVxhLDGp5f3iHxnbwMhaD/mtcmxg55PsdFhhtECgQsZu2Su6j+4c4TPPoKP8DFApKtujYpA1
Bs1vpnE61H1svBxSV3t06vBLJirTBYGCm7CJASGitEXdNr3Ft4LnM3pT2lKxnvIh8R+FFsjNHRGv
GN9h2UExpmVNwhAeghTHPRCsAPS/cWBCExkYaxcZPvLcjdkbGfgsibzSSejFF6qhb7LnU1/OYhbd
V2epMVCpn5ed7wlFIuqxymCMg2JVixKj6ZFdVJkAGyfJrf37TZvx8m2eIdt4ozXgeEFd+iwK7OaF
sECzdonPfZtSMFuTWQPwYhNR9ssaXZog+iUt864Q3JtYkI0sMbo8DtL4AM0m1hzWGqnzOW/njDHV
TYND0fYVkmApmIZbDX2zJPiDzXxAMYPh+XJdMrE7g0TH1Yzuv7BgLYt/dN9xyFsG/n1cSgyL3/7H
ACc5RTILJNWrTUDaJOyfI74iEsXj+0vulp4eJPQoTE/IlQVB/pn7St+DOHKL6Hrcs5b6w01Vs4ke
u6FXlR7NIjj1QZg21Lp/EwGEvNr64tXEKD7I6rj6gc3EwO5iBzixhSU49WL1s9344lchyYA2JuHL
qME21GXcoFjas1fLGdRv4HL9LFwnzkA3wNgenXBUUJ3XOLO7dxLGBTFTg1IxrwUAdo7aodbHT+0O
62pPmYLHzqr37Ux0wUW5mooVbQMRu0xt9yoZnt1NhFxks6eqRkLIEGOI/CDcGv9DHQAXGEP3YGfR
nm5SQUygEZEnV/BeJXgWqLFkq6FNf44dnDCRTTFjw5rYoikHbHdxT6uEQJIioFo2abeONEpea/Hz
oGVz2tqJB63Bs9O8B8Rf8Mhng+nrE7trLMwlMCuUmg7QTbGXL1Hrjgq2wOC8knDQuAvf+TxQrWHE
YKvVvc7sJ8WMPF1s27ZOUmfuhb1DGSjDvyPpDkDip6A2w9uRjE30+OPAX/8Fh9G/QUUSTCfyXTqB
7QAhw5X5Qezukp2rZ+beoTi7hM8wQt94tSYufqI7E0P6j7VCA9t0lCLDck3a81bnHsC7CvH30zPA
j/AyTZE02JeQ1JLoO57KrHs45QnUx32rCGaUusadUahfvTnODzbnb9c0kTSvWkpNPBITbbbL8w4b
oijrQg+lsYn3YQWUeoOx1d0GnpoDjlysbkV+TBaN52L+2d4r2hgCygC1RP5KcL3iKTFyidUc8Bps
FSwdmBp3dBplb45aFervJSH1X6X/mX7b5RVijgA8ZEwLOHEfgMjNqLwm7GbDdhiDu5erfX6bqYb9
Qhm72pzAqxtFaB0dWTYhcfWmXu+Xn3NhSjoPTLAaVBh5tXrFhhFz4Jpbi29Beet6Dd9z2i3OeDXA
N1JP61HJMep8E5CMRLWGUlEMJruEsR7sMdBCKmtuVhhLD7cVDxHkua50FJPwBnWVHh44GfVnMLvj
XpYekM52m+2nmJVOjXhc/gMKluQLr793hZT7HkTqFiTzr/3Ht0jNJxYF9azmGbpa0Fjsq5qxb5Q8
2CRJQRFX8tf7qFIgL9Xy1CkmuzJkdPCxGOEGQ30ZnBv5aglIkeBsP7uyPhYbBjMX/q0vBt8nnRAW
PLPti6m5OFKgYSGQ5j9yv9wspd4o7axtKqEBZkjuWEElB8wRn0GObyIJXumvUqE6++TSz1+pszL5
/k2T8lbpf75/rwpQfKohP3FdU0JVhxDAoJpE4W5zzYGJMwm1nmxj6i+gllDPgMeo8V5Qt7JhyUKx
4JUL87lJ5mmZfZ0nKSEbb9wDlpbTKhWJgKKoQeELJT8wAeDcRI0yVWqfHIedjr2IDqr4eIFC5NqG
2KMWoBRq6Ba/6qsUMBVRquj/YBVfIvRfJmgJndTIIvJTTFDxm00mps4C07vQ+9xssDf1oJZvzzzS
5dVv+ESVU3quIJQWsMBUOk7McLaKI9lNXGEcI/l9Xkq7y6gFsWUCVGYBzCu/Y2PrKqPKrdmXFA4X
7758WARnoOXz15t7Qvx0dfksCdRn+as9gnFzlTbHL5g5NSrnGUTmxbdFPOat2YJuAoo1HXPLyeml
uIs+RMPcpqrsEnQgKHfQ4T2sXedqPxLuqxm6XsZo2PjlpGpS2vXWeXe1fnSW1sBHTVO42e9Czfa1
1LgJ5ptEn5ozmBE1prTVjI8N6vtRlVxHMViziUYEaFIXq098uV+8GkFO5eqob4BLNE+8gzJe3/dl
O6KF48qPcQuaQjWZfZP/DMPZDOslG+kJ7pyMDUmsg6sD8nT8njqjWPDz4vhBnIIbKTnmpy2lrRip
Mn6UEL7hbnFW1bsypsYZ7JyBUvwm7BIKHlQwi/rqjfy4uct9CMkSO/K5K1wMCs9F2oxzazbBn2sl
Mt7YmQpEmNMLc+wsfWH94Us44QWZmArcmvQvjBZCMjrHj6ZKfkP+ul5OBw0okC/gYZR8zp0nnw3q
lUsC4bG2l2eclEx4pP/BA8DIgkD1F1ZTDPMpZqjdoax7zF5j7rEhfH1ccyZLB62uIbTxn4KlIajS
DqBFIsPp8+mF/Dmqm4SDJLcWZcfecp7rmBBS+cOLXSVxif8PTYMCmlc0FafFWJm9jzvoD/Jl1qma
g+idYSams1ctU4obIjr6uIwzWqSIV2GrCghD6iEEXYaqUnMINpGIkvvcWL2nzCtWgvmcZvaxHYSJ
w/Vi+IYQ3FiILYAxRN6PPXOiutEUgyq+5hVjz7cweBAlNusT6dsIxhu05Valrmx0scV7xFC3Xa0u
2v3L2kmi1ZHypcDCuwwr5+47JcFRTAdanwID2axcoYypsgJ4PvvZUUGko3yaEkYPWevOD1/lLAgP
M5DZZmduQuDBC/+7J9J37wZlWUnjm5DgvsghXJ8WFVb8V0X/MrU0R+WIlh8m2+iiXhWk4oKXd6KI
S7C5DT0mJ/zk52eesotUKaWxkNk75AgqON/ExqwTpmqdALIEVyppJ8y31twdGg2IIBC5wiuvc0Hd
smrQB4WeL5g7/D6ukng9kSFPyXUrzGMJ8FxnEH985AjQjzV4RjN1GbaqdYOCC/dwtWnbMJ6qWCtc
hs6llsVUVnMTPfXtrmXvtOgsAh1XEq47yjDsfyaddnluGXWcJg0Ez3DodtCTF+MKhCtWQK7qFO2s
yvkGeMGAW3PYCXTEDdTFfQ+uKdxWp8/rzQfLjVykpZ4XdvoCcPbctV6gn2WtNgTxOQDFb2PBnj8d
a3UtL7yjXkxSO4OBTdt9f07N0EexGVL1SX9aJ6lV2CngsMDbqMr8+sgI9VjcpU/tncJ3zuJlXKd6
VvJxxd/Xmp6WvO0NLj1W7U2QgYWLlMmp/e/UMgueubAtVBAochsYITdBHq5Ad6sOdBDb784J7JIh
2SowgLKDCVsj08aSAjUle1+UKuie6XTuPBx71wneWBQZKl+LtQKlbQ1J0N8Vx3EGjBruS8FJQPaL
A2oaADT2WyGakEv26ryn78LJmp7HVO9JUBCUwoPtLWu6QjbHpH+SssbAzM2cEx0zJZsxgU2O6KzY
Hy6xo/QeeS1MEfzDOhpPjizzPSzj+4pvdq5AhC60knurKaJevC1W49A4fd17ZT5W54EK8Eyh2H9u
/t7KFnci4voDpEA/+ZS4SouE6ho/ndmZIHBouwKa30x7efzpGfcL1CEAkGQUg8mKDolSA6rBba/5
gPYTd9BU2xmVNSEbDkU//q8+7v7UoMrK/4toTO4Qa8gj4fM8AxwDVk81AoqFIKmw54ZT1fKt1i3U
GAoZ4M84+NT6/Vbylq8LErE2QsHXfP+v48l+W+bmXMkqOjDi29LxA4Vs6bF7gXWOTJRpLQCSjl03
0tmGETtasvgLwI9TF8au9L4+8OE8VoJnrHFsmlTkoTfC+Us+IBHp/Ylnp5RMHvKC9oVUNT+pWueM
LkdRHpi1k78HA/hgeJ9n1UvWntP8K1/jkrg3fwGIGbNi/eTy7A43BBAdbfhrOrs5NNWyYffWS6KG
5NHV5OR8aZBBWNGxWHYxflO47nTPnt+fjKumYZS0GHyMvIj1vGe3W/+MRyQSiDfZUgk+ZE5Tb56O
227wUB1Noi88NI2Ocv04vdlXHTLzozShpGrYsnEtP8zuZpFIbBDNRT2WA/MjG78tYpjRbwnc+mMk
Drrt3HBW0DEOfffsCxNzDORFMMw0z+offVxpA4vTD7oTkP6ETdfzRwXX7724aNNkC3xH3IGe3wG4
iW3ZLWZIHIAY5hcBSGrOU3WKN5//d8QfxodxTchkQ3Qvl5HQKFP1OSDF3b2cfjp3CZEJUQDlxnN8
UNTlatcnCjlSFIwZbt5kvDenSCScwizc5Akago1/Q8PKFj5cm7LTsjvmOKiG7DNJ0WipvfdBXWdj
Q8/aHHTmXtRWxzJMc7iJmPQxGLbUFw95gQS4Y56rRtbkgIjodZPnf3IxUoSp8L4Z+1vzrDm77QS3
L2aXmRNGVLXJAnj1B1LX7DF4IHLLuYxZBYKK250oJLMihQY28jXCd57IbJmzFN+PdkJLqF7FH4s8
dBypgUH3IRPQazeRZNDSpKkJj0O+5jtxe1RxirNf56a9dhQhlYrwjvQfgTgWprcbqonvsIDsqulR
Ik9wGnT+ZsYUoNVNZPOItI2923EvassGP+HxaOEsruk4zbGMJo3utsMeJOfG74Rc0ZoDVme8pZg8
WVaAS9VyY3A0Bz3GnmEjHyhxO5co4hBjbbnTXIuktXL5JBlX+f9pRMcvExET7OQVpi7qTkou1/Zs
i0+cfirYadEPgX0pEIGAowQ50JDlJvQpckRrsWUSlYXETuoICGt0eO5jZs+kgcGVIadJDRCJmNkE
mrbDuBbeXAxDtLu418qIUZvwHXXBORb1sOGtGu4/+ITzYAXz3axAv8/neR7woUIJs8Wo2MLrHqzi
y80cs2t/0AC0XBgnBSeY3qkQ+GYEJxi0y6oODLmsPE524dBSSZtygnVQoYykiaRu2b8Lw350geq4
Szw2QzDU8tYVZYmBWMcYLZoAU+uCbUSF5hdruHMrV3qRbSQWF0GDnerF5kT2jt13ANl7rVzBSk3j
wOqADE+ybrDPEHWTfA650jpFKJNaaxN1k9WNVVOHbsXL3y+PYNRYK9QlZRLIrHu9H6pGdMI+B8Ra
N6pqr5MlE+djlJ1hcspf8ph+RDCWc4/4o+u5l/khTJU5HnCA85yki5/bE3C+6OMOT0angGmTkfIP
YpBArT7RW2mm+YNREEutpSCRUUKCXorYk30xxO+IyLesUnZsUDLj94W17iUj9e3cwnj2aR4sjGyf
rJJacat2SmInkhgzpKpntLFzmPhv9GhhvD4ouovBT3L4RheXXhH3ohLGN5I8Al7HdVJmleIkSYgk
KsNnCTQgKnvXM7nNKoWZbSn7fHM3e7N7c0r6+mqZXB2WG5eCa5bmAmRiDuXRJ+b3fcyLXh9oCuC1
CE62L4AaMq2EuTHorGJIdXl4Zl3wGJGfI6SqvnhNNhFZwn/rFRWZyII7xx1S9MtZ2hfuNS2LW8pp
+oyuPScAnCztyvq+2dxKB/cu8/+0Dw8Uhjp6PFl2lVL5bh484xdZbIMQRm7lzrU2WJFhxgJKlSTF
NekOloiWIwglHrNn1ViLQbCPIPlEG6EvbbBhT6GAZGezn1PGWeLW4LrFCdKuKtKhHXrtGn3KuXd9
pLljoDUqrAgNXjV3uRheHp0mjyV5lZrWimIUuiG62yV3TdPg9f376kXzV3oXrhjtKcBkokkotPbR
2QdtO7xrD4MijmT3Vy3o3rS3JuWW1ilwEVfvMx3slTuKva0IUaf1Wk3Uek8aqgopYWvqb+Y4wcFm
Kxa5JYOFHt7aPWiYwFsnhCmU5V+eKWo620epJSZWjSZdG1A6SJdXlDA/Dsio5Gv7rsOpUvYdh0Vp
LuTKhtKQ/pYjBJLL0lp3loLBCoB2891h3CXhPfFKOPoZAOIUFzb9m/ZHbtORYMjkX2MKTFrNzQpv
5mhg8Vk4FTGXX+VKo4/WLKx5fKlQU6LZwdXpZGUsyeKJHnGMgxtsOiyzChm+w16AGjIuatjUOIQb
CatGH36jMQXmjeQGMIhr9VHJ6NwteTMB0BpJ1szB+D6LcpVCpc7yWPlxGH3Td9oZBnDL2oqBJ8eX
vYRHKAfpettpRjYKDC+veHheVsLp3d25aTkux2UkfXDkPaYURzT+xbnE4c/clkSyn71VogFsKFlV
oIl9e/NUgtKsvb8b8Q6ytMLb0sEH71+h91KhBQDbuZpTmMd0nd4GHBF69K0MDf1Y2pQHeoOVV5Bo
JAc9G2guugo26SbP0qM6je0vyU/r3xH5ahSUdOJjvVO+iGfP2yw13u36Bj7Bdfi8hxRg5tI68SFK
nFoDUMtWxBqwnFrU58BTECSJnNcoOrQb/03DKXA/m9lPLgC1jfzyPqe27JZeJy5rr/BEhODPxCK8
rJAD+cRDXSwwPg0Vj0fcT+H/31Oz/NZoXCQcoJEsM4RzDY+biWDtpbMwCEW5Ci0Cx2YczPRWU4IK
La7OE4wfuTWxOMXy+oFi2o3P4tgLPs22Viy8WrgtddLQn8Nw4Ydria1yXRSBzVV9zqobgDysWbQj
WsGusXnJcpbQTdJgCDhRRwiNXBtk2GVDzopdJJ4qyx619Gajp6D83Vhw1cOwEmkW0eJEv78bhvoE
ju32jON5HKTdAKy5jQQuFxJk6J1tffzY+Nw5rDhB0Mjyav/hwEsDeFhP/GCZzofo/sZJ62SayQWJ
5FN8GgtEuJ4X1esSJPfwSaczyziDQsBL9s4z8xAvjvx7E43o9h4LGb4G1/bXnKqFjkjhvz4ylJ0t
8h4Ja4WBlR+6p+GaYMTcFYKUZP2+UCRtobX3ulD7GFQjOsYGhJiqtYJc9dMB3xWM/Uhlzl/Pl/u9
Olsfum/PeJEi+PhOBsFrsNbGpec6vDA7J8VwxmlJ/kzDet44THTEVk3/wJktowFFCimOzkqq/T3X
u3NRnbBWHCVE2qmHzjtJ/wqEPBsK8evJMD9ImCPSqOqmygP6EAaWscFvUUv+YVfGiNA/yxbIHyDj
dOlaMmo1iS9cWlPvjPVqwTnBOchoS5As8CrSq6xUOzGJ0n8fEShGQolxIssM2VoMU9756QZ1JKw5
f7jvsaJ3h18cwxX9HObbl+hz9JbOT9aVUlPdJoixuhiLpRtA4Cie/FXLiyUfrZz8mm/WLBqVTDDv
ON+PLD5La6jhnT1ozXz+od0hA4WcbuXJH3RcDAZnr1YZidKdrlYPeUF4ttI4ixk3aE4kVPGhlezl
E3z8/AoAUR/cZyQPsNvhIRKm9ep7Z1l8R92Fzn7Om+yZ8FSZ2ydx4fqSMhzUiFU/F6bGqMjdYzda
vbV/4JbES7W2uoSVmmyujRpCKeEHGQGh2Mka9+cfewCZNNU0B39jsw63IAs6wpCNalDjS86XpYhR
bbxr7Q2Kq681qXZQZjNxJjsmpAsCgs/UnODQAr5yK6Vrt57rMB+dJj2qdZCU6dslGA0jbhabGrvn
VMTNEUH0fQDOjauZIzD7nzYbdHR5MZXUbRpk9Jg2NXKA4eoHNZRVuTRYigD2xNojHSuUm8s0fmv3
+5qUyWLCWbcVP4ku1ThFEtFQmc38tcYTIsQgjU0W6IAuFWevhtmYDGNngtk83NBvl8TVYzLNN7dp
1arcAozbQhR73RfMwAn9OuLJsmqSdRJ9byd/1YpHX1+w4fJGrs8Rcc2bBy92F0doU0Qqw0bmhnh0
HRaz5r6jDQbGdoZ8A8QuDWHD4v+UrCoOtAW6TKR45WIUhEDCt7eJxITWJX40woRAjRoOarfPUjGc
xu53MFrRuRHUtx9+Y9KYvMCW+i2iRSVlHXKcFCSZdwFuP7JUM1L+9JQZ328OgPEaUqiC8tC3smvy
q0EpZFz9BrjxT7WDLey8YkXVAQE3bk8ZdpL76iCq3q6RrZP56BpjL2d/FkU89De9TWFJaLIhQsqG
EUGoYAIC6St/sgCz3u90K6ppL4t+mQZ6ibT734O6IZAXHzrYNgz1peuGMHUccE7w1aoCJzbugupJ
nbDno9P5HWZ+YKgGLjWj4IFFnbvV08OQf7iZrhsY2uAKaN7xsrnP/5IfUX1cE8hmM1SwIK1IM1Ey
8H/mAITde86iIh0a3bVyAnVXue4rFMUYzK8+HEk+OZrHbn5YkrcVSf6Hm0Z2OSeU5WbLfiMqwab+
YUuiKpGLTf8GlkOCIaobrIGA9LbFO4p+8EkfMxtzSm4xOlp7nxieFGiwfBBUh1JCC16S4/jtLNHu
P5AlJpdwl5zliCQa4lwtvQ6/MZgOvfu5F8hgtn/Y9kegCndeYNa4BhT5IU1KsqwvXPkGgbkAuxNt
YzE2KyXV71ylRykxuRqqOUJjlLrAIs23/rXCwoznwa8GRoond9luom0KzurnoWu2VheSHI2fvaut
o8KzQqXbsu9sZbHdN5fdn6vKMKWKKPrTItArzck4jMADZ4EqmR0BrkEMkMM4Ep2vwJD3TX9G0swW
CuGPflEPoJFgGdQoRA3o7SkRlw9BTGR44RAQymliMYgZxrMUzmZd/r1XrL5doVSJsqNS6SqRdhVA
mgtoNYM+rTE+Qd7yUIJ61pcs4Dt+2zuYRCWdy4GKKFDO4CQ3QKJxWScr6u8BYNeYe2XpA2d/vbrO
Kvllf9TOvAs7PGOaX7BKI8NIAufHchdekV5P1oDSe4nAYJ62wqwqvd+r5Mo6l/km86NF5n/EB22x
jzHhKfWVSFxWpBlnguHQSWBYAFvvDzibhQkCCgkKoJSGPrhNk3mENyW4IRWOb+a6CV+Yfwv714BS
eg34x/0SjNW/c4PWLr34TQY/fz5rbburHJgXwkeL8TStCz19JGyn0En1cKMBUt7s16btLrJftiHF
5Li4rgwHqNu3i9D/sTc+FgWDjPgrk7G+XvW2vxTB2KxudVkzc0fDJCV9lDIajZbhmKMoNneivAVf
2V4ZEV+Nh0ajhedcaHGF1TwLlKtO0rUKVALK0QEZ8rbxLbzRRZVgNFYyOnjoiSMklpqQCsKDBexh
+vflRyCTNIdkajesxGUGJDXhV5fKSDmFXLAhpdPGeenCbYU+BHETnhZHYqJKd09+h/5g+qJvW2bq
BO0mFA48+De4jRwxzVktrH+lRm9MuYOTTfbX6qHYRzqCv9OlQEC2W58eF2WAWD9Z8Ncd1hFogQqw
tvomEeQcLrhu1fmHFEb1XU2dqX7WrA+/JBrftJczWDlE+HxyDBey3peockSGFGkXQndgD8NfICK6
YSku67rvNoBwt/lHsrPoNa7jciRsUP0mL47HQeh1mLV5D/x+a7GbZ/yxHAEW8x3c8qwS/Wzv9sir
J3ERsQ5hhXBMAAQq77jK0MAmYz5qPozZB75N+nJpUImxSr56OokO7UBQwJONP7Bx9/g7PRvLnHRd
m8MqAI0ygI98YEUZNeiINfczJXYLhGN3BAbjHWhvtiqt0b0yjFDNDzTj62LLzlwvEid92D/C6tbw
E8uo650D8q+JOXTlt1VhP5IRYSVGZ9N/Osx88vp+7TVL3s+6nkrbiozqyilMlZ+aog8qYLHehVC4
JKVPWzKFXa1VoG8+prRTkYIZqUu4138NihWjrxmRd98oSH/RbRZaeH/NSN2z7yXpZLKTzrS0CuHD
IcUabHuMo+cB7bu006Y57DrlDohdxX3Q6swNArn6MrwKg7L4eYzYA+HsXwDOBW/+9unj5w6zBBRw
skN341N16mBTYQR32FthGYpv4pT1TKnjokVuGHTXTiCeYLn/14stCYcyL3tzhkK+UINRJUXy2n8I
gJF5S4IPkFuV5JtWxe4ojT4BBXbBAESwwEhzZsQ+SuROzEgMZRVhQKd3IGyTVZkpFiVxn8kFakqz
ig6wKF9E5RqZk7AW935h1h7ct7NVv2E4QGxtyY7lSUSeWhp+8sKN4lW1gnKOlzPuuu9OwPcoefsy
R3ac9v+dg6xTFqDWiYsLvYm3jjR4GM+2v/bpHKORMjYu9RJpZozmO8P08HTj1FXIou8bSJH057DG
79SmDoUAyOCJJnKK67oXiA//x6EZu7ODLRTU/w1IqZXSyoTVAa6c500WhtfzNi7GhhwmbjqgcTx6
lMOu+UYzYlVqte7iE7cx61SdXqY2tAngoIqzOIJyX/NGAgFlwoc4pnIFTNJjtJbo64XABm48FMIa
nltcsh8QBfTb+Qe09MqqNmSrAPGz203xWG1FTjdzhpiUFWB7gGA+DbFs8yO+yuOw0NfafmrJNciA
MUkVYpgOzQxUNIgDbJezMlc0JuxnbQoHk+XgNb/WEUfXtws85YCLwxHRwjk2Pc2kYlGI086xpcgl
wZCOLzfjwk3tfuFVv2wYCR4OBHdMNYScF76SKBRfLxQT+cszxnHtC3Kf7cAp7wdLfMyloIt3C3pf
nV3+hzNKb7y0q7mHQBLjxRNSVmiMHMKw6TeK/VdR/Cw0MpbuQ2o+WLzjlTTl5xbmlNgmPKai6kto
ibBWSZ0ri4xeKJ5AaI40R58bmzhJquM+qWBolVNg8AXDt9+iEzhOaGPun2HbLjoJ26dgpl/UMP3+
0/jXhmiHH4LYbplzwa5horgm/7DjKMhCpKKnNvIUUU1qobtdFiSZZ6Uio9wojcZPMseBRvq6SLcp
vqLgl8KWiO0nq1kKv4Dge6M8XNUcJ27pzViCNvnCZwA/txc+w9kchAHTWYEZvlAGQOtGj6CLXPtX
iMrwXW+D7BKbWCiD8vLrWHTiBOFsZCB2NRuD8+jND+CNJ8mpxuGcpEYasmzKPia8D9ouV5vdz5Br
fnAp0gwSzNZl9TkB4SCJU+/881fTUe/tiLW7rZ52m8fpII1ndaITIZ3AcYrMQCo7dcuhXZuV6axx
JRMr3/TCeEktfjTddYh5FSYjNvbJ4kR5sQ9TRlicQHJhBhKwZ3UnVBLOXInjsX+BqApvHDMtwySe
ZlHWl/9zrefEZ2vWzp1dZNJV34vSiUNBmGsrSEmXeY97UW0A+TYAgGe7s5aNjIM+EXgkdKgL05Kj
wOmgL+S0hgQq3W0WzfjtE/ajhvGDwdtmlmXRW/R6+5EzCs/buvG4mxcIExp7MC+/UQe1RFehGeIs
vUCIkHnNPLlm8l6wMGmI+TRNyL1sgysga6V2aOmCTnqmw1q26QbqS71Ucc4w1+TlNOssn8oQlySt
S6zrKzppJPo/jeWP8F9kz9scTelPXGD5FVyr7SC5ual1LFv0z/rKdOFbCq89LwUnRMpEqaFFnFuJ
fPZGsebcKa9lsYiMUvlhwuJcvhBuqOGuB9+sZwWHBJU+ELibi4sRZo1Re0NGdZtm4qqYWKZbwWNh
i7Ja9wE9jVx1OhaY4W2Q/NS9W/boGBSJMRyPuK0LZ5z4CKuj+H0BA25XPD4F15Zs7MCexJ0dW6cs
+bCb0jGSdiR4C/R11k964rVaOaEtm7y/t7tJZvziaj1YUV7P8WYmmxXQxqZqfeY1MTBQYUFF7oSJ
HL3S5UYX6eh9gD7ZffpPRopELWojqc/Mo8mZoBkqOoI6gXWHHMt/lSaKFzdMcWNUWcArHl1JqqCG
uYPwh46tM8ZfDz2iaMCJW4SGzNa94A79lsj9wT/MQstxtAjkRBLype81BRXF1LmgF6OoQNM6MqyO
OOJcOVGqbf6XiuwgfFPAgv0hNNIGxLiqPfKJZB3QodAGMSygYYYDEVwkDkHW8YMvr76Pm9V3gRbe
FMeEF+vuTl2+qdryfid99cqVtznB8ji5+sO0d9dUpWi7mVwmg83Ulu6RUyl5CgVJStHFdTxXJJVy
w/a9xDIS0MrtK8qNZdREhEglZCgCRK55qq4NNYnZcHEufyg7Qfo2dwmIoRFwUKVqSmT5ejeK8q4B
fstH5QPUYQszn5bg4BD1wjdr+lNGWyjKQUDgQQzKJCdmrvVHu3Wbs5ntbEVZ5WdUZi9kgKeZ6c5a
uBkLlJ3MRUSHiovysQgSlRRQqnN4n3l1eOgdkbucqXo2pXDMOHmKc51KZ/rg0j1sP4+Ysh3je3r/
HNFYTmBmZZnFVvjyqdVRIOLEq1V9WceeY3owYvCo/o5OFMWp82wrdms4KH5XugLt4S3WcVp//Y0W
OVuFVf9lx3yxVuLAlqGlL7Ii3ZAocyq+B3YkbJp2kTgl0Qn/+xMlgxIiWH65o9rTedSLPNESciGH
aYjvynEkScDe9QVAoP08aGrNxWLOjVZeWPiYrGoPxJvGSmnPNdoVIsz/N4em/UorE16T9br2mA9V
jqZ2x1baHpRgql5c8C567td41TvgP47CArmSddxNQm2nFyhz2zNPBjeRBkgeXTBLDel1X1TPHNNk
8rrkgkYEeAngN9SUEZFAj8EEDfClaHJgk3vPpbU5UQ+W5vxNqUFl9nVJAH3L8xGRz8lj6BYJH4ea
dbg5eNcCQniPPA5Z7fjlQLaidX93sO9UnBWFerEXIUyfXfZQDYdIEvAzrOP3qWQ/SSE0K//9y+d3
pODIVUTErVGAXQ+5hDZK/zBLosfnQJLzW3hH/bw1pzyk1YbnSiErWV5r5a0dONotPLwqZINZcGmO
ZvEPmxgYr8t+alq/rUN9IK6aFsdfVTUlinL/caVkCoj66Ij216qAn/iMWeZiuzzTDJUKHP6IYHjX
NdMtgujoRv//oynHVgEXD4pLyhiD3C9w5DXteSIAeS9uW/4QodoiYErCDVQBFug++4iQMF8Tzkj4
0OuZ9G5ibl7ubFD10BWGi7r/tXUHFFAmZH+2NwdupVe8JqZvgb/Lf3mwIjzqvq3Ja/PKq92fboMf
PiLXXpX9Tlo4QqSTmpPliWR9p9EdrskieErr7ACs5x3YNcI/pPk4p4qGpDJsXCCtz4LjVg7kOoCu
4gYviqJQM/EoNAkf33yEfhYSq9OoLVrAM+PbeYa81itGnIW9u8qrFGblZYM8/IzTp84B9vWfq44B
utke+Qot4OihiTxmdS/xy5bgXLx1akSvx5WLEbgAr7nDcyXk2y4fA/N4lG56V8EJzYp08JRPAQny
+CgKlfBUhQLmurdYrT50I7xG2tASgS7Z/bH0sNRrTViIfrh+qngyiEYnpH65kHeEYGrgrqx86H57
V01Q7y873rQeFyOs0vg0m08+JgoB2ngz9Ybd68HazjmZns2AAWv0/4xm6nlUmnPOK4fq1f4YsB5/
rt+oqHZ4KIW23bwhIulNXtvgqfk8IUS9xtYdNCcCOW+QaFMQrmiDUoVGB1cdEY3ABwmZ/SuR7Naq
hNWigd5hGsx2L2Qnv5HlIkVz/ccvcXlFaUXyvSZuWSkkttJgyMGoQLR7NiE8AgTPMyksl++eEY/m
T+Df4Tl4dc59col2mybBx+MPpr4OMFW3pftzYosAoGJctfu528bgjcxF03LjTdLm65guk9IrzQln
+AxqlHI598zVgX+cUuYxiS4B2EDJbNRPopAiDb15GdsV8lpLWks2GSyFoJxR83NjPGsemWFOWszb
RZRohv8JU4WrmZsdfEvsCK1GDXGpTzwCfN/TrDYI6CmyaDlWPUKZY3UxQhtbWg6flfgAW6LdHygL
f6JsOfdAUZjMhdZfGHL6LijMfEpNTwMO4BdaeDY1bOwENu02vWPK/PHaFfsUP/5Y95pe6sOtp0ZU
DnKHE98bkmDhxt+qkzzSccaQVC3L44lFMhttF6cv27SF2Lt6vfsDtsdkPPqCZmBlTwSizMnfGH/6
a4WupmI6Buyi+PMkoMImaEmDHjli6vxirlnOKrsR+EuSigkywP7fpvj25a2JyugOywugMHF2q3oQ
uqHacCS21NKrGFpne69RqdmW5A1Q7kXLejeNHIcO8AqKBC4HjDFf1ZIqIW9MYw/2bgnCthlPZvfj
TLB3wa41YsuIEiHFeGaQvHSmNe1rFBN14GHrCUKFOoSIP7jQkNMLn0yLxJFTTWCO3+XqBL7Zfqqb
aAyTcbUMjT5b8kdWzONyqS2k/EhdyzRlWuJUW6jhYDAZGStKJBJrg0ejYAP6guQQpHVRurRwPoUT
7a4uQEuziue9dM/BCHeoUbFDze2JwUX4i05rSCYxPu9NV5Go+cM/1k4vi+tneg/EKrQjPKM8kJFt
j7vKgA7uYfR21ef+udCLwoKJdDZIEg0pk+a2YzwAJ+H/WNS45a22CAG7qc6FGFBlZrcsZfPpQtB6
ZpTmc5649XyC4a8DsFxQcxbPDaJJ+UpLcWAHTYpFyOZOO66F1LHyoKLAMvI8r9f979Z5/hJGhmQl
UoTh+amMDE32MUcyFW+WCNecn1RBNHc2ENQcJFaGl/22op4YNENc6sND9JNdkG0imwnW2vYTPY0C
/W56mcynMWgRrNI0IsuhtBbNTmQ3FqWhGyBsjEJWAkd+MpWTEISiBRm0HW+1M/0nKR6HNS2TMqL+
LLdAyxFPziY9pIpMPGJ/6u8IOp92YdjYsSPi8Bm78NYOHS8LMertUMP3V8DI/+unv3BV8YKH84OU
5LYofq1HCA8+IYp6ZTJZkCAs/r8wLbWW5Fz0boxWiA8869GTX74mfgtOFweRcbCGe9bD8EA6ZzFx
y7OFbG6lNUsshIqBryCYAxRBZ1TmoZpG+FbZeZ5+vNSmmHU1S6JL9mPE7zEZ69yU2CHKc7/rBJ3s
TnxEQJioDDqkcOrDSa70HfWeiN47Osfr5lpeOnNJEd50InW5xldSpl6adlk4sWdKSwNbQGOyUw2P
WegZ4YAQPFQhKmKSK66t+2zx02ct5HhhC972Yt8I2yxDE1yNUyBSIWJeaJIa8wjL45OPPF9dPoev
3RPuXO1Z0m9xLzOB6XCMjaE5YiEn6/AGEDRsnkMZpa4Yhn2Dq30eXZkjUKfx6+XRJ/gPQikuI55S
LUKt08CTS8QZQsoYxozBJEPz9Z9fKSVZJhWDBvwKXVxBbheuZ6Y0Eo6nTjw8G/KXKlelsE+rDCxz
lAvEoP5CSfaJKCwVuXpJp73rKJix/qilIKHB3xYxqHO0qV/kTWUQe6a3aR/fVNgCSGDKtx8l7x25
MvlpNIkj75uWYLbR5ibsH5BjgCRSCeYL0X30Evb5FeouEoZJTVCkh5u5PrY8dPHSOUSD7L/SHBF8
Rx0MNwCwrKoNGtDNg2DqUz5kI8WhWC25cSSD4+c4ZQiIa2gpVz1Lr0TsuHKx+NxxaQsR4VBQAMh5
2vvoOahYiJS5yIZ1mqQrOuKmz4QHMMHJZ8O7zybL3JaF4iuyW+C9DGpdkjqTqk7ShhcQeBBnG+Im
+Z2LZpmQBTxKwIXf09MbtHm0vxDg6+URKEiW8kx2LvbMXAQK4KRQXYd17oCP6vjehnhxSD1PPJAz
1uIu7fRwMo3OpI2hyQa+JgqZZCnMxnHX/6ZuHVnMuEgTkXTR/0FaShFc0DONhhVktP6WuOqQydfg
AotYj1fz54RdKyPC2lpBFeM+GCCGVwbDjj5GrVQDHpaLaiYYZjEXRVFCzvKl0CUeSnJh6KinqwWH
IXNGsFB1tpV2zaOwwiY3eFMp03DTp7tiAtMrp/4V2VaG8LDmtafQAl6bhJ0fXg/QB5WRAIJ/EyXC
4034dXJrqT/MMjuwgdiJGp8lpHf1Ti4SoLHn1bzCIFRNRgPZDcRAr3nK7jT44GeUoXCLup0av9TX
UQs1U3dRfsqEJ3zqSa6WUnj6xnweSvfTVk89UB+QQ/sbExYg1TnKDnqauvZgkiDs6Ke5IngJmbe3
BmBThJ8lwCCUAD1jCRvVMHYAGEPtFqD+kSeptYlcUPF+vk1eq1lhvBWxpSSjBHHEoeWMsSN9Izfa
u73tMmM5JIO5Avpem/7xEo00kIvuzOlP7bTNeS7MbpAul39yz4KRXU8vulvSXnY/x1BeibOiLfHg
Bq+4TBqajehkwWQOBK/1Af+PnvWZkghspvljaJ5EQzIchCKFXiCPaEg5HKwYgxbIpGlzr4xXqqzN
k5ybQc92qsU7/aruaBRoJGfVoPOXDySJX8QMaeaLCOUt4IOEmHEc1gdt43JSS6jYtOxR5wK7mwS8
XnU+OoenQ2r5BAEvRv4M8L8wcpnsTh1k8xoUcelkOzM8YSrWiJ6hqx0mpGw2AoADOtvczQsQ5RvS
lSKpv9BLGT4kV80xT6+VD+Q+TiKU2DizQIxXzjF2xer09sXmOLmOh0gGhw84Xp94um7zJJE94uM5
njB4GxlHJTJXTwLad4p4Y68AYKeoGk+SFZSDhzuXyG/8RSbTFN4ksepN11vmOM4hFi7uLPnIqzCT
8hOz2T3d5YVJgQicvq3qYjaOSTFEMjwTARCtIxyERczx1e0G79R2VuCPGdigPgyJKNdNNZRlu6BA
60w22XU5yrRytjrYPuhmmVoi0zopXHa0+XZR7qXg02hcDp4UZS94fyIfhPqX2HnKyD44dKTddUFx
PvZQHLKiGAJZE6CB6sc9S2LR3bqMoUbtw3GVrwG7agIaHHbGBqP/4yLjeCRQLv1i8ad7GfEzsBdn
V+ygcloCDhwb4Irtf8CVtfqXH/sR41gqldtNlq4VAhZrQSYgHVdGyRBCstIkLWzeczmAHqSLzNQh
yJj1mN3kErIkn9xtBw7p4x4d9BoLuUZUHXmNuyBQ/uXuZFN0e4stuHLCk5SsafpYVtVyj2J4q0LV
euWt94bFu9VHWOgRn7VW2zONFmIrDMu78EIFYpT8mJPOJOWsEI2BWLQDrhs/cm9f1+PMhF4Y6AE4
nkzZTpTwdEqlrb1GlvqLx9lnQGO2I+/pcx42FLUycfqJYabCwOxSjOxs/J9l+9YUo5OIMCB4OpwL
H/2CX82fxbqxNPHTVPBWZyGy27C8uBAZ+bKD5sc8iQoL1/2LAdEgcWEheXvxQ2ZN6mquczaj5Ixz
NY4uZXVojnXCqFAwkUS0PhPP2hycHC0bPSC+D9YmfEHZyqfw105SATOXhwiub4Z5a4glTNQGXcMl
aXLWSfGC6OVkUYldYp0AuNAgycwyI87rcnlSL6zMiOzak1gSPTlIzb0pi3Z0f9vTjeVLZCFTmwPK
Tga6BvK4EV1fWr38KokC4Z6omeOOBKUS/fa0b506VuYDZxPcBMFZxfJMUku3uk0afX1eCFDze0IV
KbBFfIyg0JGtj579zx5j2/b2saTGsnxTCRKGUBlIV1aNtY7VCK9upHmVOoFTD3vU9ebwe7lpuLjr
QasZb9f9uuB56dkg2S2CKhqFptBspUd9+glyyI4Hh2hfhTE0bNko6txxa6Bn6cLiKt9bysH3xxUM
jbuJnFvQ3F8puzJx/u1RZP2WMZDGj8qTchlqR96mWQAlTFHhfGk8at+v6qJ5IpAsGGHcmDCW08B2
0tBBQSsP6i5VlBo63vUiXvHcrFOwBj0kAuNN8BhvKXrsBAEkKoRMuqFePMK7EumFY3I9wTova9SU
CzuhbxmJr3P/l2j6Y03IXD6onizfEHiT5DcAoSnT0Q9iAg/Be1hdbL8QUOwJ/+bFfZS6lwAA29K4
nmWrsefzFCmyzf4gQFedjdTIaHVIckgPyuGC7fTDZouK6mYQpueOroJJAhmhg459WI0JotLgs28p
vBeT8Vrja3b26t42hOFSHViwkLVcVl8j/Df8zytjMgdJVnD5H8VSDFROd9RwJWGBPecuSClblvHz
Wo9AgHZkwV1KADoFUZGWy8/bhuuVQuaZVk0nfPv6rgN6CEtY8SgxievE+rKn4ftCtL0xkjrJ6/X/
/NkeuT1Xz8E+VMP70rTVFulMswvzI7ia0fqKHNxMkweDarZLHyBrg4HanXYthLCtQSS9LzhurQs6
z6ontpF+qnJ9V/pHL0+nd3ls60JsVo61u84hd6wSCq61UMoE7HtdrlAzQ/zMKwKFq424QY7Ys7I8
oaJPc8WcG15XTenPIcYofnulSgMngQonOI5VdFXJ1XYRdJInromr1c7Tc6dzaImqShBRgYdR+3/T
Mq9GXfouYafRQtmaxw3DiIt6ngN9+rwXRES37fukEuOtm/bNU2SvvVl61rTnWCe1L/7DdTYwYfYM
Iggd/3oQahpLr7BIJAWdSRTdc1Qol2bIK6CpOTI/X4IVJw/X4PToOj+lgtDYlZC2GacEge3zwuIr
4IK3QSgZXln9sin3SfCQ2ndQ8gTM/lPUmywz+p60Y9K0/6WHFO+E+DtHqvvQxKBKCH2yVd6M2dLx
hcf6FxHEqYZMW2+RU9W5J7SkEGTZ2R5gddp5BQgq3DyFl6oxUNFUb/MAfo+4bzqBNRmy4fqZSlZp
T5t/zqT+rsg6emyslCVmpx5FoJie1kZY+iyYWVn2qk4PHiybXFZJtk0rQ0WPAiKzyFCYrZlwBT/y
6PXmwXJwQx911m1IMtRrOwGBrkehJPU6RkTPhmDUqmpiKpaYy6E0OiOuYubNCpMr7FfMNF8MCZ7x
p50N5Hvf8Tfv7/td2NP7xTZnFWGa4W4HTHIHN8GaNCHC7RHk/+gUc69ouV37Psy+ph+3RUS7rB8L
uGcrYDuwm76W321CWUOi1WZ9MDBB1OMNkovCenbjkTFQrj5IcJbPElAh86JwCPfr7zq84pCzybTa
KLerHqhg36adnliYP/sy5jd9Vpox2Ivklz9kV8emWzMDrvnq/b9yJIu71KCrSv05yCeKmK5GFfFL
vvDJwrsmYkktNfKmWHnsh9gE8x82jMKHJt29OMDRjvsbXfxVFbTkEW/AI+kh6kuaqkzGHVpNKs4I
vBfJyssM5rQYAYuz+teG6bwHJPkasyZiQg1VFh59UYzvokd75mCYUV6TWY2N/91BruFY+Dycwv8N
gKFUG/1G/Bp2E0nWzexa5Zjd4z9kh9+2zB9RY4PodVG/mLlk22j0BJTMjeeuK2+FvDWFfs8eXWm8
GoBeHHNAAt/dmz5HcfjFiTa6OwISLBm7T4Bl9pMpUKoaQ5a0Qcf0We9H2YE3oC9ids2hmESYLQGX
7QfubLsplYWKWpxcckYoz957oTLb2jRIZyaaT/oc8QBpJ/JQKYabpQvEPPkwxoHuBsBeti2fO/iZ
06E+71T+/kzByUFrT7iEiIo7zLszwsieK33GcUOB+thlSLaho4vpkhgN76F5d+hSF9EEMP6PFFpd
alELIQMqzm1RbGc8h3Mshg7PJJ0HJac5Fd5PeeRIVaiOqvzdrPJAw/7MRTAY8UzdOAM2HkFiaLOl
kX9OuqPdy50vgb2sP2Bx0AsQkc3w0FOTwrRWNrParNvMBw1t7QAikImY5BOcg3YYmZgqqqPdBMCM
Yw5giHY2F4IsgCvN919rj8hdwFNNgiRXc5Cx7MnZu1mKMVqYtKlcaCoHgfT18s7uAFqbrEEbV85Y
5G/B9WuNWDi2XDkh5179UOQBQNBE5qqAyQskezPkL31h10B6FGNyFSeGO67dIRmDClQuvlievAfK
tmtf0Vj4QK1dTc8GjK13auvTijt7uCg97+xhYgAw/NfgL3loedtuawXuRX01OKefITWZBMEsg+KN
Fs3l2vApW3MtKKHLgesj6/VzyNFKrORMPeyiN9qIi8akxHyndzvEYkXKQ8hO86Fvl57NrX0yS1Zc
HTthCgyJAg70Qp3EWZhh9CpbKeyH8qAza2imfTvLku1vj5ryUwxyrcr4wBkA+ZvU3jzHykKcWvr8
3l8q0plH2CqGF15X5MBs03VfVJQst4e4switlmPUGEoBP3g9FWMRhhezyhzc2WKUCIMyzLpn5swK
siapsfXpcLDzjvCS3FvAPL6H4m73xWQnDCUa3KV3zu8/zmnuCs1YjYo52p76XXOARvMnE1jtsEvE
E6uFL/I9KVLBCEhuTHcIEDkVBweNbSU3BY8kjkBuilkd/q1GeHNjCfB9NN/XcfjVac8l4pdwb8Oh
cS3TecBkLCnigEon4CNgWlmbHlUMkqWqNRo37lDWYICIA425TxCFcD3OjXyVe/D7lBkNvaLx24Qm
bof4AZ0nj+EMXsw6kPkf5YK7TChb5EPvgX5FaMciYkcUMYbHsdoQv2oDjhgz7J3crsXd9nCclZp9
U4531oEQlrRPqm7wG4TRK85MVVhRJXe76uCCDu/zMiY2BrXrikUWPGgRf+c4re9po7tMk6dze/dY
8NxKf7lxpn6J67DPrPztgvqh/HFRY1YMaCqGt6Y/SSHy6L/ybblf4GqZDcVFePEO0kMUhjmyIRRE
hU+dMpkyUne3oWZd/D5fbyYvfHVEIwdWuxMeJvYcK2m89BljoV5FYOy3E7SpEduuBApyKmNfd+jK
wv8l6Ho61btGArh8CsvwP4GLexPBhrivCWDuAuO8OGpPsW5hNe1GwCE4bEk2hrBS2edGfGyBRPsI
CazJhttzKcvHx3PWUDj0V0b1vjhv2DKLAk1QXmtZAuVIyjZmc1SRulPGWJ2a7EY1qbcrae1FgUht
lRYSd0ZOZL9IV+lBaknG5OejZtBypJmSCuf3p/XrsJtKoSKRSo3F3oTxvHHlUeTDDTxGfybZ6d6U
laxZz+d+5ODinU3rxMrnhYXZLHnb0YRsVRHHeq/B+TtFNl3lttwWvQnrvX21SiMrn5PeFQdlguv/
CfL5VQQOLevL+cKGT8FAgUptfoEyonmhkgizCIgwT/yyfYz4dogm0akRDWhJyzlKBrgyt7opruSs
ex0/whtZCS2rG35Jx763vYIn9DxSonx6s2Oqn8KQPMtSqz7ne0qCtIesQxfoChjAmfEoNuVG9+RN
ObM61Ng+AZJYJ9gLzswu1RSidl5hTPeXzQtEXKEyxe44B/oxvUoK3Vw0BcQO8u0+T6WPqZfNwgoF
Jju0WwSlUmy3pFLIv0A1xcIgGj57KE89J+QoEpKSoU7aFeAIkdlNQqQRQjRK27VHwcsCR8S4Ys8Y
NjqkAoxy1RpgHMKukcB9uyv8293NZz37w4lBxdbCP4/UrAiiLoOBUFn0vAbtR9/jSDZMIJT6UrK9
XIP0lbgGW8+Ds3KJMYSDhPqMUXXf2YqQbaLOPps5IWe4ZJKwgidk1wtin42+zj9hlfIh9/qojP5Z
94ePQh/q7FdlBbyQY2P3ycCzZbjAf+wTXwsEY69vMdZ+/pHLdCzMCsvLW3yX9fu5CJrB+ZcG2tXt
HNGdiHqMaML2pBv2RJr2THkGRVd67nGO3ZC9aAGIfo+xUm1U3SLgxFbEbNDBf93eCMsX03a8r2NH
ydIDihownWzS9r2bG2JbJXE7GwNnrp5ws6O758+uOOjMI03Ol9hwu8NZOhMp1v+NCqpVz2EJWzrg
hYNUlINOa9ILla6jalsWozcxWjhE8MDeRZzidYYcPGu0IS/Ww7eeVEEc7rjyvmRNRMN/8SvzXqnp
Abs9fMyncAMrw66nuDt32tciSdWEpdEiUvCOCzhJxgzjdQRbLCVfM3gzfOzf1uHG5WqAVol9W3Cx
IavunLYy5nP0/K2J0QHvyFLXe9NBIp2U3Fhg3wpK1440v5Cm/2wgP4cBi/3SoFfzvDV19mJbAhy+
ssdDBHmGKYyzrACi9zL4ZxiaS1s8Mn4yQ4Ih1PuU8wVE8h7Q7nb4LGAKAf7sHvWMkI0cyJFClHRv
I2tSJb2uZ8nZAOHIOeU8dsoKG6QWF9fHPsO7dBUgvSyCtrS/ugTG2CtEoVIb0Sxps1d3UyEbF+io
EC8MI2Phi+GhTgSEdvD5oCYETVLMNfySwqREmZqvvHu0/jG3lHig+xZIkXoVHBCOFiIA9GCTLBkg
ITXJw/rfLp5Mpn4Vqh/2fOosIKI8RaL0GEbdGd5EVAbTqYvHJ5TDAKN8W3tbgKDtWldZpCciefGW
+PHuEei4MH7WeN3C1XOFU/DULk8AwJm8k9cR72iTvrwe7jOWB89zotaxjfo7m8Q8Zk1TmkPTpENz
Ovdu6V4qvnBLy0PJGrIIilUHM0DKkEe2Sy4SAe/4kgacaEQdXFVLlKbRNuu2cDCa3OkyHozd5ezI
uo/PF+5+4fMjDCk6sVX83/6NhnQHcFpyc2BdFmU1J40XRVHPO/4jP+WDtsbW5qWRbggVt46XO2Zi
anTT05Nov2W533V6QVQgSx0YkxIScXXvFcsN5BJEZYkUSxqXx/EnPvycMBhGchCKZdYMz4vxBP44
DiHRWZV5HcjMP1G2U1c/1n6a2zeH0JARsOAI4CgpzCpn1OadX4yu0oRZ0crwQoZqVFk6Lqnhns/U
t8sbnDNqrNJ/4aRv+drvdVJdFSbgTL7ajk4RD7Os8s1rUnu+UQ7sFU5dqFkl7zgJgBGavgExYse5
Xq5/GUDr/3z8W7galmQj+vQzdrCNY8t1032VPaDvscH7u4njOyEkEO43cmp0PE9hbEUp/7XKzoyY
Kcpi8uGouV5JQ8n2R/LXKLYGZ0dJ4OhX7lMYRFpC1n1buVnbw0CCIwm737lchpIwdS5tlqCETe6d
ILKNeS3PRu5YJBoTRTZgxXj8fmZQbi6aFeE027jrkTEmRqN2qIkFkAIjgGOrL2NfG544Al1DS6E8
H+8T+yreeX9IzqZHOXpyvloe2ibgtRklwreqAdU9JNX8lETgJncJL0nvHVLDasYG7ReN+Fb8d1bx
/o/w+oUsil1XIdz+pt2tN5rNVpWtazOtRptXvsvYVSfUTPySwiLXcvJ3hAqE+fIv7PqcWecrABvN
I367sdKgEoMq/0NePTLGmdvI95nhvlTWs5ZHJjbCXFU9XC2nE1CTybHt1/kG8u9BAtJp93GenTsT
IfEzcZ8JAncB02z3wxqgMCSXnbmS8Pj6x+xwV3nczK7cwyX+iWlLoVNMOInK8OGR8sA/ATalIlVp
W8uKRutL9Nnn1IF5pRiTPLxdUlopOV9mQxnzF9bX6Wx7bJxbX/BkqHeF/ERK0QggiiYzCYyupg6V
V1mVBcq3yyODzNV4OMmPW+UQtRWc2knYCgb6bkLt6rEhBeLQWs23siSV3FZEZ2A3gCkVNP3t7SGY
WCOq0g6lVjIquYnItQ3rUrra5TUuJTTDsCmptayPQw+bXeog0JboAPwv9sWvCIS3b5aRjelRL6+5
riWjgtggI9WJgqgRDLPTQtaboSPLJwbJZsPsnTpYfoSjAt59z7eK3CXz+6EfLxMmj6dsP8SFqMST
mVzWlBAgP10bxTBrsmlEw4mT4JtahipATF0HOZnmHeeqUubWpLMaN7RETXJKg0RursdGMIIIJ5bW
SFvfN/IZbTmGL15SCU57XOOXnjais0ORyZYLSVJLg0j9XPuO2LjtB3yK8gwY7eTUNHeI7w4PUPG+
NGSJ3yefFc3OX7pi+j+tHxB6+AhmrE11BMVdBdG9x+77wtwC9oUbZHWDAEJRdWHrPQKfS27aiQ+D
DmhoeGiVf62JyK00kayRXYs1nJQ8tn9i5vnYrPjoeXhzSKqlavvnMkcSwongcwTg5EqiwiKY5nwQ
xteDftehyJexYiQ4FfX2ouE/5biQNCh/dqhYX4T1RNSD1ZEklm91CoRfQ0+frHRSprzlCj9DD1s6
mO+CMLxwqNXIDlurLyZBR4JN0jj3nuKaFepJKIKzCZ+LNq2C3jwVdIrlTagRDfGfwFsUrXadpZqA
37ceHjHTDmrMqGPrK7YgTpttsLPBKkBnU1IN6N3MteNVkWcY/ehVXsE8czCWFDVbTdrm6rVtXK/F
4/KrVjg+hkbRgzk7iWTtJ0jOLT4rJTyW0bhZbdVvwFHJAVqvUNs+Gm8P9x+t7SfU5uHf7iqZXj1y
D/dFgZuaPfTBsgTTmtxR/GOo5xhsbHAHOJHCx3Q6NaqiYqL06s21Rbdx7acm9Gacc96u7DdRo9Oe
C7sTvuvvjrFRmFieMd2MdXYQqAL1vU35CcmjKhQBg5NgxgH4qpFYMKwHxXqz0HUVs+CFbkiwfzwt
3stv+h161Bg+JKTjU2dMJsnM9z1nab296NKN3U9KzvaeoOYnVDlKye7HJIHTXrJOurOM4Xq4CCs9
DpVatHbq4YrPkYveczs+oYtrXMEn02KYgU0fOzNwhX/A4Co47OeXTXOfQLY8fcGkhexbuV+d4an9
yqW0hMdr5lyYI/4g+xtZTEvAQHOXK8pZBdH0Y8yV3iEAAEzLuTmZvFmgEoba+smbxV0TXFLjWDFj
5ciHe+4M88bLHiW+fsZk8T2mdlV4R23Y24zIC+7b4FsUoSCIIGlKwAA7R3hFOvA/AKiBPNsJvnqP
1kW/rRBPNqHccTkieAal3eybFTN6hi8zYvYsXslNN3rxSsH8/w50h49IBXuPRMCSgnn+iQEH3dpF
UNo05u+/pyNj6RnUlfbF1WoIaRudIytDYWPll3EBve+O/WYy2by2stzXPcoD7pV/R3qdp0mNLcHF
NkklY4tCKMCHmfs24X9sHk9nUKVlODkEq2MoeR97/VX9EMV6EIn2gK/DOzenM4S/xzaN1vUTff39
JBzulWubQiYWVJZGimf3cK5FLJYhPci+5yaNSoevRHpF0FhxV0ngEB0JfM6AgyS1mCcB45CyTw+M
CA2UG9ooFqwITWXnheZAdLdLLwMSPFa8Va3dDVI1Yo3L6VN2R1iXUOp+XtvRgtGgEFfP4X1XUJkP
G/K51gIuOxL7ExaG+vk9bTkjXTZec9v1ScGTUY/r8rtR8CSyphKyaLAN0sfK22dZApi6ud7toWMW
FlaNWtrdYZ6drijizgzFazuHW7yJbMVtqrk7FHRLxJWqKkLsrffT08xlpx6Y0wVzuIquyKm8j+sI
H14cBSQvYmflzxKJ80xvgqIZ4XqFMzkHv4h6P5Qx5R2ly4HFL3KRWH9xJ/6ce44/Gk3P9tQoGiaZ
FBLchEqVWUXNPXRgi0ZvMbVTPp0+H2rd7gQp/wi6krswDKClFgd9IXL3ruC2RLd774IjJk246u5J
i1C5W7G2bRD7rGS6zRD1fnOUjiFnIHpjNyntCvhtNqsANCnpYrhw4MuptrmSKzyIsLH7zLNv/zzi
u/r+iwummCu3SzRJ6XmdWDE6RaqxWzv+Xq9FEcrjUbPh2TLJMMqnrTdF8xBIgeONYAludwZjiSWk
fFbPe3ZcT19k3qvkCOIo83AsLG0vwe0v07k8POGbdLK0ymhCB2LlzfSoosFhaY5rOK0ReFtXfM5S
txBuoLM3fp/q2bv+js6XTmUHKJ6sToDrRWj5Kab/skIdAx07UYRquQqdbGS1UVjTXE4GACsI06kH
91dDaLFEurjmvFpSlHGrNo+uRvF4U28iuaJ8ZtPDy/0y93VOHfDW5LNJI3p+AffchLyker6+SZIP
1+da6k1nZR/uWZk/AZH1a5BQyP7LV1AZ2aIHlWFkloJfq/rNseDYNibcgnwdKUVE49urty2ghbmG
Gd0yQJJv7Zjyp0CGAbQ1syHd5tTPZQOh/k/NGlE0mce++rXRACLZMAPaCWPmbYF758sH+NAF51SD
Hw5GO+EZJNJOrACzKe7B9lDwYquCxLOy6u5pp7al3RT3NvNl4O5XMHYS6N3VBIFd/I9Pw9wrSx/N
Y16+DXb0O/iwgArDudxqRL9Kc0DXx3E99dx9jDNmfywgZRy6IOT9jMOnqmZpRur3AhxPftjqtPlP
rUgqdv7WZfGCpvUDy2QaV0F70jUrG1w2UnXLm8NCT0WSno12sCRJ8/P8olSscYuTyfUX3Z9ViOwH
iKtQkIhLStrcHmTcVCDtWHj1OxFE+ephb7Lhgwu9NmVFFRO4XtofszHRdDUViwz2e4LWajZJrOc/
AYXq0O6EWNG4WWCdGsodrtpKYKXKUhMzzF3VijIEH2g0gdLRWhoCsc/nFjmyYwPuMbmBZDW8CprQ
9FkuMk4VhgxusgSJZlrLqcjypi216c5PCbzO7xrBeBwJjOHQGYBj8arg7RQ/nVsbAMScGfSPQmi9
lpcDnZ7WzX17+3gUBKE4KqABoVV2ZxRWTDwvB45qKw86NickZvbqkvSREPddnqpBiIlBnAdo9xYJ
R4XOR7BbTFZMWMIegRaL0nNy+ni4pYcbzDv3GOUXT9qbpnPU9u7Xd6Xov0pDB4UQP7l63qAVkUUB
E0b3K9VhyuNUpNqf9ygbPH7UaPJcypOirAfsKj4arMU2VSx/g8+dk/q4ocYBA4Yv3rozR149Y1Xt
Ch2QHnvVp7PgLdo51LMTcRxI26v+FJuViQedZwQWvHrIvaZdvvdc4Ihqf+hwgo5it5ZKewWnCpd3
/IMsQMSwz3QL14wBuzGM4TWdm8HITvW6kjPD6JIWIKQCQzlsLE/St2BFhHmZWkkW+SQ05bKY89TI
9s1UU89hl/VXcZT9SBBhHHCyvRu2l4Vqu8YGvHWrGIp0BIMRkUpUoBbtcgosUWAKtMpxxG4O7kTg
BTHr3vqBj5OxKIPs4yI8ODMnSGQ8KRO93WZzMqi5Sx+x9Gt4qTD6EhDBaEnI97tcX/1vINJ+h7YA
BZXoKWjOlNGmglJq8EydZIztehE6ypOAIfnaoBg+7u0PAlVr7cbFgwYVdJHtMmpXRD8D6zEV5QqB
5ovpbZIbItS+3HMChONrjbCoy9xheIX65XADXNCTSgNVROhPijE08iNzeIBbVxEaCXo8O5VNS6mr
M2m8zYrnAc2uL310s4n4U1AzSCUcnCDIDGibtr+SPCredBUs2Yi0WSXn3eJuxXF+Fq2J2R4WL142
OxX2nks6Ed2/64HND822oYa9IbaGAaDWLRqTUtGy6nkLtw1YC9YuyRhzN61Jc5uCKINDRFZ8zdZ4
BjYHvm7Wf7++WcTfMqC0BQDS9W9rrTPohnv10SNBmYtLRlay6+jG17isckLWWdAAOEA1JzZTgs9k
Wy+yXkgLIPWPd7aAxYTt3dTZrnIiH2bxaM98MvAcX+roheNZGni4edbnq6zu058ZJLaa/Jd0KqQz
sIiCPQuRVab7ZuvE2ls2c/FNwJ6NOUBLyP6AO8pryOlmuHkSimjjKOZnx83C/6NDZBQad9p9j0GS
B6jBYlsIMH435mryfH0ImtDrskPYbE2NWhTCA2z6EzvNs+h8o0FK0Nc5LlTL57S5TI/YNKNN54vd
qKdMmodXzFU/3PeC+i9GfK785pUAc2QwWNAodngwAokGkCFQh4wvfGxGq3hRzb/VIVrWEz/mXhaf
LkrevXsmgOZ0fjpe3leBYXIWP+xLp28SO/q5NfoLCe1eBKWs53E4uGyNSVjaAHByTv/DslJZdsY5
jSz43bgqodoReUsUFDPt5sIybGIVwm5zBR7o3NoWR5mFDgSb3QiOe+pyOKfvA61oHFiHQdW1ITvv
1m6Mh3CC7BLPuNXU7LHr5cLARXEQmb3czXNuF28hxYyzrbe5kuTml23tYpY7kHKoxUkm+wCdluKW
haEzJ2uFHCYXcDNz8KR55wKxoqHB/SxsIKCjNp4F3lmmUH8z8Vl0JdYoWUWTV32OUfaxlIOaHaM5
+IMISOh1AJhQnOwkE5Id96uQXJ1PRh0v/u7me7T60B7kPBqwMVDp9hNnEgc+xfIGnPvf3+TFOWUB
7ybGLac1Q/IpZBU03vjcmhw/ipLWimyY9qY2RlQkDPWnHcfiK0B5Nlp2lkQM1Y/sNxxOzI7MOSiz
vbZbFbBJG7Bo2m2+OPirHdAIIvyiAH9LYz9AVOw5+2P5eZrYgi0iqfRw6DJNemZ3srGLwmDn2R+o
YmD5DDjfYLg+fzwC/wkqokfKzuMMqDFS2uI3y1hfmKY1GetoC+L5GHVJtTlIIHeYA1BWx054vh8p
807GwuYIvcE4pDy9vd/42WI5G3/VG9S80Wd26Q9jIAB4jPsJ3b4Degp9L6KPNjywZbnPr3cmOp9w
XbbTVQoc1+2xyD6vVhQVflPRF2XCGCfaA7sol+Uh4JLFqdlVKJ65QuVZG2xy7RH6+5Y4NFiJlsTG
d+vjpuLr+pguNPYzYQ64keHUXHf1JNGGnfTc8FFzDhHFSmwzVEftgfjCu4eYArReOoDEwMDl4tp3
eioYMA9j5UePMLqPMf472xPOWvrIb+WsL5RP7mNagNJqo+HV4cvTN1c/e0/pp0gJNh41VuGm79yi
GiqEtQF9RAfxdKu+b7LizxgmBTyB0y004uR2ofRRxiwvJZelqPpNtIoUfZFqnEzEDjewGSX3HB4D
TxOaRPTOwjJ1voIjzAGXLkVC5nADOp7NTSCS+LWhgfdoskonIsd/MK77Cis25Tft+BTrmmg74PGi
yXll+WBr+4inGN/lwiPAEZFm+J5QR7KiqhMGiPG1W1rm4nIBHAP03+E0o6hHxzyhAcdu/RPIg83u
ddlTKUAqxgV6CkhF8zMeSR2/kvXGEx0RjC/tCrHcA3v72ugKwccCdo8LGw+4Ki2nkrw0h7MbHyvW
dPDdz1nFLudm2ijmP08F76Neud6kaoG6LEEs/G1Xxa2h6siZous79V1iy5QF/5gfIsB06NV2eAl/
f+Tv34bfSXa9znOCdPojP+tvGIDIfpd82nADxA7BV8s8sy12qwaC6/8INdZodiArdLe6ZuB6iU+f
DxDdyqoRBlwGzrqQ9mHoZL1M+lI+BFy4diwsuaJM4vLD/bQDZHBBvYcCgwnWRtlnORUrm0rESEvi
2OjwB/bQVbE/RFgiPwo+pnJ1I+sFqDQ35g4n7DApN/BoOo4uNTMEyPTtoUOhaJ7v1IPgrOVnIi+/
Z3Jn/PumTNOIBm56sd54Cqh7DXzMMsDgv6CEaG5/Et3yIaSR6tmKGAYtv8XYnBKh0ZzV/8VKayTu
Tk2hD8MMv5Pq1kcmSDnRzFl/8m/qfU98ZP0xolp8Xn3b51EMALFvCCT60ILNkiX6V5keyG26KsTz
zUy4tSa0cROSPJHhSJbbWS9iUGerARgsgYmE4AG/iQVuV6ZvYEFraAcEQGJcQvpfv04IInexD8Q4
ZHtehkjqmOGFX3ufw50cuhaN66iLtksC33/qhaVj/EfMVZIPuIdPQ+Iu8Y3/sVvmgX17+PFcDdPN
EsgjB6334py1PZJ1q+JSeuY4B/njPyHX8BIVUP3ZmdvZdz2x6c+P5U4aeAXfcehuWXlAYToir4SI
3MsRhWl9FQuPchrpxlhjzUgNQwbu77MwPz3S/+gFAkX+UwqtkfFbroATbWJ09fnhTzgwrIeq0gHg
BrXdbR1yeISR9hYQhDgGnrGt6oF7yssqklzMPZ1Kbor/WZAfiCuDPEFmFQLpJrTpJS1MPaqmnZhe
IQBNtH54ly9VP4L1SKR+ESM2A3ksKOYRsjOZRGAOiumJXVekA8jkymS6MxELmGY9xEhKrzqhbckC
a7qUvkDQS+LkQ6qAkFuz4rEvlFBrn+dSSDPTmCp1HWVJ+y7RcOnlCkjKHDTb/kWR8TS7jzQ/xCw2
o+ESHsL2JH6u4PVZDLy/EkYsmKtp1TOKmp6kETh2woU9V9vgNUwdSA0HtYer6hfVFQ+L2v8yFipa
b1ljh+hrQi36TjM3/Hcp9A1GOmvvCywCP9ODeB/No81+cwlz+8iNZGU7wwkoBc7RkBLmkCqlrkND
JEyxhhRCPYf71USVFGNne7dfCTJoy4Jck4oGpBb4o6AEr2rLOb2YQAM6Pe07bHGQtCgTSnIx2bsS
OL+bjhDtPmkDGZQSjeY1RzepJpYZE4V3KBHj6s4NGvXUJ5TgYSRhN4CkMCRSrE9JrzzVpShQEUUV
sbL8NKIWig3copuaoibaY1qerdDfpQBum9FCAjIPd/jWH8CcuTAeA9AEoMf+Qhdt43OebbQMceNp
fKBdTaHydZ7gVlgxXSsYJJ0MvxqajVKHOIUO6WqoHfqMier/8WtW4CjXXo8U2lePKmaqcisGPGWg
KnqvsB6ShceEv5BCM17j5UpmL5oJgyRJFEXl3JCT4nKTuY0a1E7dUJrETWqZMO76TJMwNOAXlmpV
e+NlxmPmVnLv7AngJWrstUskqRwJCqHVXVU+oCIgY4YIY5xumQSu9xZUNmc0BvJT8MBFE1ziOQo8
/igyxdtb6yK7e5qtBMk63sWeiZy6oqobcuIqtPGOGBGzl6P13fRvb+SmH+9Nr2FjOHYsT1fuExQ4
NakYjUEq/iLX1HnhOJZtEVu6dnZ2BDsvaM2v4dsDcG6rrXZ9ugGR2Ms32bc1gHs1w/k8a2d485BN
9CnJFWmWRcxE514yzPGrNKNnpq98FLjuvV/8QVmxpQjtrLb6RWRG8rdT8Wj/hwMmyPf2s83rwkNV
UlxvJOpLLo6Xh9U0+X6qO60xd6InwlAQ8oCFycaqmncaQcjKb9hz8917TfVkEBuh8Fwne4u1TEur
9LDYlWH5WN0pkAgVzS9KcXUYowOt2LPkdQJKCjSqkcA+eu/FUU7ouHHmC5m+AMNBfIsh3xlVm2+v
/wX7gNqNVAS5IRD61DV76OTEutsF59vbOdGUuwwJ/6SijcG8Y2u0AU1Ni3pPwMJG48chP4iGa3l2
xtnNEZub27NAA8q/wclVAT+3NAh/8LEPuj80TWnZaA6Uq1/jXGIn/zISb4J/pCqSecoLnWZoq87f
7Anx1vylrSpQOcFsAqlLJeYw3yvgFhaSz8XA3jKoTbEmFiF9LgAIXOj4wJ3pFIPjHy4oIqnrl0/w
Y/nS0DU191tvobD9H/w3c1mGkn3DZCSaBfMCzTP/VjBfUpGkJLaefym3gG5nN3CZuGz8iLOVSHMU
3jgfxbeJg+P9nh7r+UWpOOLOZGx2lxx4qsn2yOPaykaGPPdwt9azsNYJ9WuqMiSukSRUMWmJg03K
j1cOKn/K4wMIPB3alrP8thui20qTgBaJX8ne3AHhurAt4adqKgMrJ9nN1lzYQvtuUdq+GvU3Z2f+
o9ZTtdF000Fbl/WvcCDCbQt7tBBNurUC+US5wC5s1COt4SP1vvC/6r2Nl6ZUWDtecVZdgZpyFqy7
OD79TEvN6P2Q4PmEWjhcdqvGXEPVAXqT++T9KyPchG5eBhkeRe3BoGL8XG0YH4Y6/+nlxPywmE2E
98nUj+DoIgcHBXuuWRd9GyhSGqX/hP69ICfTJh81JVoGpEoW2I64x8CilhqlbB3sZQ6DNlGFQcdW
LUor/Y7eEENQYr72K1KX21ChPjpiPBZQBdgiZFUo/kc+8XaVALOPZVXbyyHacRMKMfPld0raSHpz
cchgjx/LL0RxQB8EVF6phId4SBwJ+iHlQbwZpE36RsMjhagp5tMXgHRKeX6gzXA4CPUzWDnvTJlm
zo+ZViaYwxNFoHAJio4fMj5USL+okgDBTM9QMiP5fkTQM5IAhuLelT/KmlS3DjInojbr9NEMkzi7
tGJ3yHP3M7m922VXXVJI+muS3jJJJX9w9ArdYjmPKAMU7GSlxmHpGOBdf/aqj6vNOD2zyLF5LwC6
ttMhFWoF2XrpO52qSyWH7EAF19WvjBxU+ptMhCxas5fj0/OATDep0x0vFsrIAmSyWiWPmzAbS6fT
hAtLFu1sy5gA2RV6/xPjyYJY/CXWL+BNgM2B8XMuF//VXQDcMzrNAe5F50F6CSOcSYjU1KECqJOr
CYrc+cw/xfm/NsUNsQFXHTrZNSYFqir1Pif0CrFZM82R7JpRKcGrLkbhPDNFqGFLTz2BxRlS/fuL
FDNmj8toXXq8zCSkn3okKsr/76pekmS+gRyLQpynuf11ZL86as9aj+4Ln4UgndU9ZGdeoiFFGtbc
QPnv1JUBs9Aunr940aGVkaZQ+8YWJpRzYfWiEtE5cn+ShhLtzDnfO5u/8Pl7K0vywQXhijsTCsI2
U4+a7VElxYXolhHQ8i2aJelBk/YGC8vPPnSp8+6gCfFs+chdyrGctXro7q4Kd3OQfAkNbNX8lO1z
T90uCcqfJWQ5ZqFmKH/sPWTvpE1jYYHGFI3JaaAJmCIlNofyg0Gbjajf8n+mtzXivouK0ioEho0x
3SVsH8aLrERe03ZigQaZAUc6cpqe1LEFs75yLVjqJ7ahFgCuXC29vZPIafTg0nSrDj3zfEYnqHVV
k/bN96Qk/tGPlwsKVTrQOuKXBbLGv0eoFGOa7cD02s9GTCf8psVGD7Nb7Cb9FNgtTW6d0KpU1hFv
dkA8CR+zXy0RSJ4Cvivx2fKZsl3BQYV0LmFb2qQ2e7CwOoom8GPkBr2qWD6mPOLyv/Dt/sYfhfqy
dijxV20S3K1apcORp4cL0bGanZbx31n9KWmDq6YTKwW46c0ey3f2qyAlYiy7W1BbS7iMSX+tDZ6G
SFXlbaIAMXt93Dm8xp0OJDlzOA4EX8RH4Qh5cW7YSPSpgm5lXqbxRaqlqnXPkctXTDC9zBWdymBi
Q2SzgtxJwSrNNlaZZ9ssn+qLk1z0p9YeV/U2H7I/XjmbX/21wBEg7dvLP3Oo3FJH3uowOH+qpPXZ
fEd2cuSV87mzb38erTfFBCqxJadLWKa4DhVNPvGSRNyIpg+suq181DiM1fEsnaYp5RmNrSp3o2/h
whmTSVOvPTT0VsScRKLBnlBM32WoXp9t7KXj7ldhYFVfiZ7+g1qnN+8EgBCUoRHy+r6jaJEgJo0w
/wuJpIGoiz8vf4cJhs+PxD0t/SVPaTkaYeFA77YJIk5ro8CD4vypgPEiYk3qs5I+Z04dnXXFaZpQ
ZD8dyheBJ/hV7hSTTA8T2o9+V1PZbKW1hr7lxA260lS8+Z3Rlw3pG84p8vDpG+my/shKYjTDdk8g
Rp1PdXzAj6tsF0EZH7kUWLUufe6v9ZrnsysmKIVh6BH41yxDBqj/lBtpMN9kxllBBFrMQD9snprq
JxktoK80SvIiw+gwn6Vp9NJC7QOAYldUg4MQZUFFR7g1gUto62hniBX8cYgfvedG2VHGjYH7pZPO
1s1Ej8tYkv7bUhV+0WJ0HR2nwjQidXeXx75Nouwb4rAD/RRr7jmT/3UmLn9R/Mgd5Doaik2nEAco
Coup8Xbm7TeNErRUpE1WWwhUacKRZ06Rxw06egUTCgZMKO122F4jePQxIAwqYgi0AvpXFF/B34eU
tZqzuF29rtV5cP4o4glvE+r5Iu8xwkWX62RKC5+Atxymr90g10KcWgq05l+mKN6QEqg7mUv2OwEZ
4pNg1EvIAGBz4X6r0j4XQY5rOgGppZ1UsLhnS6NO/GtWBTIG9Od7HnkK/TeKLTR3Iyz0hMHv50jN
QttibB2o2aYaiXjcNoxPkQIFbjTP01YXpmwXuBan0oNI1k9KsWo2YXRhf0AyFus3qLCeMSUEkeWo
EA2eWeE7Vn8vqKAdjrOOnC8Yova5wMVRWGuH2VrgZBVSb3J+VJR/ZThZevPLBhY439IZ1c2RkBc6
BLHkocJ0cZnloyQDj5yo3I+N0WVEQJLQ4xLQ9bnlc79ukthjPIngcP6RN+k0WgGfY3pW+izpbDlq
mYMnGmF10Dt26pDo5ApLGeyDt2JQWLLhQZoswA9IdnDXKAbvSNI5e7AvQdCvWqMPmET4kuXtwQw3
TXmW3GjI/uyUUtK8HUWoTzB6BGaMQctdp3oMWPI2V3z5BnMX3eKO7+e4rRwq8Ivfy4T2AGoT2sze
HF4v/77x6M14j5hRf8Uf0oIeArYIyFOfctWlbd4eG3XMYDnFBNE630r2/Px58Ow5YNyUZWnC6T6d
MlcJzirC4zNX2JvaUtPY6q0R58wIVq2jC1RWtwNQYSX0jYNsbVRa6W6B1r60fvvpDHioBRxeRZ9j
xKt05dIDmnJgzNOsEJhIyaiHYd58qN57qUjHGgN3MkUXB5MlGKJQbsu/QMGcDYaK2nLKY2cG41TF
oGMi8i8TSXjo8u3HOOjlTXIjbeVBfnzHXOc4204EeuS2jaVbCvx4PVpRN6jPmy/lMU4i77B8K760
b0SrCVCrtjBW4OtrZKlwwA1zniZCWnTlZPrWraRhUPlzZHBP0sRXvu8J6fepQ6Tj0ojyTKvBtoO3
rK8hTj8cZaXh34m7byeoSTryILSSJByaOXWrIJYODDFW7IbrX5pwI19ILIHJq9kjhi7wRcEDNFGQ
CzXwMMEAAj0BN0zE3f8t0Z0XQA1TfqYBmJVqsMVACGBQLGWZbRynaZThOpANMHA2zmw2tI9gj2bk
16sG3BLwpa9LJnGVWlH3U2aoKEpgMCWACO0C9F/V/aENrPvj+q0GfnwgnILTX7kqUeKogXV8jI2p
0ZYIJX1YuwcDHVxEWcsgFN2uzK2qhiiZj3nNFNA7xI4MjHwTpy10WrKjFC/iZ3FGLluNURbn3LA2
3Z39mcVEET/xgZmmeoKDQUxn5CwyHb/4oABUw9LJeGh3nPqIIGHzWCTUo0w/OSRwJw0e0kPz9TqL
wJ/JxdYMqdIoUcOGBfIGKbvJaML/XZmxg/wsXFoszOK/MMXc72axZDLX8Bxh3hb1MAdsRi1qurM+
YTtDxwf0QX07YvNGgc8GRAxATbrI0CozV55L5inBiCKHF9POMHl2YNXZfh7j9WeoS1WLnvhM2j5T
jbzGIgeh3nlvi1Xio+hSs80DXAcKQDtZwTskB6TwnV6NYIkXb3rxiNrc77IW8x1Cvte27qHXJ0K2
YBohXAA2gz5ZDK2tn4TZm4FCM4i9TQTr9aKatbJPjEs7lmqhQlb1Wr8ea/RKwVzTqy99kOac0clE
r/uVhF0GR8z+UqXWwpNBkwS2Vh8io3/oUbzS5JngUrAqZTe2yvb+OKcx1UxdpY8pkkN9fhbrFT4Q
6PkMW+XxLV1jofOeI4cSzPPzTpmr/hdXp2FWfsM6vjLGdpoqzMCobMiIoCRTCv+rZU3SJJTM8+kj
nXjI7eApACAYs+mx6/AKtrJl5kusedWQAeGWNMItu2asm66hDBmbd0L5H4PNyABl0OTIFcHFOMEV
V05MiwTAL+zUpb+rago/9T1rLz2u/deGmo+Hwrj9Z71UXC2Kp6H3x4vsB86dz0B4RfSHx7tNVooZ
gOjEb+vtueYS5LSGX69wpj4G/beglGm5jDFptuhtok9ubrVvrNyjKmF6Eas5p7lTNWGDeROxIqe8
KB07fBh9uw1ebkDLtBI4chLS14hJk4eyW8SmKwyzVYwwttZVy8PGmbSVYTqOX3sZt/WQgQKBCfmb
SfPjzYcfnuyDOEco7+f8ND06ug2IXeoQjRGXGsb/bsZAHA4LjiYtlALRTefOlwmgrD55irSXk0e5
QRDj0Xa2R/J7mv1PlrVDK1FARF3HjUocFrgRAnw/QKLPtNP4i7RQnYkvl7hB1CFqNk8yKNggeL3z
12YAf2zgKHu5k9ZnF9vgXZqo0s1xnZyfU095lajJJ9K+e5UHFsEYzE91ys3fK/Hvf/6a4C5prjqy
bOFquN2zdN2wcrVtRR7jynPMp5IsxqSNJvL7Flg3mhtWdd42gEqJoor7OFWDcxLyseyVP8A93IuF
dLP6YuQl4o0dbbQWgf/uwwndNx6IBct0ssnSZii4UI22ABYflO15iWraG7V91Qa87HtPG5gEfwaj
5XfLxBGeZWUeWqlHYEvx34IK0x0lOzZvmKLowDoylXEMfsRseksSq+A8mAWizb6u6/zolXiUWQ0S
IlY4EentyWpWhmY+u7f2KyLLGp7+a7Vuz2dobdqzCBp06mIcSRhqpKCfPmuHwY72rImsNhlA6Qsa
giL0JpaVpFB6kCTXpYiqrcBztAHhh81km8/Kagbiztqltw0r7wK63RXJ5YE6fN3uWXxW3SS4qRps
mk9WGR9snBND3EZq7qW69h2BxjVzLIAeEFQsEYyiizmcV+pR6mf6qIk1Rtwich4Ha00E61QQv27t
tyx+V6DpGR3VNKljYBQc501Tyd/XwkTXL0YPitK8eHgEqIO253YxBIi6quGWxcxkv8E8eZneuxo9
fDgChCmXOMnMU6hIPfelCObnMCnKyYWmrLQZpDrRjC1oYifjssWUCFdGoM3ykIjy8lkW7YU6uGSE
wWehx6SZkDuI7xDzr8XTzd5l1QwBrTOruB+fHfklBSx2WpsryANbPxPV4tK8JU7FzhNiECu+3Xs6
WIn489xcHUK2nwL4vvPBSHPWCinyGO39ErNM0N35SdbzABKzNQfb2ANGL89vvdbhxzDM8OtfTfzE
vRfoMoL5boneUUG7UX9jOn5fyZpqGlNP6t4jlupbm9IXZYB9uOtapmOrF/fCvvjbGt6+NIFZ/6t9
UKVye+ZC2VRMYnf7FPlue00KHAQ9hlM72XwZnwRhcn3I14CDxIpPPlvBKffb2yPVHMxtqfjCo9v+
iAmXk1HWKRf0bPDa8HZYQu0zwfWok5y9NQ6LwtlsdxUbhfRV+WqV0uAgExR4YfOqcUQbzKo0vB9u
3K7PSin7XjE/9nMTbsdqWSOfSKcA234hJM5SHgNzt397EuM+chIkcknbjSuc7z7IbhvNnGDrH9m5
6Px7z8eFC+s/iTNKsidJV9Z6M/n852X87lV3ymtgbNhmfGPZXvyftoGZiuFonP0ukpFUZEYm7yrf
y4j6kkAsCx1ywdY85KkTLQjC4/sJlMZDa+8c5Cpu7zjujNLBjnT23yElVN5uGUK0QiiUS6NhqSm5
DBx7OTpLvFzDa75KE/FnaVGgxZHTqRZ79/mqWEpUxwJro9/ZpU1+TCo5jKs9J4IHpc99YH9t+upB
/p9AHiv3TlhC1aQFt+R7ATeBaA0lMgpiQANv5VvFmx8zLb9tgBNbLfq91bjU1NlV5FwaGhdtAC+D
zM83nlh7QvVT1lYBQQ/XvfZSZ3uhkVWvMNXFqHPDh+7PmS3JhS/GC3rBt1A9ygS7CXlgLEBFLx6p
nU/9pJI8gHDdFgPx4NyrK6ZBEPCT2UTrFc/5vGUk0ux0oPTV/SaZT5eVLZKv1cfUxgnvbwJf7YOp
A6/QBb3qYS461G5Gk08JWmTKM+dlBeL0DGLMCW8VmuSt36giRkqE1+Tgeep05A0qIPdVlJ2TEiwB
bsJ610mthjq6hlC/atdUUdIFfSxSarLAeFgt5ecUZPkYperS3zlCVYGYCAGeMrBkXxeWYnbOBw9D
HjuCpuFZ8Fw4j5XNnQyvHuqnyAvDn80WbNjDY+KpsHDVXER9KDyt0Zf4HhaQxyNNA7Jk6fmk2u7I
LyhZ+lqme2y3Zo4tkBDpxRwuuLPLge8nq+XcYvTXYt3x2Di3BeEnH0OqgcQHSIFO4tym3lf0Rr0E
Xg93waeAhxIrhDUkj2iV4v9nOu5Ms7nFSA9LmCzAcQn9a8XY0+Kr+nEysQWC0wLvByDbF0J9HiEG
o2lN6n0q1YzKUS0vVL+RmtQiL1YKuDXD1/Sa1Tzezw6H39JecbPMZ1SNE0OHXa3VHE760XcBcFka
aDaAo6m9zQTN1nBRuRmJWZclAAWdvHtNl8yiZBsgCXlfg9QQOvvXQjhQI0T+2o15X7t/gb1evRHX
uJmSq3VqZ5Oiir8jgWPYs0rd0T0PC0mg/INRDsdo40hMfZufw95tDp6l7lNG8N4pDJADbv6Vjk4B
JjP+D96InzK+MMfmTh70FF9HSv9Ecznp7AEnIG3eV7yxddFstzjmAZdhxENOs/XvAbIzq7s0KriH
IjD0Gm/4TsR0EEHGvtVIzDZVvaQHA2KSXX1g0Lw+5rALMSSJ/gPu3HFd305MWUmv8MVHFtxuQmEX
guaLI0YadzjXj/ziNwrqnFWCcT5eZu0yrDrnOL9XUpGZp8peYsXkCkaWv1W+nXVsm0mPgY08J2o3
A/KElt9aabMrPjOLXEHnEinR23H1sev671NGX7c12rPAfLiQ8IvyJBQAwVvdoqq/1jn4zR09RhWT
K9snNCE5MeKElAik5lbLsr7TqC9djPXn/RuitbqEndc0PgUNLWfpUm2tUIFitQv5Q/wVGWT7TT7e
niyOF6NkwhYv2lldOSvkPQvD0n0sjWgJfd4du+o3OqF7Jbvf7NuH2dHupd4TC8az3OVzlhBKcjs3
V9Sx0xj94/225hH3A6X0y3Zv884igPZqOS61XqsCbqDyj7gl/c8ZdqXMYcUpJwN/5CN+Q9t0knyU
19Q+mwY4vg9y3txJClDKrkRLIvG6S8WGvJVd7OoWwtTIP/llS8oIZO/Un4XJ72A5uySdxlay22R0
Up/3vncp3Icl9BCEcuetMIXpmZ78PB/vCCzbVT4J/6jx4dZxNSJmiqyzuei8tykLipb9DOHRLqtW
zi8R6P01XcJFzXcuMGx44HHbf5ok4SVhRut9UlRDEG/dn6fAn+PM0X3UzQ5MgJyNjNzOa8kL68L9
FxU2v2NeVVrpka1ubnW9Qc/dyNYi+SSXnI9XFGpHerRwq8B5ISGjNNGu5HlrEAScutmj3fEbrIj/
kaEG8JKS8k3TYlZOwqESXoGCi0532aYyWIQZrVSr/UyhCIppexyiTrjubpeR/q26BAjjySImkd2/
Sf5yLuHG+lH/b0dD6ZlcKsszaI8PCK4lAPs/6A+cj+VS+7s3dmbq9Vlx8AWNy/AnWggEr5s6yt8d
hiG+pBEfK3bbAs4fdhKyQbdsmBFSgazcsSUDAVMwSolcVbGuNpOPouZICGvnNZZ4fUTio7MZ/Tyu
UuWb1LqjNSHEiMvh+BN/ON+HFCdiObdAqTZpLCjRDU/13pafWNBzL+HeJ7JAOKUzeyubSmUVC35H
bzGHZwumGUZt/QKBgNrcI3G0pnCqGPN8kKAZdOuLYpEJVSzXwApGdIkwii71v62H/4gW6BMzAC5O
JRwZ0mbMmKBKGYEJnqoySBMBC46xJgQGTOdmFCB1GUvVoAQb3T3BRBbcV43UA/nddHZi2jd3vGgf
+O9oGzuIn/ypaZ0x++145HvDP0YaGujy1J8gWs0Adto5mMrEg2WSqAbB6zPQdXNaLp2ynMm+3DI+
0UEOgVGe02WHKCZUk1AbeVvqYUyLK37Dx7xxsdTi6M0MvVx+uAYBUkwVhTtnrV534LeiDWKO+yeJ
3ex+jQfF4UTz38J7m0PlLSl6hyZ3oZfQ0Hi7vf7uq+TeJ4hy/NmtwCA5uXSgrpYqrOp88twniiY3
uFZtekY1gAxI43+k2/ddYnkEcEUOlfwh8i9EhZzHSYiaDPfzu3gEISS1twTjQL7ngRw3+TQMs4xN
73zaG+NL0zqidmTV0SaouBY+U/h3AZkQDpl13G9TBQoaAajiKBj+cvCa5mA3WlXgtheQGoUZgQg1
tgG+5F78dR3JdSf7cflJpNumTQukN3TeieAL8ppllCf97Rw1/EeGYAWXvB4Vm4+7VJYgbxy32Q5z
G9BiaQ+8Mrww6pwIs8ViSZ9gyhiZSTbvpce7O/wiHYFG1wZXm0Bx2l+/GGJ/vFgOn9ltxX8qIg1B
y4FKCNVGhVVEsTT6o09+3iy8TPFQMAAQqMpAxgcVplrdx4BDYxkhMHNos5XWFYCAcWMqP4u8xhIU
u4dcfVY/sdY9rWv6CMDhfXExhBu7zXZvJyy+UUDizqmGrONpLNBxqL+sksc0XtJQZcMb6nv9EIbS
wgLqpVzs5JwdfssEcLkCLTasIjXMM+WHerJJ1XRLTm5PD9pSiR+7lYpNgnI42TMjJm8WHVdSkI82
UNXsOEPcQypNkvNv+tfwAZZoHApNpHTyPAoJD15JAIg4YhlshBUEvwoe96vPbPKPsD/0KvUJeG2j
CiD0mMqI6fDm5ZKU1p0LsM2cUNPXuCv/VtJTSQCKWe879/itTN8RU5+sefl2T3STBwK+7xavkLGx
sM6mpXEWHNax65F3ymyNPra0AVYFhk1lBvS7TiAQdb4nqis+rLSslpTtB6tpSwZgc8VKHAE4GsQ4
aJWkW7NmjXEzb6khBU04e/iyR7J3BqYSqBQZPpjgtiDXn62Ov4HxxdOm7aF6zqqIsunlaENkbA1K
ZFCaBmXMHIwrDo06INaS6hxCR+JF0GXEo9pAJyFaTKGBC8FnxHoPDDklMeGNN0z6W9CyzujBMrFo
Y8Acg8xUf4ArKbXvy+PYYXVRAMOklHrfgv+FPOlHfyv7if9sqfDdHOpfUmMdvbRO5R9j2Od+AT1i
Wc93v/SfgHWQkh4O3tzIIsqRIPa94IKcpEw5flTNd9Dg5JOvMAKxg7VRFdzZVbtmXEeU85RkvBCQ
KyQSvz9SbfMjQKQULgfSACkDuKKudKZK85xYGUbZMWd25IJmtSGF1omuGI2ixwBLYVMbqFngqrB2
3uAEsC/ejazLG84qG/rzX2QeCDf+Pt60IiSWNOLhaCaSJ4EUZD56fa9w2ihINW6JEDqN5oDiNb/t
wO7yWdiwTHiepoGDD7XLRh2Y6uTjvPUEjD0CY+SrXWeGqmfUhf27I7CVaD4PuGx0IVyMV5vCdqlX
CC7kzLjk5oPSPdrd9+1e1+J7b8IgSHBSps1wL40CnqXeoaMYJ/y3d+fF7p0jc7QKGuvgB1/LxS+w
omA9p31D9nXPd/c3EAEN6tW0/00+VhFAlOdlou5tOXy7BWp60LaRUdXkXBbmNYBAoFuivD4ZO/EK
WM3UsA4e/gypwZ6amrHzahOSzcVtGQq6ZcOnfWCLxLVfqE4TAV+pTkSD0MGXECen31CtH8VmrIt4
OoQqKvJM4M8XNXsH7KLHQqnQLMnfY0/a8V6XywRE8pYJ4ti7oleryVWFNqnLOeoD1caW07Xun3GJ
bKqVv0U4d2MCWLLHmRZG68R0uPtsJpFOJp89PvyFDc1XJr2HoKVuAmw3bGnsEaD+IiyWFRV7IPxH
UZF36uHR3awaDDq0GXR38T4RD9RiIisNYQBqPV9TYaE4mLjPkbmOLG4LDVP+TQL8QeMDg/yvupt2
wVQJ/bUG9UzFqwfYyf9fte+fngcwLmdgv/KYOl1Cev+j4/4ty4Y+uOyE3Bm9Wddz0Xf1cPW9LugF
fHt8yjniK0ab5cGCHtZRZVacM9b9JH4P31xAMlVH8Er746kz8voIstYmLxrcUssXnz04Qj7t02vu
5m68wFKKQl+S7gbX5+so6/U1mvRGM5lJ0I+IX7mB6EkPgJ3kBgDixtfLOpR8sybmoE2Cj46qdLO7
zYK46yO4N4UaHsB1CJN4zfI2xJ23ThZpV5sEjarem1jx70HJ3+uym2hi1cGbKiqi8yKzKiOwyF9a
PFYAGBDaqGB9zoIfkV6AByIKcvKDQD1FmHB81sZmO+0LZW94lZoDIXyb8VNe5jsGiYTA4YWQklzX
RG9tnT6T9Pn8PHlVPiX31TQpbdfzka62QELN5Oeof9MKkiJHbBUlY6+QY6sO9QiMiDKNNOhjv7Rg
O/brlQ1WsBI/DS9/cYoynWxLLidptKM8fEoyEwxc9cJkpiMIXndetG4F7jRrbL+wpqiJEXLy73Q0
Kg9n3LP0NXBSJaU3QSzbOIAgKYaIHDwAwoijd2vWuCIa2a7tWNisjSbt49h11GuEF/2e4WR0L7IC
YGXhy87BExXRKGReurwD+D3XzSlt+UeF7rOWBaruVqDL/n/pRanzCYdEpA35ownbI5h6qgjfsnuK
eLS7tzoq751Cjxu2u/IxqZ37KPDYiIjmtGvVsQcL0YvBLXeLXIHzbzedtBZ2j7523ZYC84l52nq+
82BCOyUjNhFPTGF/aCg30IbWp77yyaR2RlohNNBqEXeZ6yoYHmRvZj3F2eMC3aDFS0yWLCC4FuC0
WJc9+2PhbYXljiZvGhtM6gks60HhxYLBvN56Sh4bTCdYBUB/V3FOvaiDizhPM82Ajg571XbuZjEC
Fe5BuTmZvDjef/Z6X/1e2yZHjcxUeLJekusOZNJqbdoxBvD6FH6f8umObSlXE9qO12qe2j8e+iKE
XKIJI9J0TbQ8vzUbaheXCm9N/pSfZB5DOCMWzlUqT5VVm1RPMGrxi9g3zgMd0tmCk1oat/KgYTYD
qDTujgXMjd9irSJhqG89kFFzBWPkQaa8y+bY99F5YmxXWOLzsdgMfCDFgNqUuOZGa2E/kM8Y4GrO
VKkIZqC8oiKUm750KjC5vgt06MDwwPs47xtQAVM8ekcJSBKrRSCErhmZbfP1SnCVwIW/xE14XGCP
4NxPdyiNda95sbVPdi40yaPsWzP7r0kAUYQ/UCRbOW08xbvjNzl9Im4WPVgYsYX24ftd/5pB06ev
+hPIGQ9NGJta+FfkZCFxPVcL5Ofb1zg41XkxxSlUHHPuKbwNrfZ7VR02orX447n+jTscdofahhHc
72nN18qqmcp4PYur3gqgJbBySEMRtY30UJtNZYakQ4tDE78f48iTR1xAfBfrT/3zf9CeZufquraZ
Q6UXNygMd9gMwKNCvOY/lcr8WyErdu/tKs7u9hUNGK4dC02vXZO1xfXre7mGKKPgJLc8+Igjk6+H
B1pM1MNKhVoEIJ7rLvxc5pzPkRcq4vg4bbc0exvKxZDUfX3U+LuFis90Cu3BMDU53j8HDPi4bvor
4OVSczT7ZZ4pLfVicLESqqb6lsBqtW4DhatbOhF9TJWNSWdbrcawPj4v99YHrB/W64V4RxpkUut8
YE482XKNxiY+ZRmHezH5MnLTNyubGyROcvFIZNosaghjwlPP8E9U8elLSuOtzwgohgS5lpvmnsp7
+DYR7VuZgtOPUv+kcz+NvF+s42pAxgKr+5C3GzFxx8KCFhQRtDzCk7oBFz3Z1keAMY38an2dQ65j
6tZe+GjK0ZdC6BYoQOlhxeCid8q3QPkFXrEHQPwt9Kz2d+36B6LbyNk6efxOxaBX6H4KN0++i06k
gnz0n94QiTGpDG2JdByyvFIs11VzlSIcqsoIMd2Fmuq40RgSo0LwhzQ5X1LjsZer3kxRM8+CH2YY
PnhrswMLqyjrANbWD8EycXj0oHhCA4auhb3rxCmytJPS7CB0x2/GcN2aXUfnh4xAZ5+997G0G/dk
NgfbpEEIRsJLco3ZjBYsnDTDgnmTOTWS3gZT6/O4uaPk1mZm0Mw3ugn1dcFFtdCuBW88Ycg72yIJ
43tLAS+r3h5YHiNDnbIJXKFkuzSYkC/fF2C+DyL8GilEAs3B7sZRA6+HNCWQ7uhEAzNydTjr90+G
4qEfGSolol5MhWfUWT+Z63y4uUV0l28mXS5VMFAPYeoD9RSJhmF4CjWqfxNvIyMDRiWLRBHcAiIT
58tHZTIjJFd0MQpDmKwVI+1RKToZeLgBEDZM36UePcPtI0t/wVTEKv3ZqliI3Jjl6tfMf851L4du
Z7yKOWWAtYVAG/2KmEI9s7JtOaoKFoV4cYfFjUwWdlsY2ko0BcPrwg2ilhCtC1DqxUrlEF92B3Yp
mQL4tYcQVXyhfxZheM8y/TgLbzKUSS4yVK/j+Hsu3z97TJq41Uy7KS7jpzm2AG2ErsACJkwoZQwL
Ls90NemK8QvQDrP5r+8RCn+9romKGDH+HgnESAE42osdcFtDwADoZbMwvN+W3gyAaSQ2ElNRUm/4
Ntbb6JXtU3KQRYvD5qza2CK5CyNipknnWdP6xKowpINk0Bju5141HUjK+w2iSbY4CEIt03HAOlO/
XYTGfHITWnArvQkmV/L/rZC45yjZHPjqTYyT35udXFBjSGtG8qe1eSLuoBndWiwF8TIiL+BTVMfl
bfb0AvbVc28CtxELgvpKsQyBN9+Tg8kL7IBGyQLToz7CW3bEmG24lgdMzwNBihViPQbWWz0GQa8C
cC+HdJfUMigKlm/uFUG5pPN+LQk4xCKw7UByZrMbAHGWs+vhGRcXbvRI4xlwRuqsCV9cFGI+KkHM
SgoAPTSt09YAR1hoPhBE7dp7Sv/ESdGheKaQlzpLr4hwr7iwpCaCoSyz7yNSkA9gojG2nYdSwUE+
L0/qC0Lgy9qCo00hbtlKCMHECMtSTp3awIsrQRlQ4J7rH69lZNwPZf7TKLAMVZ+sar7XPqTo+uKu
d6QWzU7pcACnzVWSgDsRmDoPzXlTu/Lzfww5ySwiNXS+QyJYGyKMtHNghE/8oSL9RkvcMry8Rq5e
xxPL80krmHme547Ai/AYfFEzACSwFUimKqQe2H+E0gocQU+xtg9HbaMiniXh0C/E2cMDz7JpHJWX
jVstaLmkoLyJoGc/YTFjhcG7a0Yv/rcFXjX4Sx9EDQsDhQRrJT3RmivrbtzetQzPPlUZMUjmjk4Z
xHa76F5mgfa3FCHIZpHoteEwWrN8kTdnmE+icn8azioMlnCggW5abfZXS3E95kQea0YecvGJu8rp
/0s7mephgzr8oY/53FU/ak1dNP3/bJT/zwACYCxdoquno3MZo1bqc6ouen7uSRhZ4higoJQpfdQa
odvgEZOcLP0iga5OQwt884+xHaafHRocTQUHnf0cMkrFHFPNkrWBgNIBEsLczuFethcL4kjb/SRF
5Lp75JaCAtYNpbPb8ebUxvrwwX2OV/wA1X2nrykwSsf67ly94umFgFgloECmq5+B9In+OZUeQqZi
M+X7+FOHQti6TxafwtmDu4FXvkxk/V/dY2271MYWYzjt49LS9WemFgHvqTuJLbeheSoVLjYnvMsX
tgHhl5Nhy+1dEWZCOj0h/+B0yV+r1MRiwyFOJv5I5Vubv7wqpG4IFg8LsEgunqhABT9UPP1VN2ZT
IOA+WeTi1aI5Z9jeE91DdCoVOAwDPkMz8Ne1izwpVvgfU4osobrqOMF8yFI2J/JzhmM9E1YAHHOw
whKA9OW3hFeljtOoplVQ2SvJo/DPTY+KxSIg/n4CT4YJcKTCxuQtAYfb9IdKIlOT82AQuV+APQFf
UbWb/1N/fgA3vC1wnNzpKqypk2iPGZ9Md9oIdwVnHmt6Yy2VdeMKjIvrWsI4ZLoHiZOotBLWNK3Z
Tpko9pobsA2PQFj27R7qa5U1pkMFJyMM/SzrrT43jKnDtp3PcvDNd2g/v5SKSYm7nXECxRIkcoBV
XJs0DZbk1J4NAquERrY8j036QbuEywE9eyXtpRmyc6idWQrcjdzjWoq7e/LHHW0rhS//AysR8hZk
d778VzVeFQ1ZYFOdGW3iOYgCsQHNvt+YA9QabSFUyHuwBbvoF5H+als2+NwEGFiPiXIx0umFCrvy
O9SSjM68f3I+kw/5SLCMnO8lFhdSFSBGaAXlJxzDHQM57hCFJVMfb4NTG4dW/dyQGQirodXmoXlM
LVNgdEb4/Q/cwd7iwg9A/9iscQ5ozt74pQL3OrD9hhV8qasHbhyNCf1VTUZ6lGgc/nnV7Y6J8cIs
iqy6mjV+odMiC2rLjNkCxUiNbHXzpsbxcSTagsFz/YUqnFCjuaOxKlBU/jTyF4uNkyiOQjpQ7unf
OKJ1RAjj2JTxSjb7jUS4uOGeDiL2oX63vho6o9UhNF096u06LKyf0xD1qNUpBKTM29uFRm3LGB4D
J6613s1+ojHH7DqHYJz9XcXpw3JTsHjkAAOqPtYr+y8Z4wglsUpGD7my1ZsQmGPPwqmW09nXJk2Y
eCgWkf2+JJ5pi86mvfYeAdOMAub+SaF6/tJHrdP6Eb8gW9M9bWE0MpntKQ2MjFBAWkNK7xkjmJrJ
iIB+coJ5gEtM+IfpsozwE7u6ufDiW6ILzyJwAcaBwqAxJFzdQTXz9ivxibLZrh+66KMg1O28FkNL
tKu1mqINGMkDDHHdyQR0S4/VnjwOJyCusYICfYvhi/1rkTGaiSGhFg8JKcCKkMvp1ysYvTMsQV9B
Rdqp7gGKrL3EAUHLBX7E69zGPzRm1yz8MtMN4EfWfLfQ7iMdJV6Fa+dyswBLvs/vmarQcJMl24uo
OUP7/VUI2KO+8YumeyuVZgg8+bbkG4SvkfOVR7RoJri9oMMlLvhsATXfjAAU1nGw6PxIOGmdC4f3
wFL9B85zklsvZA7JlcAYCZy2x49wkKgXEk62VQ0SwqAbtzxO45pTTx90Go1ue1eQwOhFLm/wHyfB
RmQsPT2QVJ++fhusnrHDS+KqFZwLOSDMLxeH8DdGyD/5zzwt6zMe0T9gwXOeGQmEU/dsI7hZMXvC
URQKt0utJ0Scl7DCgJ/19s/z9RvwgEGxvpUz8HNrCbt48uwwWrbVCv2bCdISZ6tGX+dqz+ZKUDHr
oqtTH0ox/+lQ6kyaHv6RzEdUfJAmd7JtrNFsmvu43ZEo6Qw8f3W/bxwXMnbjnZrYcNePb9xBfMdU
PAs2QTNaxDlObYkfJnMkXG26A1tWE5LYEtq6hlZOg+ufLpgtnDkE0dui55x5KShDkSiwglzpiDXK
oUStkeyPR6cmO2OZRKfszko6mw5gzJ/h9WCZKJtKPHX7mKP/Q1Ke47dQBFA7LDWErsAsGOVLDecg
o+Rm6L+cRsX9DJ/Jj9y2oQJWSZzFen0NO0Hj2BJV6DjlWkgCUhyLx2g8skkvCkJQQiByorAFV1Cc
8XnfBCSEZe1G+PspS3oNE/Ry0lfEhlZSdPUBtJ2s8giwm7GD4kGUIRIFFb8dxqqfrkB5YHpmlbj1
50LtAtj243VdUAriSspp6utWgIvcUqoqmJNSoMDSZ1ro9SYiMdh7CgNANHj5kCGI5j/SloMC5wKW
/KHn3sAwOuP4z05NVDP11pkR0fDju/nuFlI/NY+FOPupxlxzQyC4eqA8sb9k8Zgw3hsIuK28jpCd
BfFG02XQl1zVsgyi4mkgosKyi3Vqx8IA2IOX8vXFGE0G37huvEGTjb1ZV1JDBQhWlvfvbf4fwYbC
l9spZrTSG+Gb3MdjY+A4Ae54GqyqgJJJ/b4jn9vignFpmhLvFFzDgHWgnUFT+qd24/dA0/b1lQcL
8S5oUsfxnpRqJ3O2edQksSnN9mOyFTMkeQdA+sxl4VvVxo2IeNlm5MnXdjgUO8nxqeF1GfhAlxd6
y9QRg/wyIbO5a3Uj0LBDDrhp2aVfHnzfV1OrtuW663jJsnXHXGVl/3w82qSRXe6FwnAVv08zf9gM
7CmltkaO5sUZ0SDON/vZUvRZNngnollvNfcBEtaVCxQL7KAu6FtUC+0i5PyRJtHTs43xvKxLWdvz
7s0iAlPbFRg83J6lAyO7xQYqMb3pvKLxFEvFzwLXEOswO22wK5xKBrQdawqWJlAyRMBVHBKQZRgJ
wvuIZzlghXQ6vuv9j49okGOuLcxzQDGnGEwblUMpIfoo8WGHmSGfGB7wrarhWZCmRnZtD3emS6la
NFRYoDZF0s/wWOoAY85McTdDS5JgwVcdcWTjP4fBouZL1vzkiyQwjKMRT+q+1eaG1NkWQ3eNzuCe
3wFNLPlf+DhUNkEZQPo1R2zrZwja+w5PFvY5ERRSXxhlRYeggNPeOcsl1o7qBeaOXEz6CnT1TQwO
kTKIaVUFiijNu4nSIWm3zQTXSCjDpg1wGZD73iKCM0PVQxLZLrEZMiLdAEwY4m4kscqFPLBcAYnF
rhIv0cUnOozGahAgTtlEHDg+gnHKUJ40UdXGyLMqg7duq/vb5FT9y1040xDT6R1EiJyxmfleTKe1
3XkWbAttmcJR0OfF7z0Fm6kHYKzS0vfRtPbuxnKWhTsLopmvb3yCiA1uCIjxHAB3UbDfuABMfP0l
/JYNF2Tunbv7ufbXMWvYzlklkdFRvJsS/jksQVXa+F55zp2nQjW/oBE9YD02XHy2nysTSpPq5Myg
X6R+mymef1HkVTJE+vxpVTvKABVwKJaF4/HV3jQGHD7gzUtSGEv8i925yXsibLv9umoqBEoPLfAp
nQlisM8SpvS3Q2UkKO3qkctph1Rh6SkCajks3DfIc0pU9hGEb6nysgLmbyWlF5p961KuRT07BDjN
yUxlTOQjpnPGVXsxrqoyf5XGmb0a1RozwzN8fMBwHj/EmgU9VOLwg6L1YYFmKBPibCsRJzcQKE36
m9WCmgS2ieVtq8w9HN80apOrpD4L3+IWx6BwgFBwR/uP2sFxF/SW2avCeDH7tp4B5RlO9DR5k4PL
w3IH9EZT1HEDOiiqbAmZbA7Ojf9uW+bL4V9PXms/UqwMfIVBaoVhCInJAwMa3SswvROLedsokhuJ
0S0+6V3NUD5g+k83+lTQ/W0n53vKZ5JgPhRBdu565DiEVwqN0sAa/b2XyuIkgZ1m/RoYeXClMbfn
WRYqyDgWgSYfCVMOjphbdfHnVtFuzAMgI7QSDM2QL+ByNLwuWtjWT84DuW2UvC81FhPVMHhY0L1C
/cWNaksx8UilZRnYK1ViUB6PxsHFtLxK3nXAu01qLvmKALJjuyrfV4XSEj3ElvuAUbK8u2mdBngU
LFYyQsq7jpYRgn8ZzWoEvf4HoXyigLo8lPZlEXvR6jgub5lXMNDyzjmi10+li7rud2ci6J4e2Zkq
Rm5sWTuVXu6f9wi+6buSHCKbYtB8lTnbROX9aF5gyOELKe9Po6x15AFHtCZmIWYpmiDZJjswTH2c
4dAEiuXp3WHzIkQ2ckD4uyGQR1VaOL20omQHPMscAEGUiHYjQV9/DekQ1EgGkFnb+aSc/wMB7Wgy
AfJiIV2MBgd8uYhHMOBk3bPkMWymY0ajeImYB52/bWej9vstoZz7zZ9HEytV6vFwug+3OzqOBoF9
ijAIv9RW+VuueSBnVucwoTjH3Kbv2mBJ6W3zHJ3EvptfO5JRC3RqNDXImin97jHKqW6/jFDfZpbk
R7a/+kDc5HYlyp3b0Y8X88+JNgeK9QTOp8IoXXmKMRKzWhRyO3qjKOiazXGeTyT12mSJ8O0nwWIa
hVkdDdT60/H9Tp0vs2ehB9SKzd4xa6XKz1D87MABRpLLI190gkB2x80Tlst3qpT76ADHKD9SFfN3
6qWzWVTZ2PkRVZfk5p0i0fmvNuPHwGYLYKSkVQBHpmn0CCgvMK/DCS1GLroaS3fB3bW0o3QzC9qr
i0dicHNa/B3nOq1CTOLyGpL/HT8h7MVdo6LBhfQl4Jxs5RpW+ikCsefNk7K1GWGuvs49SK6lKGN3
NT2/4TLcN18Ic00mz+WBPacCEhxqfHVEssyk5RXPODnNhMZuomZ0CKzwbG6kmYzRIby1ZALh7Ae2
Z6BH3qPkAkGub4MygiE/BpeK4ChqcFCqoOEgshW+NLZj4CV2i1gz3Uj19j0XAvPFA0R+sQByJMaS
jzV6ZZyuQEGSxlF9UxqL8Gc7Z5hqa4WEb/mjNZTQ8bDroPNs/sEGzWJaFlEUFEoMXF9QbWiSb1of
/4PkBfSCr1GCQ118z7zHg0FBPfNejORPeBSIAVqxRcdCn61EWDnHOdiD1gE8VqoRQvmt01csVsh2
v2grw3/L6HlGUbk6Yhuen3QMEmzPC1ygnJFVRYfznxT39BTgGltn3ZJ8UQlSdWKogSWOkjPTwbuU
rQpEJZoXg5C51VnsCrHkpOsSkplU8vHyfFYDH9+SUguty5frwveexIfiS8YbAHXZ3xZppO3YmEhC
11uIKX8sXmKZMgt/6AVD/7ODwZ9Cmr1bAxTMcvdblUh8aRX6wbZHy9ikEoqnIIiuxvKGEizUNWc3
T/SUwZnmx1kCSlXWXJjHexnjwU9JLvsSTsgd2nqPt3GiRvFlUVnYO2zs+r7IOtAWtN3AObWYfaE1
5wfOWF4dfJmX5oeZudpu+XUGs4zuwRuuIG3/KM1QKSEAJ+zDboMFywhC6HucwGTl4jakfIqN57GE
FG+nPXo1fPix8jW4M21sSyJVvwwNLLfTV3NX5zVfPRHBCwX/gqlm2Buq9vUWn782UhujG72eKeIL
TKwrutqnYpfWAN7AL3RvMmTt8bthnHxcXu2E51HQUPX73Y7XymoK8h8dnzVKtMO4sdmD3pl3XqRw
Wskpcn6JJ7Cyvv2X2ojykjLGq8hZI7JITR4BYGOsgGf+zhq1xI/+vkSTLgDEdxvp1Vy9kDoGiS9b
exjnTAa7iHEqDkXK4QYOUVkrOB5P0RPjnwIveN57bNzTtWSK0O9PPAu2g+8M+IY8R1nC0yaSSLEi
MUFOCp0WbEC+cmjMgvmXjall5TGvynHKXcQuiE93vXTbYE1uIp33oG2Tqdzrd1SxS0Oi0voxhPHX
JqUDp43I1yWIvn2ndwwWDqKzqyrPApaB3m52x0b2PKSEJSiKNSGgFk5/Duel+eGOA53R0OHQK7Ri
Zjg8WXqrW0zJbqWtC1XCPIHH1COhd8fMhOiCUjqyNuc1oVct+kyd1c6IOUf2eZUxIUknmqF1OmhY
27bPF0odcAvVk/fWZVlJkLj7pKeZpy9KVq+Cq0aWfs74oiAyPwSz1FHdEaTVvYnFUCSM4svRBpjK
rxKV6pEUFYdCRvzmYOTWC8RPWAYNt0xC5mNFHcFn5FEfxdiy9ety7pMCC+jprPN+m5o1D4bQ5yyp
YckzGNFTE53ZufwOn+KBQkZ5aSRxaBcTRVb8D4P5F6E4OI5tPcMnHYhZ6vmd88C2pD386Sa27SJM
tTQespNF4xXrpNhe4hgHqUP4O7yalyuvkE1pdmIBl5KnbstEMTsR4Oop/pASCh1uPOn3sehiKgEI
kLerRiRPrV1t9yX4OUM1UPjeEdxWKY2YoZ3WuOn6gtJRvxug2ENiQPjqUmho146KtKgzXQGzzwGL
dyUS3DB3yQ0DwISFaXugFpWN3yujAwvwfbnw0ODCJ7GIN5Tcd0PZA6Pt6AQrHWE0TnTGQuSyUZ4P
CzXkQEeNqUFlHGM8uKwGglOUDl50JVMo7TAb5yERvPOkSNeuRcfW2dCdYXA9vEdYEXGheLmixwLu
tWfuz/VeVCc41DjY1cPkjB3tzR8fImM9cp/CD8iUQo1iWPSSKtUSBlh1KzpdQVBK1wDhTCJYqf1i
bA/KJgSE/1TpG6NC2RQPEf2MHm0e0SB4nfTdIUTF3XS3WhfOlgspum+8Tk3ZWatM7IDxmeoOrt7S
+Dw0GqA49IRR1bBOC8nAiy7ZQbgmGZo2gMg22FP/tL7hqQbN3j4X2u568DXXKe96arxND8l8ptX2
nrDHCV+EASIUHePK/lHOklbvicCMJD/vdZpYM07qyqzZCb+BoR3tZvKAnZqbhS38xX7vHGerkkqm
eOoq5WyW5wjV4PHPSzRmqv4vBdRqs7Qw5MYVaJzqLsJZrusDoqqPwrfhgQw70+GdS/VroBhtclsb
mpUE+dKhzfHYzSpi1G8OHmeaAyW8KRmpzqD+yNDTpJXbVDS+Vhk7NaXcvR0xP/9r09jqT6DEvOXv
v9MgzPp3ikK2jmQ4teo1WniDDC+FraalVBcZuIMbN5Ot5GqYfIkWyWkA67si99oFtN6EV7BHmv2E
hjt02wzoWdYpby3zzQuqjP0Ob9zfb1gWSPPUv1F8TBD6f2w1rTkYv/ZxA5eZ1N1YKTgZEq5XB6Fd
ysg+dA+fs4udkqkXznS55QnMsjuZ7H7laTxtIdehJ5UW3Wt5HOSugdoDNUcnoVthPd3oDy8vp+pw
gXRNeaIEVOqH3RsxjNtUQwBh3SXQQJ0k7pl+NvE56hQW5yjSiD4NJ0cQ2i+88gv3xtjB+lfntZSA
yuJWpdYL60g1YThfYZoFya/k582orIlFN9YOOfnoTHBrP+lUvT220gMd6iqPYaERIx9JadO3Kwlu
ny0jo2fsWBuBkYsTk4M1gHt04YMn9KPukbsN8Ct5MS/+hOA70BGTS0lIc/eczNQQrlmS9kh2wK0z
FvWzG6FZZIvJCgBxoy09p47VEIbdUPx83h2DfffIQN+0rmxtxDAtYCsH3O+6bZK7NQeWhjjl+hwa
IdUn5V0tjZi43pGBmnmDka51XWRsuHZR08KPPZoc5CoieIkEItJjjII7LSHX7U67twQqQUeBkz9N
B1I5f8IoiV826UD77PNDq9Q8jHSBoKhV4bmPmjOb6Aw/D86zfjzkuJ9dP1QCCngcFHgSkjJ3CjdF
D8gJHIDb8D5NhBqlrItAa6fzS5e21VyR5aRTacvpL7efwkTCfrzDnKZEnUchDY/rtlAJLr0Dq2/+
0CB1t3W1OfD2VtOSP6L1MnZi9Ypyi23OfzD36yuymtedveoXRGAQNt1NeSyZvt9JQlbw0/DJTlgx
gsr+9rFZQ2p623ovI8dn/bXOPIO5M6RcAPP/Yq+JJxpik8ZViHw42qqeen3EEObDUtKZvsNrG1Fn
gbpdwUj01qAMp89R6XxcnJO1vdpC3PlbEFHbN9Oa/AGtqTQ2+w4X/p6Mk+MenlPRqIIWLsmc8aFY
HR0pfVMPHm5rR0T0w/Js52coOcm7M5UQgur9KZ5AbBIenA7KNP90hlRIh4px7YYapmSqVFJd9Knu
fJiDJd5thCX2EgboxwpL9K3JJQICoj0/0ZfbVp0CMNAcCpSFhH86H+RnPwwUjU9zMODezDCFr8xp
R8tlmjxkblSruNTyTrIKHyRCPSx9vBOo5/nFBF9h9OSJgQUF/j3VYn5lD8gs+VAElYMd0lCunMUE
MMHqhES7dQtIuGR/DseaxN8NfAUsqisjCt2AQcsTMLnzLP2fUKECYeLYAeoR5N7XjjDu3yYd3Lvi
8rf/IzJHGp/SG6pLA8ModD5exRifBcPVnUgSPTrtYRtZOFLA7Z/lcqtvJUsPbq7OPhCE7O6I7cYt
mbPCeJ79bzoTsa90Wv/lIEOWcdXlh7NKt6AgBKWfuV1hJ/x0yPGeoIsMeXwUtQz4/rOAwm/6RF2K
f4vOmci5n8b3o8hQ9C8RE1fZpYd6y2h9/HX3j5f3TFbCq49wLN6UlbI0hT5yCHGVyR07VsCn5DLQ
26r76xTqDwaQcQNIDFPVkGTqExA5iOxTaBfhHAQ6lgy8KKs/W+uY+kKxh35TuiKCUEqhCTkKvAJW
zMtXhROMs55nplRtStObowk9daZmcMLpHgiQyTUQhNFgZkRhAO1+tjHHr3qzPnDQLpI4NnaeU96T
0kFfnPfWqCIgr/osGDqHc7/EzQqfKbmLp8Ixgdz8RCLETJiMDZXjVjeYZhoj5ri+8xf/8/tWOYe1
ovfEMTmUhSCwcHRob77wtfxQoxNz9AU6mc+eTDAlIQCCHoOK63fQ+ZZC7oquDseSjtbIMaXc+2UA
RIy0+sUPrZfH1RCgHS8h72IKS/pdOmPJCGF2EgsajPY/naT78H37e51VHYC1fTT/pu0SnjKsoi4W
PBC3dSIh6hRxQnP/oXbiQioolKkYIwjQgzxDtNgkZG6ceTAR7PE1lRM2w5L8lhRkmfDI6cl4C0tG
6I3zi7Dm+8EFcOHviRBJ3nNhdnfLuZM+fe3QPsf3knmUD/o0Iha0pURL/LLtjUxAB3/5378ogsVW
wQjc1EONg2sJyuqC5Hp8K2WTg2FbC5aSJS66anfGYR8TRfPKl7afJ6KyRkiNAa4QkMEYHLg1Fo4N
/xB5cuODD/DiQdeB60+Dx2Yr8bT/ATx13CEztcBAjV4AX9NO6fDWugLXSjtU0kquuw5w3Lf/719D
YTrDcBvXecnF5Ow/1hI3RWT1Sau0nVMKHLlUeJuK34Of0IlMeNKWr5wbMER4YwqumviFu1lf+M00
iHuStU1c2SPHLYT6i0yNJ1eyTccjAhgeHQhs0LjBrCI4f6HznXkz7sv6qiP8UTcY6kazzeBzDYBd
juZwow8ZAVllQ09vMwBJmojbm9ZzZNHhTUSy6zXX9+uGJn2D8q0smXxw9KxpKrOjm92AXVbjHyT2
TlNZ15QM3fRaQYIqAAHUqDYGsJbFt+f17EvF1qhC01PUBoUkZXdTKtQwg3bnX5bl5Ik25Fe9877u
bsG3a7eK7IQS4M0PjqKiTXtx4DUOQhMCNBdMyrSZ103Sj4y1J9hXTqZW+RNTqN2EFvKWm2A5h20O
GBbhR0frwNVt8xPFazvmUEzrlroRZGB6RRPTdELWv4DUR2FW+AHQEeH3KBfApitisIECvf1s3Rou
eiVdj2X/M1u89l3n+xe2EYBwgmafxFs0leqGuQbIKdKhOZ3bdJ7f/APC9Y0YO5xeZ7ajpfKp8e9u
OtpuqvRWOSjqBxIw/MeyM3WemFoSXlxhF7SPkcGroCgsNt+13Qif+aPlzLEoXxFIeNlycAFOm542
b9O1BdM9cIxxUbF9SVj4eQDePLXfxYjfcfbK9/zsI0mLRoief2D//+KBlRbYNf6+xIxPez84ykU4
fYm2D069de9cGuzscpWoLXg2HvKNDGyVEVOi2GTuT5wRwuSFkdum0xW4BoLzekVHhwjqFYPTT0ZT
tzDpnzbl16e1cjA3M1LTeuxdD+PuTSsTkSPT57KOJlJ/ANYAMh9A4JJrDUWYGMX57XoI9L7QMiT+
b1DqaC1eexkco4gXbjK75SgNx9zrcpRwMI9fQwlcJ8CPzG2xdfJvOVV6sDFvjupFvOvnxuPHxPzm
5aLCMZLJgteq2evj6fAiuE9lvg37DRcaoowgkoLP7iqbZpOYEdBvdCxQI+BBOMo1+3eD1BfHrGwd
owx+pI9ScYXWmH7oVcAh8+N95PDzcQrf2xE4YoO3V0jKC61Hn5ab/usaCq+1hronMiUbvvQFMwEJ
oWsKEg8kkVYgMz9Sf8EPMwzQPcORaC1KRudJaIlR4ELdkVV8MDhE7VP+vZRPdQhoiH0mlkImOdxR
Et7GNNWdAFmQsreUq64DI5FqeBQ04gcKVtTNKi2QttMg2wqG1BDR9sULEztGUb0VYOpnvjqIAq9A
RKPN6O4blaOLM7u2w4A2CBzU2pkhoqSweUltWS2dn7AbNwJVmsNs6RB5vDoAiWzZf5b2p6dXauWf
SYfDM9osutaaHGRSp5m3I0/FrepRmNf48iP6aoP8O9buDLAiBbJlQ4W1jttAwhB598eFEJ/g17Bw
DqOJ6EYk67u8JKFcRclfKkgUeEfuoCi0zgHPvAxiBmiWsjU4eoihoYpKfaVVKp24xiIO8FutXjLt
IT1zXP8yI7D6dqdT29mIxRKJRcP63qGAqhfJGs0HJe0m+U8f+1OLigCrL5Dwe7YiBUL+1uQp0lPM
0oQ5LwleQyA3X7IonzLLjurwTfTH2ecUoKlumJ+tWcJ5gtlttX0Pyj/I6Bv2bt1/tuDo3nyY63S5
2W7M1V0Od3PMmfVieHqAPw8CMbPb0q+mDwmlDB/uY8UNjKz3lt9g9rkdqqz0jQRh5CpuWWZ+D/hR
5og7u8z5bU88HwQuCNcQzzfn1/JQA3EjicscrddGVLk7YI7vqy9NhOXggjhFFMOBgNC1rL8wqNXt
az2rqfWBVF/p/eMRIwXTsU9HGJw8EGfjVgCbreFgXzjHKDz9tsZGpr8U+5p68uVeBG2AeXLUYpik
fOkstPr+fqJ/eM1Dsaygfdlle4agTarpFXH9MtSuqMWGE47eWkae01/0HDnAltjs1CK69L4hOmPV
w7F27zspdZ9nXhCmqxkZTSgYE4BwuD+gzRssUoJYKte+QjBHG7f8wtplKhseG7t8lqRs5I36KVYe
PL8nE8zSJ+m6om9GSl5oTeQO4BMNg8lBtSt3Tsy9u6ZKsmry2N2ssxqSgZu91s4LuR9hFOb8YFPq
bl1Avis5Uqv3yypNLpiKRRbm/l+VCYYWg6HKLgHE86zBDcwuQGM5GvgX4bZ09E7yNqt6Uv7CLKav
O6ure/SwI+5GV11pIzpgK6logF2cGTn1jzQtL5EePAy3urS0QrVWNKeHAsURW4qD7g5hbohvGN25
9Rkq+h8vCSEdADqWe5MyvjUvjINYH0cR6gi7wtF/A3f/XcxJPHpdlRfXkPJh+8T56TTksKYtpo8d
+oapuutukFEj/ZJj+r6HyWwZLGuZboLT4sX7Eq1ho8UwUri/77pua4Q2XiB99SjYoWR4iOQSllh2
5wfodyu32ILXtER9pJLGb/p/5C592Rvos138h2dNaeMIX4Dqwr7DUdrxHNIO9sI4WPNqUrRIVAaJ
IQpODL5DB35l5F5LmwR4rpQlhlQwq91ifEqux4Te6sTXfkQqr+rMZI48buzYRZ2N9IGlZDSuAR/q
QlzITufuI63v5BGn9xIfEZkhI08mTstn2WTBMXy/1hLEG1vBhsYe2i+uDef2Rwo0x14QmLTxAtEB
T9db5owJGpPhCA/PCoaqjbRikZNfjFRe6tYnA2bz661N6TicVDembskskrMwzHWzHmAmgLGISBwn
ptP5T/t0tM0VLOVXfHOX3HM6uaIUcLHq55GRSVXx0yVb4IWkLKRUpOmHXCngzI8ctlF1jC9+tBSs
4gq92ukAAuXvVmHTYFhUTCBxlt/Za/gz0SwEb27wMHFMHaUFzoVhb5y/EABM7aUQTTH/vCI8Ezjy
9gnaHresLaKinMtHMxyAPwpk+ZbV2bliJvH/VhIMWpDkzEzKr56HBqf+Y3I2hllv5CiBs6YAsV7m
Skfd9bQ9ULH3K9v+pWVCVzoVwOLp3cRxN1wVvWj78lYhBBQOciGxfzMv6bFjlkO7JePFNjmOftL8
XJKh1q9GIe/GzOU+cDnRpo6SG4qDJAZa4Gc5t9vQN4NnhgilPDghW5ylZC2sq9jVtAPVNzimx/hH
c/xiviSVdVE9xt9TYXBBAu4ViQJOP+TDquj2QyBD3r3215WvGsNYwKX2KGN1YslkEooYbaqYNww3
rVKbGTq1pQke1obh5DQL2Fkr7SPWuOmpgo+vLO/kI8vIgMgdUCvN25+1va1ykYTm0QjWEXlK9Ue6
/Y4EwxiQ+uONazScs6U/ckO4xrrP9/kKulOTV1oEUgowL34nDh+iCSo5Q7hgaZYANN7dN1iaDIZC
mC3NA9wM85dFgfopP00AEmxMs4hIS8XzzmwcVVnb2tpSJsFMZ6nTkCf6c2PyRH3LszpmhgaXlf/k
O/VEHaoMS33LMJT3Ma5txb4nvlO36I6Hxkvv9hsnXYNWXoyc30mqRSuO83YVojZgiX3VtncxRCK9
ZhJZrSB6epXLLg3qaFJLexlEv8i21v4rJC7MTKBSLyknhZOe6ZOhK0sXTEXO03FVGkPt+vzNa2Zz
xbLRtAokaYHH/RKTH20PgWP9j1dqasNwGdRH9eowngC5TKGCXuEnDWR+1Eni+4sIIBaXwou7byj3
v0ONUeUYHvkvIXg0EMcnJgtAyePRowz3IUObCeUYEBh9nZr/vE8QRq8fEJbBO195uLKag/gzM3wR
TH3bm4x0PhRLmpSvYW0PE8CcX/gugOvhMxojjYYQpZOZayKw6uZnTG0UnxC9Cdp1R2sPvKYX9zJk
axfU57snKDE6CAMKcVKIsNIYYw53uXmGcHqPaxCIhOO7vpNs4EKiAP8Zitlzqo1Jv4F7ZwF6ulLx
FabXF4O3y1uYxtbJ5G0FV9cs5SI+VmjLgnIO08WGbzGuIC1JKzxbcfX4bRBKoCztHJ6te762dYgO
QQZ3i2rmjPtyuWNv5m8xZiKu/8DxAYSxEjCjm5s5nwrah+41bwgSC6nx97VH5CfPcXf0b4hcCzMp
RSX3lIgVHa3kPiBUxC8cSWsAvgTAACCmb6wmOjw1nvj3vCfE2WffgUwByiOg/KnJJft5K+z0TC0/
f+blXXXOnVuyOTTQ6w6GEStaXFUBiuHIse1PsxyOGOmr9k5ue2cz55RhT8K7kkz2msSnXEZsgRdq
JqzlDR/wDx6JgfESoKM+4dTv4rDYYqY93t6DgirDgdo4+riGG+xOYP5ygvi+BKaQpY2hS9kF/RkQ
sClnU7vc9+v6bI6TlfucFDgfEGm1l5+JsfepS8yFcUfqIIRzhCcDOz0GjbtRshfVL7CHIPf9yGfq
GKJoIT5BayjfeCl4GvuPXWH3hShgLUVHvwuGIZbWIA8bAupOp1viw5fB6J8CgIwsBzX9tWdEyVTc
PeFTHVQh1vFxkksakvlVVQ+6KK1OM9KIAJSkQsi2tL0KRhy95w8kOGUoor2AxS/wen+PApkY9G8n
KvC31T41BqmbsFFcE7VuBXRqB0iy2PRQNeegXQb7YComyUOLETrWlJlNNq4fRvBAbDeERpDNbtbf
MvCa+MHk3kpgiRjkqcAlC3MbCCegJi2fINDN3DcOIgr1YJBi5scREUV1P7mxhX3+HOmATL58Slw0
PdtkXTzoAfssJKMsaEGeALLGZeYkjGZHwsZb8syj6fWOImXyMm4BFV2raOEHr9wyBcBsFHg/xgll
qhF42R+Y2RVYzARE0hd8+jFIREPMneAIn7T/Ns25lz404hgouM0CmP9UXEbEiC8RchFZbBuAjCCX
LR7fsHVrmxEyYcXT4vgIS5AqD3M0qurPDh0ldoQ/4NnVRmVwDQDb5A3JbEwe6SHhiUsMDpWurfD2
Xao+U214lUMXCfnxV86PYi5/77fh/YWJEmhQ2lzcc0uQf7Yae4rQvBHyofks5W0IwnETAzP73Dwz
G0TBD/y1K3xcQ1AoByL3zX2IDaQnoadGpbCJGgEw9X77Fsr5vHK8jEuVQiuDNEDrQCcFxtuGG+pG
Xrg91xWWKNI/Z/HOc6mH5bMEIQb9driF0WCZRe6NI3/qPpciinV5fJ5pMhRGg1t4OYqfYIKTg2rl
XalXcbVTw2A/u5tz7Z9Nz3BtU+GCfxgY3RowiSCez7GMGRFF0qZmu9xAQ/By1hSWoP+uN+qR0I21
BJYOPgZxn3MZlofe+3eZfHrfkMK6A4r6Rh2q+QQ3OrYG7YXkcbCrTt9tHoCWahTP+GIBsQVO2+Ms
f+/IsEmqRXIIls0ustsibnTAhQiZ8aODZe0znd1Er7OXxOuvsQsQ2K9Dup5Ye77W9zJETwDfkC8f
+BuUYln2vz/seGQElWqJsAvI7V7OdRqCchI6VfvxjtOFNOVO8VaBmW64xYFnsSk1zauGD3mwc+57
Wwm2OQZFzVyhGpGE1NXfUQ0fbR38QLQd+FT1vO+kcjJIruo2pJm/PbOo+zwfWPAP9mggtRlZpHaa
EEDVN3cND0Seq5q2wablpTSbFzUcHF9qrE9zERHi4rZzXzg9dhykYTtyBtuH/22HcTylKbWdrUFl
nJBJrKSEao/ETAZKm8E01UQcER5whVHYe7B5/AEw7pxqN4i7HaU9rOGrqD09x7nDOkV9MzBJX1mO
C/Mh5Es9GtcYIShrgN0bNBS9Z8BKfSCO4x0exU+LH7EN6HObSzWVg3oPyjWq84XLe9ZFlowjnOc4
OFB+KE2+VJiOX9+oDFQo6iUZ+DXmetXyfefpj+M+RR7RXfrdEWknN754FxU78WRTVYL3Lef/z/nP
hNqkR9GympOy2q1n+EH9nmukHMoVVaQs5qAdPZsSnadLTqdffJPbIAh3Q4ly8L15/3Nz35EGoK6M
9vrVsuiNqQbzIKZOhOnwQm2kvY0jGCXzvQM11eMcPoOBo16Bkcb6ewcgF55espNr9qplhJjnnJ+A
1yV8RjWvqLowJUa47B+APK0BiSaVg0v+1ySX2/L0xRoiAEYjb7OChGHTz6EiSYC5z3MT9MwIkwLa
Mx4FFB3pTGcombsyzdor+20ZgUelk5rUeYpEh+53dD4ANZ5WAmrXryBLDp/kGrGntI3wdyMq9awg
1ZTc2mm47gehXXZo3iEu0fJmV4VV55iI4e1PcrhHcLV0kV4TZgkueXcSgflciomIKQFCclKUt1da
WY0I39xgkpZtKPPXhHeRTg32owCqjoOnpdXsf4nMEyBD1it5AzSF6InHBqPLC/JQnaMS2ME8JpDA
mj0ydjlk3KtXHFWWEUNlhXjNtob5aE/FG/Pege1q0FrqppHgKqp2oweozyjRFCJl5RZQg9TnWp+M
Srh7zNCrC72kDYQnQjWGUZWd+xPlskOzUgrFSnRuLcuZm/GI5DsL4vJM63NJ2zYjTr34mnY2z2wz
L5qtlg6xzoy7rUj7qTf4LaONhQ+LKvyjGwCHA67sBx7ucK7IxBAnUjkYv26AoUCx5EsJilWht4wD
Z+ZuEIELlOSVR1RR++Pacq3iXrgZIKYkT4VxVSIEgvyhv/zrjRcDIOwFBRaYZ723PelD2zJJfmAd
JcR7XABB/FYe/fYJp438xrjx3DlMKjkG5xMl26EkyhCYhU9oouIvelhOq06fksCHGRuy0Quc7qFh
IlYZVAogDHQDqgnjaYXTLqhCpc2fo0GUpT0To0cV78aAOz/wdSShkB2Z09vd3mAU7vGqi6zRX+lx
F4fIsnoFLLE+jjL8j2Nb1oVRDpx+xj0OthtTt8dOpoJ9HWsOQNBbW0U5iZYF9i7O6j3BMm+59+lD
AbHQLesklDE8iQ0wZAgS9egHgywFoJ8cGQToRm1haJyEp4FhmHvCMDrJ8rBrIDa7pUE1mAMbJphU
0QHtVOTqweDiS98QrogOP0WHh27YQA7tV7KdsAX6yai4hPfwcaugRYScRLhzMxsc3f+worC/v6S9
kRoex5F0X6fqAN4F96mKBM8T9n4w+w4rgQVKYVSHbK4O9v+dZGnjRHrzmXds+d2NZLeU77+5qEYJ
DdF0976sJinO7P88W6fajdS5p19HEhPz/jV5Vj11UHwqdhJVbjXYH08h171vH/SZOR8j54Z2IJOM
uOjyxmYxoVEqaBDeppYxejslBKSkuGt7VDd/+OaZV60Onxo1hLIPK3xAUPeL6AupJIOi5/AiUuhQ
s5zsvPsQEqUhVHiW4HG6nZ1JtVLVjQuQCFhtrOJAJsZiH1ZpNkIZjsaCU48fuEpf4UkGIS7xetLr
4K/s46tVlNs7os6nhbjQc9HZf/vm5BdmzFmvE1D5Z0ZkzZZHXK9O2PXJ+oDZZxBdnHK9GP5UwJWJ
fuX66lpL4aT7k0sZdhJbCHiRgZUxL525W3MTFZh60Htyq31FPniUsNGtpHMsfitg/y9UEQQTHo9D
eqs/6wyHVT/uWYU3jPyBLMPgHctWo+AZ3lQgkqliKUwGdbA1V/zNFxrzWXo7//ehgq0bX5NTHH9Q
DJKaax7I5+QfCyCKlwK0UX7dM/csRy1DF+GMRF78Vp4WPq6+4gFRQzifAXovkfUstsvvkhPkWNqA
zS4rUaUiEko9v7KdS9+qzN38f7w/nBCWUzBtdJYC213kNChd44w0NCZpsBJhMLiO2TQm6xFWKPwr
caWu6L7MDVu+yNUXyfbIuhbvMJ6TdkZB1tFXBIDlm5Q3cfhFFk87RO/lZNBbOScNhbgmQ8iAMoeQ
FO1BY5c5j4rGGgxdUiQEXfe1Q7gCQIS0NjuCY30ulQwbBY4N7rgHBsC+ekXJTyKP1MOp8hD4oAWs
4MWrtqECnFiVPC7mwv4LTZGAGD/DhQWMwTAleP0hNux4i5gdZuYCBU+KWuVwJyDfGTOXyTAhwuU7
4yfFJzNMd+u4YW54gocfXUSi2eohOO56TMawmRlGPoHyrYQX4/z8DH1TkNh9HYUKqj5EnseR2kUZ
yJ3krjPBs7hxhX4o/4tng8caekZNABGaJPCbSKXsH+Ibr6AUzxnDPOHcNqObp16lg3+XTEtDR4LD
E13IxafAcemhBRR7fz8wOaRgULe1hFC77dc/xXlduF2PnkVu76c1Ry8bfawr8KZaPLojOYel+rHE
q1ay4xvYLUXS6yhnIyS5Gb5I0ZmCge7pBpnQfKJOquPx8Nh3bzu7Im8Rr1LxkfmeOc/byLKGKdnV
sbsjMeySsUMQF+SCZE9HM6rLPe5jnQxMs5Y/VnWG/i0KsTaKF31WQSNuZfF3k95IplkExi20OH4T
dqgWUeXs8Ik9s6WP1tGJfifaZOxrNjsBgz+CrUkmSTEA+fM8cQSOxL54pAdA/yUcwq5sunpEkIWp
Lm6PY8Ke/oHVZBgxPy7gUCB387F3WHKxN0FNYIFN9XZg4BFeYcjYHDcRTOTi+fK+z1mWqhbRY/cg
O5SilkSHeUXaPBRWllVtHPyoRULkmP9P/CcRucYkjH43wA4gzUtr59VVYXVjEqWPog4eQIcnael3
DJEerpMYVjyT78ngeDLSM4vBqa1JiU3WoCRs/ku3JJuxUofCFBtE/JmzF0OV8e+0kquyKRszdb/M
JsQFcp1VChkr8dlWNxTxGv3clZA3LBiSGNLhYfirxPa9WHtVLbmCjuPY6p41bKBN0JV9pLLWWVBY
yNVuCSuBB+AUnL926pyBJBFWBkoSyj6PfPSc9ZkQX270IyXFToxKngFuHJeYNsJGVL9By3gkWa1D
q1wKuv3zqVDlbJFvDKRfwlHCuWUMxcUi7u1L55sfc4y/gBGL70SkDnqfKnW5rrf8+dev7A6cGs8e
LKdgPtibWEMg9SLkwL1L0OQCg96j5UUZTLNoNckVNtbr7abZ/+woPjxm/P+kaLDacl8PRwzD0sV0
IgrBLXJ0qb9un51xZl9USZwbsTyYATKwi1jvzrsEwvkfIUrWrPebipAOrCXZT/xtq/FCvQmFIrEw
eBhAmJKMd0zOTtQrXHd11MP07Yvcx3QhMwcwPLtFNYI27bjge8gpXmXVvWK/n09mpktuE1S5lH0L
Afd6hFEQlZMgt9X3bgUUgv7XLtovjwbeOGiX9nSSyKeGT8tSBfg1a3Y7MpFSqAJIHhvJWvXJw3Nv
9QdI7xGfvod00ETDy8d80WLM+MoTYjc5nLd/bhmRdiRSTz6Otstt/TmktLHZNwsqSEbZSagIs+X3
lronZwzKjDfUz5Bq42aloKQ2Veq85Qh0AiVAoGaVuwrcJXxezw/pHhMSvlG11wg0wqg4KuaNYXM3
vYJvvrlghMoA7djlSfecdB4YqlybbDAUFVRp4CclwUMbH7DftyOdKv7NSO77OLUpq+tsIvPe92GL
FIe0OEAC4SFIwtpt3OOoKKGpE4hqnz54JaFP0CO5duNRp3VTzWyiGEpQDyTXjkShP1Y1Ot4VomKv
D0Ytk6aNMJrPwQZIdkbEVpKDhlrm4zwGxCsUTjZwQbarUoh7xUkybRxAJAfdujVYQlwp0wd1Gm0i
EobHVjoXRSCwC69GfAsdS00jYGycWOW7hQ8vTjNj/uSstimTHxXnlYdjIwh097GHnR51r1o/4HJU
Um5K1Ok2jKLcIzMwWgWgcD7l2CBfawRxVuEg2p16TXY23x12lvB3idRlL25msj+1eLoYX05LqbsX
mj5ukkHWKnWLichM+LH253SEAlCM9Yjg+IxUbeCSw2swddC3lVZ34IrwY3V4gWsuHOugzRkAHu0F
yCCwhyfQ3a/r0drGi+guCQ4G51UsQmNAm0zk2aCLUlLsHDhOlEtg41o4/JQRlXoOYc0JIRKiEs9e
JaceUHs5eDCW95pD+8SmUGmvhMDYiU579ObYmq8/NqCzkOJyHlVIJd2bBzCJLDgQjXCJyZ26RXGR
aiLCOqXz+eVb3LnEhjAFYTY0+xkVQgBBYNdD4hXERk2PDB+KHNjW1HG8bK79wvZOsN90ys1raNdw
vlnVszbacY/oBz+f/sjItuQI+GHMkak2VB9car7jIIMgkTzZkuOdXyC/cwSBCxTEmG4LHocl1d+T
yYbIv/wHB4wg4lkfkZTXbRipaGxQSIKasuHtuO1bTHAaClF8bGYRToycHRPJH94qECYl1d0IMQjC
pvyYgl6NsNM5GMg5WJeSivJl6F1yIXLmlL7KjepfOxFl/xtaou+AK812IqqtoXgL+60AvcmoDKmx
YEya0B0uQd8juS5XbZqq7njJAtk+i899EJi0+uLYs4ZrVRGDm/Ru9lvfrERcZtTMJgCR9FG/OYFj
a/tLD1NkAxmiZb+ARfk4/ynNqcQLLjpGeR+6qx0LEiwt9DFq/cgiQMMD+jscJUY/yg3R5/wZbiBW
9GLebaosahFOklg3Z8FBUk8PNlmH1kMAIWESk+bQHrMNukzEJzYY2eMKYMNXei0vGsEFf8GKsUlI
jyyGbP7VSQhBLpCCSNWRhKTomgViRtpeikuQA3B25BlW3jyqSNI+W87y4rvYMgHoixcL0VExb2oP
GrBJHWKphhkyUgLCQxy4CJWd+VkknFMJTHq0ePqgdzbW15QcBj9xOiyUctGSsUaCQZ4dsMuy8YRU
bVDyF4VIapUiVYt2hXW6nD7AEwS3/XsX4847Qde2gZPnl01fKlU+/Qy+piDiFcLeKWjCVHAwn2eH
GEhzWLfD3GFDw9UIalLTFyBcW5QjpHPvZNVPXCJM3j+rzFokxGyNYQ6VotFXiF1P/mjQhipNsGZW
hJEMJItQL1OWt3z2a699Kjt9Mpa6pSIxFVgyBZoGu1YiL+36tT2SIggc6lnBt7xgUeUr0lZ5zIoS
yc4HgejNonqHgf+e8x1P4XuXtSnWs2KAkEwIRha43d3HnpvwKCoN/dz7k2j8Cqtwd5Up75mzIKZL
MYHflu/r5aJlZ6bieqpeMk0Fxwy7tXp/MktQBsqgDD9l2/1A0G3hkyj3sEjLSE7YDKObYxKzTxC6
Ovrz/xV1gEZMaZ6ki/DHfQL16jVc0xgzN9vZ5SMulBcJQpbw9T86+r+9fClZ+zSON3VoCQOnlHdn
lyC1/L9MFm0LgM1BvVpnLJvohd6Rryl1RhxSk6806RkVf1W+nWJkqQ+xntbnE+dJEVo6kCuUlz0c
PCqewn+zQBDZs9wBKiBHrl2zbKu+jRetu4Q8Aq5uJuaJfuMQbNOTpyP4di4XU87zVsB3SqyXkpbV
iokU8mvNVQRZN+LWPV//YPB00gVbGJa3YmGmvOozYgCvIB65r8URvMqZdhDjClL4Lptdls0kcyhD
6HK0h626JCVwCY2R/zMbUum5fJe227QTn69lTM2rU0HBF0REJlspCECJXpxLNxlUWE2RuYMQ2joO
9P+noc9o39yDXoBl1m5fQXTXI3AshgpGfh7KwZ5w3MbaWpuoEmGH3a2R4tVgz5Nj2Fqa1WlXxN5i
C3RQY9neZS+9HUqlwMehhM1d/Mz23XqY+7y93qoSmuDY5+6m/s6VgT1rT08NFMoF9QqUOjQ5lh1s
B1ivUo+aOQL7TDcFgqwkR9PN3O1z1GyogmqJ8DVWHzCvnWuQ4Rnh1/8JfU/4l0GhoVKx1XUNm3py
UaFxO4kAJIMmpCAe4Nfkq9E9MYHO76TMnoteeiXWtx2nueeFB8+kzaSTKQ2P5N3CYPBgeVpxgage
5zFctSCRTw4jc4PMrerKW9dcr83ayImvQRkDsIzjJBx4oTjcE7iRSubsr7psQ0xEQs39jQk/d/Qw
o+qJUaEey90Q1U76QVn/bB12u1bpSakyrlmYgIWE4BtJGu27C2PgisYplYarUnSrD6oJgD4CFPNk
JsV3KL6wrqjvsPGVMautTjyah9TcSiKr/iz8JJ2Vk4VFNI0Xqpogum5Dw56mRUN7MWvKsAwDkIN8
lU3H/vC0YNG/W3axBIBlBsUQpjPpOrPmKZtVNfGgPuROM2xD7rYXgQ6oGiAeeNnVXReYUKB2m73+
EgjEbnwGv9G+sB5NOjvXcEFxUwCS4vxyrq5j7V4RFSAyMJFq5l4Cg7nuT+i2Ygmld23hmVJPGILR
YDkdwnEI/KipfQf5s/DOfDtyJb57WvZ4byejiDfSVzKvhV+2EXhM9nP4gsg0Zlo89A8QAVV3PWNh
6RrXcmSRRlYd2LTfE7kUEcJBYxLDVRulvYG0O8GtyOoNFW3kG8ftqZaUMIck3hVuDMBxOZ12EbtB
siLfbxj4/5ShbEiUMwW9fsQd+Li7Xa7YmzhaZozb09jRSgXk+QAzN+/YsBc9TvnlIlWZMlGr7RPl
egNlvSoxUpO271maEyjNnfjVVCHyY8EPdwLprGcQqEDQ6iEHVDLIpXPiE3BU2M3EEh4b7KOvFryV
UMbDv9RjbwUco82rrsQkrVUqCyXEpjJmA3eX2fte76GPxBfVkw528i1+uH+SJf0tlEsdpIzB5Z7e
xmg71eEGr2XLnJOaLw9za9Q2CEFROy+dZ/lpi9PWojeW7Kcwu/EAHfo5klUJLvjVJd0UwIDEedLa
UlFAhlfoalAyPo5Fzr0Ej6ZicTWXfOqZBSueWwaFZLKqt8Fp8GuDjuqkRYoe+ZXTpTQ6a7w8UqtQ
rc6arWzRr91fHsoigTduOoB7iWIURwvFnH16se+n+8fyK1nziXwtRaznDUIxTuVZAk+OhCq/YP05
lDkQ5VrrZLLRmuAiH9vTmlqGZEI6DYJiPlSKA+VR/CdghfaNzpvQHmU63da5ZFPdvhmWuaFz30RQ
O28zduRrtqg74n4f14hWX2O/h5mS4yQGL5YLqlUHKazY2KYMJd//kF1/kpMy/Laz2x9SG0AzKRRq
k/0U1t64Sgs01azFd7uP/uq+bAxwmq/hwjitukrLd9BK9JkEJlWw8dy/6LrmpVBPWJA9cWuD4RbL
O6MLkWWpKT0iGGylgnVBXLkoxGnYc3LeUi69eOywfeN4cHr7zvHT8Fw1HDWg42bxtk0FO6zKEbLz
xyf3G76pYkIxv37l5fpHHO61c8BFd2qFjxUUl4aCoKDGuLf1ePfyS9hP/QD/gKtTldpzcDKdcHqQ
Bz3nXWyiOlHdUPzUrd8Yf6lSOxT1eF8HvFHkRLQwptxh6U1ju1RMcrdMnFTPLeLTiKHQOMc6S6JJ
1bk1YIKoKHnEfChZcx79HkCq+Noqjhe91KbCyKL5RM+aOQ1veMadZTVwoBHn0Y4XUFdoNDN9/q94
SK4EYzraKvDirqtU6SXn66f102XT1+vKemSFK3X9jvuoNhO8al09+H6+CcMe7Nm+ZDdEOFCHV5O9
24e9XoWtuhkzStz3N/DTc1PJTdJN5+VZzQXSJHR+F4MmPMVZAMh3ksfgNh4FLJN+1HabJcF7ZamW
rcVCUzgR3/p5PUFUCTXqCGbiS8JOKkbyZABwkiqNz97I0dtFzko7rq3zcSGS4zQnzI7xEVZNziab
WJPfeildFOUJPef7BDLgqb557PSzeF7Rqebf9qhquGK5wpjj84GmuFH1OvU1MvasdwbCgBFJlU3P
RNTpuFAGfuLa1y0tPzU37rzkN4c97UBaDPAVj+p+5M/yWzr+kyfErfPSEnzPLvnjt1l/0FfRccUZ
sS6EaVOvYLx9nGueRa8d4D5UJwkpZLwpNyBr+je3fc5oMeziIgGkwSitqBdB5buY/cJAihQeh8GK
wTzHXmqTMIhwPd2CM81w7GJVj6s1eEOyT85yyyIK5l5M4C37Ol3jszT5KYVsbdycwH4+sZB4CEQC
Ecs3m39aclVLnrlZvMpnm/HmaVSkuRF+6uFoBrDkHNJBV+JLpapWQSRyymAIuTLrjzxRjq+lhVLj
/EIH+paHvQWWd+2qJx8jxIgFnJU++Ie/n/xWdYWUfrAzxUJegN2hs//lD4aS7m+MBsxotoUR/10V
CYR115qg3HhgqgmhDNixGK693dGc88Pnqh8vGZYGMo5tgDOjC1fkl8VN8q/xanguMgSMTJE1Xnow
IEGtwDGEF0kz3CBJsB+x2QzspQsBhEPsDiiVROU/nAEQmt25waOo889iKh5dfZxCMYaz8vKfHBQl
xyZYZekWwOsaIcg20msnQ2VpIodyhyoT26ax/O9Q6g5zN1sYmjMkGx6A4X0ePB+BOAPiIDfavinO
dWTZjb/kNALdGPB87GsN6Cp/N3FFapx29VAzXf6mNoAo4+hTuLfKBzVIk/Q2HfZ0QhH+cdPT6CnG
HxIQU3BKKatPDU9YKzAwGjnn6aka9XzlQFw92D85pJNo7t2jCTJghBfoz9KJgGMXmb09HbSXePtm
q20xQqX4er4poxG+vWAN5uHOcwOa4B6w5JiIwC3VNX3nTokUF6DtJED/jA6BPStiTdjgGvGHRMQq
HamtLwyRk7QvLZ3HIEGzrecf37pRtACDUPA4UMehyyH4T278kDKFZjYTHuTEdqHV0E2EHgj617Cc
1eFFEAIQRIJEYWua42v98Z+XPmgmuiC4zO/GxL3p9NakESwHbN3W2jttdg/pF1AHhgiAenRvdRlo
ZeF0qtrYWJOuUJuAIMPobNleezb14WdoRCma4UXDcx6Xc/4Kpr0NBkjm1irFnzoCXg3Bzb4YFl30
Gvs2vIvUe4AUiDz60QsFAW8DmXm7d33vNbF+ETcPp8SaJQRfYLY91dLvgxI5lQ/3FC0WfiqtOJEn
q5pdMzDQdlHaBZhzveZM+2A6QJz6GPVuZ67T92dLi/cN5BM1Dc0/dQUrq8GP54fUDu/YunZNO33o
S+a2FxnDvziUiZ5OOB4+IIFZJeGcUZQB7ec/Z4HcWBeGIdeh+gojeqgTgWVtUNMUHMHsLCMI3C/n
E7Aq8E/f3PXE2wvXgKiT4/VZcEnt6g4QdA9HfmtSfR8f+Aj5oCu7PUjiR/rKOk3tUSCPCKOsXWxl
sXtG9/namd7ZGQ8bDTGf0/zPGrPeFD/Ucn8pou5+PyJDbNWCfTppWMJ6DAZBCgjIYbT8HtWQauEL
bDVg2s7jwjqQ4du1bveroqJFS2iRea2+3sffqGiF/FfcKwOqjJsl8kEPyYuRHiOGi5Ocpr8YW3XX
617aHWvVblZEtXN4lOGVCjTmfteDR4ZP1BgPD6NlY/X3fGtRIUZ+dVQoQH90usXH90oyd5lFlwyH
HR4BU8ZKb1bVmIt5KqfrJrUGO1a7KVwQPFWT+qIpc/bhKUDMQ4etrgvZ0lQ3ebNDrNXb7uOu4uSH
MEDJd9dYjEW/xjKS2srdMJdGh8ra2pocmN8PdBIs1R76m4YZSrPYnCkzdvt6ky9TyvBUoCMBY7IK
48SrUsl3weHbjTlit0ktlvgtyv2IWjzXNgwb0ngLcET23VgU10R6/tG61GFt5/N7fKT7z5Z7kfFR
kg3SuY2laFPFe0tqT8xInvO3b7JpwYkDYttM4RcKaZ4w/QkeVelb5FeXQ6/85s2V/10zyUs4lBo+
WVaFj0LquI/osyL975cX/gobXSQkv8dqkRlsZmbiiuRt/k+30zDgEr1nECbGPgSyD3dNukjEYZXQ
MzrPtlfDWjdZ0IhT84tUTRCCa/ITE0nIEI17281fbJ49sbj5gZ/OlC2JA0Dm5ORG3wwoE2+Nkn4T
AfRrGBOxKq87ONIunMVZ9U85AWMYvuA0HVg494LKQLz5uSWj8pN0s4FVoLWaLzIx+JxFq3+iF875
pe71TmzNzV5y2YGbHiRNGu0Wve1jDszvY0L7dtqkJCGnKRj4D6TdUo+BqP1IJna9qoqvGYLQd8QJ
4no86hbjUM8Yd7ntB3BwfkbAH4bVAr6+oMnqqLNGCoF5AJ4zhW55AhRIjZw1djsGOKQXJfp4wTmg
oopJahf/WkEDevs0PIm7sAq3SOFI1eVaF44RQNXLWY5uWRtvXmZrp5eRzCLkKYDZ6Dy7R/ZQh8WA
JX7s2tcvtPMdIPCg74/5Pwunqp1pss2ikMBmW2GxaFki9eDKPV4FE8xwRoKi7BFgPK/gHPtp5mrZ
P3jmRbn+6HydvlwJAp7PGoq+ogOpOPRzceUzQEenMOLLSXjIUF6+kOFfd0eBZiG3MSGrUyO4ohgX
go4gxrQFImAh3OYvDhyjPKJGR3u9R9fqFjn7MehbEJkdJokTJTgsqNpWaN9hQ12AaRlF1bqBNSco
46rHxTdmKLL+M7sRLxrqAx2bIiaxHEEJhw1+uDG+3a6WvfIdn2awhy/qYuole2zulwF6xSXoIpXD
vuJnhS4aGjDREca5xSsGU3gUz8qf0CBaca+9soeTW3+vrF+FmlPmedjmXuxCGFG/U+Yq99pPDEsa
78lJdi+RCg6sF8axoNRwKkyVOIiAd6t4ccTpnrA/N6GkQxf6gUSgNapqTEfhb7S6sf2wnF525EZv
PbbdFQ68UOCK3Z/pRFETHWRcDjwkaBDf2yhvfFV4AbwRMg8YwhRBupxucHlEVDsci6HFosGJTSuq
4LE0RcMqCdx9MnUn8WCmirK6MR3J7Djb/G32NmioH6Y7gPUJ++vq61NhxLoevpYnZwG1GGRoFMFQ
a7PkYgvO7SPlhOVUMNaAyHl08BacpV+/OrfT9g37NcUT3SK9S7BLuA22zuaGFVwAU+TG5LvT+JJ5
W32CfPOd+EmDgL80+d7zv6GeBaogHfw6GJ4tpO6ZBy7nhEb/4t6jBD6SYPpJO26JqhJZhNYHrIm/
gJyLPFLwwalpomNJymrJfPf0LzKRm/tEfukqyDn6vORBF3kjb7OQtqo0RHFDoSjTiTdsSGuXhTko
SWWcCiCd97Vb92VADID/RbXVkKh6xdfisHT5+pWfvUH2ErrwRcJwxue+p+SRnV/p33J50VNdZfTf
pp3TiHMU0wxXKNWXJXvljYtVXNnYDjauwkeGzPmZnEhe1wxPe7CYCF9LjSFqzsuzVo+jS4Y2PdST
Srn/mCeJDx6uR6hHvJTGLXwWMVxz9EWyEM7TDJDxit2pYQwf+a2zZ3LLBkGRUdHldjmIS/Y3RCTv
mkKCCIs5xq3sEeKg3SR9DyqfbdUtX4jdAc2oEnFuo7jf/xS6g2LVMTP7/+tRgXOc+xl0XXGdRtM6
W06lh24sMaWD02s/RNIBdeKp8Xt/GA4y4uolskNiqJ4uqXIuUUdDxSFRyyuMoX8+dBjx240761Lg
AwyluQmPzNHoMY7R/LKOzQFc9kBENlc6thgpoC0tx0QeDpJi0Ik1yyIpweTYBYc0gAjF0D4teFCj
hqFX+w+e9xVJ3yln2xOt1YjmtLq4OlfW05Gta4OBQd4yO5cKle8yapkRF1kBZIjVSSWBD2HKUm62
pNugsm/xVcut4ef3zkRvIlhfpSMkwWnGfsR4PMcHESMGOMs50AwQphPtbT66ZWHHDMnXGxNjx6cY
J9JpRD9sw651ZCFdlm4LOXzl5tEaG3Cb9MC1k/BHpqeztbbwO/x0U7IidHcdfhsxRJ4uUxwRsz1b
M6CDB29WhQ40aP62bn1/+y3cMnIYohlrOvBJ5qENdwzz6jMfJNOHtLC628soGo+rYRmZPuMIXpM/
GeplINR0vnRnHil4CB0tZyBgpDQLcgVRXJfkxWY0/ZBPLJAQeuQueXVl6MweTTDdSEdRRfIM8flN
qJTWM5EdtjJtEf1nGbq8hZq2JU6h4zBbShyuzAAEi/W+JWjGtUCSfAep+1ho7iE7eGfbOunFog08
gJMtIv5g/CwwJyoNkc4JhUAPXeyx6bHaVNXZCfMHYNG7JfXHQ2RYh7k+PEW6FRCrb769oAEgVUzp
PMbNVL3mwOpyevBXm1hCDBZAANToka1DxQIH3VlH5YRYrtDMDRCmRo1FNqFEbkIcPUGfQ7rW/JrK
7XDt3KKM0Iq6boMUXeewT4u7JT2ny5zQjO/NJfmxKUv7ZOzhyyCdU9t1P7q1yh9odz7tj+6qGc79
oEUYgP9QzBtTCKqmhfMBF/HcgCjLQgVnFDJr0e6kgBBm3K3uF1ofHiFvXtqFcpSlDtx4WqX8ty7r
1RuGGCpAKXd3/olIu0drR2bIH72RvKRx3IK3IP641dSbiz+eYk7fH6U8Fpax+9lVlKv6bOGBi28O
Fxgt+1ksrQXHWidmStS+kFGW5VoDT8uV+PCXAlywcoTQ5OtWNPMvTy1dC6PuXSJ/N3nKExddats3
xwymk4QbSv7tO1Z13gw/DI0hMz77EtPbIJ9POacJlAc4eTj7ngYzwhstt91/VyeuTZXoqSHRihhG
H+nRMgc0zN10iwNa8dYtJNnDj1BoQvuPPgERSXVwb5oqi6biVLDxClFhlY47yN6R4km05y9FwXFG
rJ2Fh38c49SX2hbW5GnUYEJtXd9awfv0Ss0Chuhos714mVT9/26V+Nah9at+yMU1pabSALfCwuqQ
8gcL7Go6DNsBxK5ptKwDG+hsAim2bor1XInU8mqLxwxzfuRqUoaxKK7eYwX/xR7HFKr3RLD4/FcP
nuOFmRY1Hdo0oiiKTfrMyILN6zaz/X50xEfH4fsItjIp7odY2pkjArxeQXBasCjVtTDSI/CsMeBt
rIWpDd8lA45juLwKB4qdKezLkgNucMjU6jduQDqncDrqZOqieqqlsJnuoiwoD3lgS/lTOaQ468Xj
VoqVyy0OLUlHFWSQD6LNLOU/SN5pb6ppVAv0vwr39qkD3rn3+yxxubOJ49kTg+UKTNzp2KJZzVsA
ICAbt9I4moGbWNDX/Dp3jc91j5iebvN04MeBhGr82wbJPPKD8h26ZmUl2O2fFP4ToOUMTGKKJ+Ow
2Pbsz87McqsG5WjwL4PqgNveRVVzo3Ay+dKd3Dw0N1ZQ6SYR9M+ybXwLvcOXycunwsjskLfpa7dl
Dm3J3Fgn3F2lGSS11foAzwNsp0VfcGZO/DkgTZG1zPhY2BKfedhP98FSysEiISTQfnagjr0C1/rL
VJAm3b6mEDhOdc9Gv8b5Tfj3qGtaRxMXhyiQ45ulMkn6Iw39IGftqzIIAoIwOMyDjBE46wT15w3v
iWhBUpO7z8HvqDXWyvCI68wJ4GR90gUWllsPR9rxjrLhDxlQyGlpGhhD+4TUy/LhHlE5WKbuw1Mi
j49lSLMRkn6qOZVzq7Z6zNjAF7tfjE0FNSHYn+0wTBz6BT21u+Rre7OMgkPRGSZbNt9PLZbhu9Rz
lbLtxCiE8YsuExX6sHirSqTT6T5BOn0s33UR5uS+4LwXF0viuDRuwVvPNucQLwt38btii2umbplA
bGBWxrUUgKa6AsxeWL2rwnjIRvxnEsDhqvSUdfVMMSyYgln+UbGNQ4Sr9MKQsZUYlB+a87ydoStc
Zm1OuHiSZkAlq3vb51CZFb4mmU8OA3UqA2D1aZkaIwiWwb+ONwCmTwV31fkPo2U/uQ11P/9fnFcA
JVqK+ihSl4kNNAxz3vvEUovDwK0IzUGChALUQpD5n1mI7/RmRFbSbXkEq0j/5h2IiEqVY6bc29QN
45pJPUw/J7UrBSb92O7T7iq4s1S/N27LElr66GN2UWKFbxtrdz30zJfo23hTDD2pUoihR6YBZoSn
BnL7zxYVR0XP5Ifo8QVflrwKIs8U3x9wQSPl9/GzE7yCuIyEmG5GOr4r7mJudK7ucUDkPbCMVO7t
fqazUmNsEIfzSmB6qR0pSJpIyNem+BSDmHgJnVuKh2qTy0kea+Fe4Ml/FnmVgyl1bT9NWxPeiQLB
13dJgK3pW65391zi791maW9Q/eVIz61CuPE3rZ0js4S4SnEBOdAWebFpt8sFXAKoBLgBAWI/Dd3y
WqBJHl93cDC89x0IjctL/BMTj5gGdOiD63HggUzjSLw54WMPXDG9ECG96ZfRhv5ctYCwUysTM1U+
wDQYMC5w+f690HrzbCAE4jvI9KaWD5JWw88IOJGkiF7nfLh+x8jiTIZzMcaUt+RTxuwkQxdhk4fa
a9YFXAx+ClUh1LmE9cYkW2kbOuoXLsZ+6GSOvKPf4RAW2+oxUJs1qI/ufPBbewRH0jZ89OtQGAgu
WOPunA1ZtKNMfMT+2z0x3qXDMiG+8VYL+51O4jBV/VeO7/XsEQdEAWW+Mg9rrI4kW/30vqnoubsf
iZ32+xPdcHy7XuW0usZhdu2eIOqdQiHmoZNUeeqIONCtyYF+q5k55zUhUTV8+8lPMs6kiP1MRl35
S/trAl+xnfl/oRRC+IRDoQEpLwKUG3nCpXDNoI8/ngUS5ti4v9wUQXnxL8iJQL8OcWELeIygmffB
XY4+71anRctcCgvlFn+q8jHVxhZijHtMeKSy7+zBRZZBfTgPKg0K39MDeVHJ34wc/794xjJ3Idyq
2NF5vmEp7MfJXe0j8Ut5lDV1nkLHNvajs9Q3cnKeKxozMMiLx+ae21Mn8G1L8ElkxfdhcIwG58PQ
mZz4RJ6k0TanQRyemUyPYqxsMyyc7JvqCMp9cmuvtYicfETnmtVcq9R/TdH8cGESXCymA0dlUng0
t0jsp2PVU3ELggpBHtvHkqeGWL2pyQVngMzPZ64sEWy8r1xuZwz/tCZeTKyxCGFl4vPF0Oysjrn6
8SzaqK35wad93B3h3XQmNCHuC4nmiNlPUGjgqcsd/93vk7XiQbsk7kruvZ9GZftxzVe4WJfvyoFM
8FM+rJSLQqmt+s15u90XsJxyhXSJooqOMYYJvcEBImjOQKf7+ugNHzwTKb5ni427NC8tlx9nmHE3
zlB7gur70BZqr/6JH57SsSatvOgaYCqi/iVTnTe4J5/fI45CCL/XxHXx+lU7eAk4UyDOgMrzQdiT
eC7FWriB9FWaSjlVV1JG402BRO9jvn17y+rtigwQkLXYBYeKlWYaVN0RmDmB+NnFkITRIZX0h/jV
kULJoeYyKXVEX6UbXUY/kQJrNacWHruBFRdZlJQSBJLKFUCHkey0VFmX3UL6mqNlevVPVpUB7dMo
e3vHHR71X6qpELooKysXOwGJu+H+p0oKcFXvwn6i6pA0VKk4lQjtsAEvUleRezTH2vSThIgUu1jK
Z1ZSLTc3WX5akaN+ulmq9Fxa9lZ6gMSDykLyTxeXsTfd1gOyDCScBmz4D08x85li0Zmtmqvl1rA5
fvwqXd9yVTbDDtRdNxBaMDC+9Hqr9pzEvDglLFSJrbuqoKLZDLA/Q9ZLbZw1IaD5THw/RfYYwWAo
x+A6nzcdRPfI2iknpLemEgv/s5qhy0vBRQasQJSDduqgXj2qKbLN7MiLxilHb24VCSRI5JKw5Boe
0Nf3GWv19inGH+7hlr/z++CoPOfDIAXw08YVGtTXKKOP8jn9dAQaxQihrmOuyAfnRcyM2DZeAx1A
QbfX+j/f2Pu/JZLhma7d6i7BIfRfaWpPI4xlv6Xtt2FHmuyFjuNrypdBXzh+UlXRUs4y1afW6jb7
3Jsrs4ZZzHBbAsDNWZ8SKqJLqBMI2KMezXDoNIsafHQWw0CqBnqeAy0Pjy8VmKSLntw0zVw8aFol
Iw8GBJIdO+h+nENUZapbh6cb+U31nypv/rkN4kWHWviZBW8AA5Gz5jJ6X0jV04/Q+qeVH9khMsFf
+BpJxlr/yoYiOKJ4adm/WoFDPgqK0s2ycR7Vz/7YhrNRI6wD6bIGAjzYsbgb/XaToayNj930THND
UfGB7HXFDxKWCAv8tr96Z3U0D5U5TY6xWtOYUuud5B5ZvNgJ/WfuUyVQdNLR270umYh4cqFptD/d
UxYVc8Oa/593rLIBdg1iHjfIdTyECek+RuEr0MZ7PZpZXpejQhwzitGF/SKNJU7tLxun/Wam4V8o
GO44REh1K21BCfmhMJQ53PPaPmWOkEM5OGykTXY/pNII+QYVr084wcgETLNOZiFj9Q/PEuhmXAe2
Hr8na08liyteZ8L4yKuJY7oS7DjEmk4gQ/qAYb8UlnSXYj6ZkgmxhNutukUhrIxt0jAu+/U5icdU
gpsN8J4hmeB8wYP4xaiTa5iH4TRaayEdtOsWO7atmOxRYcGq/arTYiVCaHeB3EnItAamVLKDZct+
fuTYDPfQKXkWfiuE4v2EBjurpOC0VDX8dKheNZTmHg6ZfIqHJ8PaP7j1ieQCqFT8baEFvANoMkMN
OSNGMhr0GptxdP4bk6JmYjTqP99evEX8Ds1tMfZFpmabNuKIbjE9AZ4BaY2gJEr1cxb6u21ebcnw
uSsSOkZUsflVPGpAniwiVkq2k7hrA43igMNpAcSNZgLno1G+TRIdn6Cnuttlk87ndv+voyE6ek3F
YaYaBHjydo6ewby8VoOkHxhzePU/lJYGpmSAqyV7JTDcGlYzp6WJSlquzsj9/wyrGNSabhYsYj4/
YRoSGJhUlV1xoRIpEYv4tuWUqFbOW2fCTwV4x4dlMsl7hHQYoLZQGY9Qlhj0CxExu/YwcabEo9WC
Zurbv8QUIF93euRqRwDlDYY4mioxoBBHAWwft+N/1aiLEGhLSN5pG9SHQFQo9dMRRLKBr3oXecnC
5sgjCBuXhJwP0/LSiC+5vB9MhGGTE2U6n0PZkK8LgA2zbaPqteS9c9xP0MstGqtT4cRNVOFPlSk/
UPtfz5Z+QkCTPnfCRLWxeY74fF5JTS0LdjjoLgDJQzMmUp86FgEwg41c0ObSysdURD1qWeCc5o1A
MHuKR3nvSr0eqDVujkZpQ305eIAS4qzBVxGhmUJ26QfKww0vPCrzzLqWPj3uDZMh5mUEKyqORNQR
csSEwFXM8dFGQKybN8Ckd0DRfP7/wKy2TKefJi0lPfSRn8mC0uoiN66NhZwXy3I95tq/mftbegPa
SmKzYHK5OprozuVaQtgKwK1dxBml/y0QlpxSI3m7Llg6/3eyCFpWiapu0rDJdfLVEe3Q/u4ecqut
Xfzt5llE2GhYb5zqxS9WeoB6HlgxQ72R6kSF3xitasB8zyxB+xh67A1QjSKN034GEKC9BWHUz3GF
BoUu/YjQnTJa5UcYtgT3qcyg7aWW25T7BxmpQvwmByL4sEkS8sGXjs0vaYsW1o3PpmC8QHU+ZrS1
ofdtKYF3vjNsEnvJ8mvC4WtrmT/bH0MofOG91NBlKFnVnEmGCTKK0WpT6aYizLq0Q9r9JIH6l+8X
Vjxpa7KxBZXwaqdR5zK5d9UJqIK3W6jlUwSRy1ctwt4CdHzz72YXFMabn75UW/T5DWO2VJLGkbYu
YrpW/2uaCf8qWrLpSAiJPK0aR4YDo1hkOLFnwf9Xnx8CxH2OLN8L0Wks/e9mSnjd/IPQEeqeec53
xuWO122heNwqxdhJlDzNBpqN4ac7Gu3fg1Fo63b/t5LviYBZ6GDskDTX6Kdj5y0LrFCG6pAAsqj6
SCJ8avbwnRtuRYgWuYIh553xJrgmJQq50Mv9U3TxZksO0jry17M4DWdyxdFKWE99BvNdOKh9EcS0
vTLaqZBPJLNKAhT6js+/SmSGgQNMko9WH5/mmGNQGt399lNlM6Di6m9wvI59gCltDshWhovuffzB
bU6y3z+fGMJkzYae6AyA43/xwPXdQCeE7D77Z9MpPZ0moTzA6T55B5C0epFU7mrENk9kHFUpajy7
T6PzS7WatmlRk5CXVx2B+X3mx4Ubeu29qnTv2e1VM47XPmXKFejn5QMudcZBtbtUqODqprJL+SwT
SFCV1BK3K7mkPEM+WveGZPiirLyNtlH9iDXxlzR/ax9bffa2jLx8uBW9AW8w2hN/Aq1NFNyL08st
yWbOceeqeRcVb2YVO8C9GHcXyP9X2WiQqlhZzacRU4TujOwB2oNDu6ISfetocVQZOiSMc30oC+Px
U0qoRbAOYztpeFR9JtQ2mKbn7Kh/SkBhdPn8NEZJgePmM09KXHSRKFcZyiP/oHDwohwL/3IGtBw+
trF1s/tBC3SzFInQ78fdiLAKeeG5qRfSRwAb+Kc+cdlq7g9PT2Y93y5CV1CGAfkoz/dzQXfYwd6I
fC6sL6dxSwMDsGWS+uVy3JpNf2ZrlAqAIQTDIzbAJLCu6loeV9JN+oGvQ8FhmSCHeRdmg2/hoowH
we5SEBHVdd0EInBz7mdS8LNAqOTQuFGhddPwFcUJUJRVy5MWekUlM+i0+aNA68SO42mx6mhd9S4b
tMK8ZckiODakbpif0l7nsksQClqXma3bWaoYED4+vcuTo6qwIWUKOJjFkox4XRE9Pm587nBLD4Qz
ac30Et7/K049RWQm0Bo0SKAI5lSbpQW8T9HiGre3RNlnc68G6ezPQNRkMU6AUwgWmj263WXnUtjp
iLWH11fSAJSC5V+4G6BfHoKU9TTDruGaQWYMNCXmspG7IaHxhCy8FZBnUVlJVhiwJy9gU0kSQZpU
ByFwCrLKGK4cFnkVyGlHwo0tFaWEu5n6qtkIJQ18pM78TJooyeFu89Q98472Fc9DXiLjKhrxNKYe
7o/OnQ8PPIRPLzGWzyg7CzUORgIZFc6ZIS1igbP3gafmReKQnDudCk4yf2rQnxjNcxxLy3wPO7sN
HyRde0PdVB/LCNSvcRpw+azxNK4hwTeoPwomvg9WUuGrJ8bMGn167DKiUVw9Y5iQHiqXfq/PjJKK
HMcCvTA1lOol7qeqw+f10FMCFq4OAL6F5Rg1htuQ5U9PoCx6eacdxt/3Z0TRodMdMg4SliGImr01
DzKjS7FUPxkN3XSom07HDRmSXT2B7aXv+xwC/vxXvZx5vLM1Ozxv1VKfUridLrkyLtHxqxGfh9xy
F6uJq22w4NqGx1ga2kIQLnGXAdoi+mkS9tmgi8lPyS0e/ZJCbHq1TsWowTDgbPcdaR1T2CJ8l/62
uXg0rZ7rchZFq/ZB/8rwYYj7wUMn9QNlxzAE076gdkw9yfBuWjWyKnGR4MAWp0MRwaqWCdW80Lu6
AGne+i/fEv7duKkFMyMrora1HLf4Vnrg8Om6ByC5JYSdqf37Urz3cEBWjARw4mPf8NWwyBPHIU6c
lPuiHOfEgOc1U9QgnLzNEsmHof/2SXe6Bvr46e9Q4jocn8wjaHkZ5OGyCBir2LexNaSvk3zfHvnp
8qNIMEMHM8RoSplTGdF3pqQhaA0RwfV37Bdt5ZayaAPitcSHQwM/CYDibz+rYLr0YCHZIbX2GNIz
LlFS+YUAGQDIqkaR7fuvGUKt20EWOLsFUEGBV22Ga7SB9VdSYdXZ9hpI67xfQcWtlugPq/6zdMZb
YTPCE6wpEcKvtFrIUAiGquq3TQX29Z4OyoW4KWqLUH2rx1rI6+4+mhXqgYD17PS+1pF/w18UKmiF
d4SS8Q+Wd3i8KPhIE+Ujg4vYksCaSpVaXLZ5t/678uIxF69vq1oPmmLt0MrwoYAC4On1hUfbaxRp
U+yOMgdbktLbkdFQY01iUoYgSN1WV4kzEFnZ/NtgaXdoLmFNbTQEm+nkVdDxXB96tGim6aMuLSGH
Keyxl0bKROmayFC/IgZq0xyZsL4x900iwYH9cDbIm14khBxbvCQjgg5hhktRnkRXSE6Ui27MBCVf
G6PfBtK3arupeAZuT4zc5083Yp2gfkX7mlZFEV9lW5rfepF9v3Hr9mDnMDiKlaqmVi0b8nAMSTxg
5f6p2wPF9wbOnfeHpsSvaTkPB6cM0ruCk9oqgkyHdgQK6/bA8STWSgxRlUWeQL/qMGK/XW2iHsYC
c+bncnBzRl+0b+B+gfHvECA+x9qY9pAr9gOWeqciAGzbWQWrp6ocQ7LTRC4Fl98bz4f4UeBdBwsn
Lc7fmCaBOnODssYJZYwPe2B5oDjkpVySPjN6ylzT/WvVtdzhjGu5Jnd0FtnquvzkPEJRguFpBVX6
ryP3mpu+NlepITJVHn6hW2BeLfjXe2/O/AJKSM/m4GMjWQ8cdHPsQSj6XPPBOJcsLBGA1s2djqXP
ae3F8qXCdpltRyUqBI+wQqYwkV5EMI8trPqd8gPsrx658WQw3UhS02v+y+ohY8+illz6Kt4C0HRG
HP24d3+Ya7q3clyToNDFBryz25y8lnDxQgovYD1MT7UMn9a69NDA7sMfHgRaCPeL8fYwkCmH5Ksn
FCKz5EDw+Z16P7ZWT6kIwZ4uMClUgjammdgpasuKP9azbpIP7e6LsjYSWoiaMGjk9ZGvsyHnWL/4
55iyHzpYwz4TG118nxi8mWPL+yWxDeJ6dMMIhxIU88ZYxo1M9N8LbpCJ6gGNCj+yzpQoz2ehfCTk
7GsFrq2xac2yriX0UayD4tjKlvnZzlGWl6jTkeEM5wsTDxAwdrw9RnYYL24Ppks+DW7FZjsACAZA
ZnBnYM9jJS/y3Q7n34pSIPpyqFbcQ2aJrovjMLGsQcTZi/8STfTGIYj1CNMrJXKNtK6UNJcf2W6T
9LcwovZIoetBfvcTWyUk2BUwbt3I1CIqrwJZiQgWbmHC1xyzvjlbIQgsXvCvqXF6CPHNIsxMXKL3
tzh6g9xwba0whIbbRdzzjDg7KhJRzKl4RKTOkDh0PQ7DldK22VIXO3z25wE/P2kPdWdCYqIPwjPJ
pLR1PKr04/LMt3moYtWHpY77L3zcuj0d43cDIznljsoYJ1wpHY6Reu4jQO/nO011FnSyjRonVEx6
IN0c2hSFvdZDA4YpkxkfSKWCARA3PwwpcybBC+TmJjkdfBZsl48wQ14XGjLrE4EKQ3DSHNGWaxT6
zblQNzTfqZWQem6Ho2qd+5JRQ4J4xG3w0p852Mr1steuIUvtXY1bY8Ql/gn9z3d0Kgam9H8dmofj
woR2Kf+4OcYl86QZ4a2+UktTVfY4HKAPuuY/XuFxNQJg8FCBRl+C8tvoA8vBobaVd8PbkwDPZbGv
C7EA3btgS8bQSTkj1t8Ovd3YXFiYk/b05lgcDvwpq1OGlyGcsAQoDa07kZBai5QydWyDvTuZPgQj
5712G/xYwEE2XoT47wVg73jpXmQ+ty+o0uNJOMaGxEodbi710HnIQRtH80/1VOXLD7dZ1mGHiYBM
yl2r6HN0+1lhY6hkNtfBJ+bJW91Kwr4/IYNoG8lOrRhSv43NF9gLmSwBvfW75uqRQ71PRvX/JU6a
brLJwFmAbafyOzT+RODV4AgHAVqmdYNuVqwps0CmGjm/3elpmonT7oknBaJV3THfSykq58n1rixo
AJBXpQdT6bIc2D79IZUn0OjeTCCXumx4Q7svcB5zy86WkzAepNIe87ENvsjJWjezNT3SxY9F5skl
d0DwcbhSExLDLizrjXzauW3BjYLO/dGWb1CGeXK976SmdM54WD2CRf34SqbaMJLYO5vJ2X4kM5CM
U98YGt/IAwxzEtVkD0oozlgsPJJwJh3NJuXkzfsc4aSyp9EQcWfN26rudzPdf31m15O7LU9ZYlKN
DNciDh9hsvKUuhz+1BJNGQ7qEaDxu03hZRh3jo8I8IYFPRFOEf8xnoh2WIumku//EKOnx2/e88wZ
H11fHFs4O1qBsiV/x1lfCZjfkHbW9KVFkvuiuYg4pWntgRqqD/awj16al6z7zaPolUc109diSUxy
MHFuyxDWVCA3SLMWE4AxLfiMpA9FehT6M4cNInqSVr7lULqmAz+/3tot+VybiequsdAN9UVoIPgL
MID0mKoM3qd4mekSIh1q3HfMTAwlcR8T9+1mh7byoIi2lGUMp6EBW1ShFkL/wxJHdaXjQJDnMqzC
475xrFgOchC5AIme/x05QjkEnH8/t2yRWiDdP2xO/aBmi3tb8mROQ3epTkSo/MY21CbcGvEBl8Wn
orJFR6R/eFpLQoe5UAUzsPe2TjtZTBCilsZgCAvbqT3nn4BKJgBw+bKwrL9LCNcNQQGKKxOmZAJx
2UmlQDFQs1e5NEKslMu0wmhbEg3K6seHzxjH8fr+rNknBkXGCEQUOthC4xOL5WYrQCrR9Rb3R6GF
sS1m8CkvA61FyLKs3rwUjmyk0gHeFsuijfvUlng9UHRnAbRTYkkWR2SWLS7NmSDVYxOK5rQbtbuA
KT0WE2TsYz8VxTCN5Butzy6lFbkYLyckkyAIJgm3qGS8oOaYH3iEkhEJqj1itTRKrhIBDvZzTmFt
ATBLxdORdIWQCD9w8ZN2KGOfNmZ6h6O6uO5hps43s1iLsgB0kw6eyk/x58bFohb8FC76kpVf0AfV
E7ZwBghpRJCfGe6r9bBSM0qeMfNt/Eh4XLQgPoW0oyhtmorHcR8Hur+4A/VAraYsWBiEP+7gyYmg
UhSQUKroLZBcFXBmY/oM7bSzJ/O0+2FC50Y4HRoeCnfJ7aCesU6PUa+kPzTYQT4Fqpfh/Hmh/XyE
iNzjiP5SAJ5xt4VPFTsqls+ouIVSTe0118cgtOM65/bwlhunVJ00vbZD8NfCIWERguvPQptP/Dtn
X7DuoQE54a99rwh3sz1RW5JYfFO7ESU9C0Srn4frQ8blVhfbf8w89uM57kICXVUfBSeK6k203+AB
q2Z3ZnJh+E1+uNsT1pofBH72jgb8ePqFw5KqPizVyy7MuoNjw5VNFC/f2XwS8yOH2klJF6H9lSuO
xRVdPBHQxRr5EmaNf/+MIPSdqoIo19Bne0+k8jjsfIiMtnmVtgGbzNNBTmg02vyi/mYuuqjHdIsq
Y+erikge2a7in3uW3t7Wf0Vw9DJf86DHlE0AhnP1a5K6nZyqj00Lgg+JsqzlREyWaRVzwwXwga5V
YUr+gPssYucj59HjUs6CFHWGJGF/2D2PC1Cp1aoup8NGqh0l9SoeIFHt1snq2B2UnHketrJbO7zu
Xjlqsqb1TtgFNWv4u1jEKOw9mtsYS3SfqydGaLo/k4e50PW8GVKZoTMapss9+WMhasMBAu1c+RKn
QJNPMrosKyELQcr7DtKPN1Nu4QxgYZLeA5D8i5nvFlUjnEB5Gv3YQeL+RTcJ/sq4iNgVupxW1QDj
3Nsp35aJAHPC+Tw10W+Flw+tGWPi2G/SsAxQGjmmzEw+U6qzY0gpskvWs2faIQtcgegdCSXdgtFb
qXTT6jdluHGp2/OSNjBj4qulkmmuBxi+lmG3z0BTGSXn8b/VCoVqZ4SVmY6wqjDB1o82T9TiUUVc
CGnNKq6gayBDA/WcCzmX3IqbYtGHC15kKdyqNV4vjUHAIDGLRE7wvyfT8JMFiVrwLkN1yFolvqfe
aGdYAA3VKQ/sTtNAKTGFWW6afUGsqG8wyFj/jRYtGVqJktKYm2DsTSfwPWionOva2j2g3qkr+pXP
99BdzNwX8EN1go+j5j4XBeIV0AyteXhIqmNrOuk8ONpY0WrWAa9PJtZWiE4Ov2VlMdFI/Honwcw1
pv4M8plFsxSjfa0fH9goQJa4JNog54x4IpKs3B1HB/eHYYqRjsTnFj5sUmxLlH0M24yBIdvsMep3
4UezVuNIeKOC39X0t1W/Yl77XnUJsIvcHQF5wLJrO2KBqRY4Ulx+okMI61LQtPR5G3lFm5uft0fe
t3ytUvEY0Kd0/YxRUZmBibOhHcH2NP5iWT3L5PB0N6IYMStmYHyIg05r/ZmhAhB6an7ml1LPEVjT
4uF8jVXj1Z6OE/QNugO+zHor5pLdB2eRAQs/2HDVPd4OjD9oN0Pc+HwRVFhJalNng//7z61VDS5N
vrxTUaZBgpQF3Jb9FerKUNVr50rOD+8JyayUL4TGml6/6LN2TkaK/bv1eaZyVqUX8phMn6PAj4Vc
hamgvm6IQEbLSPTaW6E/3UUKvFgQDnj0h78qWLrr7bSWpoGyIlsK7LEsKFMs0jGJIDTYLaS8KafX
gu0oqU6sA0mbmPbCLUQCqTjubIRXKhjDCbq4ypBIXAZobmj+pJBUa6sYVpV739S7YCV2L0tOK/D4
X+AkrukIqVaOswvCoJA85micPhJA/Es8C1iE3Zj/JGewCM5NOLdcUMjI26dBvkMAhW/ZoHZ442At
Uv9/C87MwB7oqPO1jMC0ugvAMbBJuVnNomWiT0b6QCobPIVZlYelM4DUmdjG1EvM2aaza/e9JNqE
FLJ5CRGNlpCGIiwpstLkWBt1BS3dmVeXcO1azbHIXCytqX0tEqtziw8ZoEc0tqajNpNH7yomZ/Xf
q/yHVENicj/CV54NB5kI4lxvNXpfRD4AO+EjkubB4yN4lOma4FJvh0pDdAPyedEAIIRO1FxszFKJ
MU1qdxGYnccGqNIF8RMBml0OxurkuqFKbU4EpP+QgYjqRgcy1i2yGX5MIEnEgKO3xUOwd9+d07je
2v8lnH2yIzA91hLJmuCfjsMqBBx/6JexugmLcty5xlL0vNDQ/aoB2OOK7fbsuwJAI40nylQhlr5d
A/woVE83p6yEcvPglfisiU0pMs7vC7ZS3ILobDSXZ4AwxnfLbi84yySiZIeuuUZngmJr/I6Sn8FR
wEyqp+lfnUNkGWmhT2n/386X/lckTn1AdIz46QIespjbKIDP5H10zuOr7GrgVUM2akF3ME2YXVai
mOzcrIF3v6u9O06YUj/GPsXDsNeckNOFAi2hgEN2FyTTckys16OiybrakCDNPkDUIjwX8zWjiV8i
Ubb4XvT905v49m9v2IiWa482mlvK2aTQfL/YqqijSaTu+qetraKP7kHxYluaP2zsiFYcPWZgWVEw
RcHacUCyp2LR4WoD5vazpZGlTdKMP5VyWSEwSjmPXOaCnbPRDSTKYCin7046dHAhhl8OhKGRLZn+
vn5AfExdMUX0n1OU9I19NnIK9cvegpQhyhxQXSA4X8EuKgXs4/F2p19+P5rrL3/510zMOGSd6pKG
kGZcDBMp6sMOd0mHhbXCloBmITCIjeooKpzQqqGbyxorwR0BH2ReS/ZPMoJVzfVda3nrbH5ZIirS
euxLQQ5uPP7DOP/zJ/gZauVrJ8NiJF+dRsi03FJS3mMrU71cUe4FGbU71Q8CegoJWaX9aYkVt/Ly
ZulHwIAN5EhyEs65XAy1h1Ih77R9UQSC9K0O0RepxThOBpCrbpom8/wOKUN5YoQDX29YNje/+jBa
umd+Jj+D76NhngMkEgzCcZoHU6+/GbfPZb1TBO2MovmI8Is+uiyz8Wgz8/WI9F2VWAloINpZLHLY
vqniTtCXciY2fTb6Tj9oGCvnY0bVuvhGxDInjZ8Cs9Y8inV4CiQtgcShfHlBCYMePdtBl2AXqdey
jLz38AIz4R8XbpVbpThMmXp5ZFquOhDBueSmlEAhR0tvHL+nwQp35IkfxXXzkdFt5HRvs/4QWQvy
zyr6BgsqI1lkYtH6vJrW8VmkD1knoy9OEGwI5+ps93KFhm0f1q4tkvvPnq9r7evQ+trTr4mVk9v7
zJ3Tz00OhzSmnG7z5ObYPyuGghMT+zpRO5iAeq4iDCw6LAYgQpd0scNrCwhz2eKV4Zv94m8TSsZM
eUuJt1ddf8dfjT5ZUeZrAZs9EG359QaI6QKsfCnW+OlxD/LEj7eKcgdxTLVB5Q7/X5/X2dzl+/0m
Hra+PwFCxBZO8EjoQGLlzRWCAW8Gz6BgtquH0lIdCK/PiUvaYz1F7fY0mmpZP+dHeFP258IVRolC
dsomN4Pm6ssxmj2uNB7RpqNNJtFWpMfZa+zyvs2DV4DQQQTe2YOlN0SDGF3prhDDbVh45qwcymh4
ANXJZlgvvRCKrhMHAkgq/7d2zYJM7mbba+KfWk2qXI/RukCQX7DRup1WwY0Bn9GjScNpkcpXw6uz
Twpblw0liUkqgOVAFtljHKx9d/H5ZyDCu1oHaQzIIG5Ab/1kPKrd2jmU6SewxHxiKkGls+RpgXNL
CXpWnPjLDU4CA+PXaNmXg2pe24V1l3VB0q5Im0p4WwPMxYEu9teysqKqAnxj2KfZFbMzI1QmwWL8
PKPQUokPi9c3nDTrsxHIAj9gBkpKYnfO17QQDrB8qsRintiLl2tsenk6nb6iqOpdSeu49HgtT930
3xjRT7CAXAb3FkOKiVG5b9vDxjzli1lWzgc6+SylHc41oyiyRi9mnGH/w2rNtuTRQVdtqLVXllPp
aGR4qDl4dcUei+Kj1EexM59qalnqWq1tD0Yqhyv9blyVhY89zQgbr4lSwznD+QxXdSh1LrQxXnd+
8u8KvZ/g9kVmi0Rb90//pmKS1GMOBp5iXmQ17jCxqoTDpD9wKLUARxGtihbcPmu+YXhcGa8nXJBT
KSPnhJpipiPHgGmHweG/ktoYa/gnBlpP84Unj3VmC/PSoGs3iruT7fMNAnqtXG3uy7InXlnjF3DE
vwFitPsv9nIBT9SlAl52sEI7VThnyPkp+79p48fM35c5SBUOXARi6HxjnV+/RbZTpgJxjK9kRjGI
JeA7VtpYmJRoMJBbHInp21U+pGODGy3JryYKl6P4DHxr73u/6k/V11syHt0Go1fQZXyCoSltqh79
d8RX9qRB18PslWc13Rb73/WZBArAgs2IjpGnf8K4P14lThFU8mlLgPzTCpCCNfKjG0/C4v9e9U+Q
DNUxJzSfb2H6J9/dCWX3+InaquerROQQ7v14VePkm0P5OtW3M0d0r+qVyWrfdF6oeHBJbyV6bf/H
9kpdMg0nhmWX0s5QNQ56kg2dz/Md1PezRLQHBTqzms96q1zpqjrBufLoCC3MwvUa2gWRDqGsjAhE
VEoVGev+r7bX8eIdQTlyY4d9FcvWkJ/JmuEk4W+6BguLzSDXPO/XWChmJxANS7F4BmhKPdyqjAF4
oH+VEdhLc8KMc7qMSaxZXTT/pYmvHGNrsAsImEy3aN/Vc8G/hOhquZuSyn/nzkpah8yKPSqdZs5Z
j8JpXTlTOHug+XvVyv5LZBJM40kOsWblHMPKN1yuWBIOCnxvtbqm0+cwQniKGLQQN0oGjaRB9sHw
/Gkb+J71k8hfWJ46upArNyikJf3UPr/xsibav10v+WiQFHUqZlwNIM3lo8YFGBftT9TJarHFdM9U
zXLW2QnuxtbhbwPL+xST0cKkXeFZTZm4RrtvKbVV+RvbehSnv1X4V8X6frIm5MC1Et3o3qm55eut
kum62cddumah5Kd11gKNMe7kOSljfIfDV0xEYZpXOy/gImve+xJqV5I27iZXxO497ss1/IzJWO6N
kvcLRIhWXAlQTjBHJ6+VSqxq9Cw8pkVGNFh7P9izE/tGZ7CD+AFDyFlLQ0k0fWiNqojccoQHPMcb
zAGvyGMlmPLM8dpKkQev1D9jop7Aa9n7wJPlo8k0n8p9qto1znF3mC3QMTsPvvw58mLtyLtE1hF2
QzoiViSlEVzNwHSekvbeEUKHPm1yLlk1rHTyAjYFZC7zsN1xEpkUPWyb08EQkVM8MPh6Na1wb8fg
ftutfRlw/VOkslTTSklq+9cIgir6lQ6lfTatVR2zdNzTVfTBei+cF7BPScF/kZtDwckxupgkrkh/
KMfXkCke8HdXnQBeqQQ3AT3t+nIvqME6lM0tuLIz1MjVCO+vN0kOSQzDHFX1PZk2bltPYf3mvC5u
nowRCNivizxARCZdvN+gLyWzV7S9e2PflfNDhBmg52+90MjqTHIjEHQdF+Z4L6GhRs8fvhx10FWR
xTPJ+qiPU+71dPdRcaCmv8Z6bXvJsWruEEftiPFOQtt1hOXORfgiUHoEPU4T2KAyabB5eTO08QnA
+6ZUXq5gSk/GNJSnXRupU7Fdk+KrI5C/mcnSQ83K/8OO8lhESZm2MC/gyi6PIZOf66+QuGHduMMX
2ihnObHEamsawdlULWKC9ZqF5xPl6srD+Vx6YUoeVLIJWwQjR6FdiMyCMFZmAD8a/OHgUdTzVB2b
jCWSN7/mU61dIYrT04ekZglSXAer/KgfGvyTWhFDvGrLHC2XpPN3iQ2+sjesjrgr1VqNCfDMMASF
yPpyZHaR8AR56wMgpgjU0Wd0QLS8MYTd8hTpLclS3p76xYzJ2C7HMKpMv1lDPNwY9nsHzfDpi0bx
MWMQxdK0LMK49396yXdynJj92oDvouy98WHnAN1ikKly8q3fFvnH0ZXty5PceR8wimvAlp5oEQIX
6XqrPUZprusEsJmZHk57bvV4FFC6fvWffzpqairXSo1I2NGzRzNf4kI8t8sovSfchCj6bm3HaWi4
sPkrtuvI1QsCXeKjP0822wMpMqZUPCjfG5mdihCeS1AiQk8Sr8MFpVxz3btAiTEANqImne/Qg/S5
zg+wKM/1zawY8ErNCX5QWNuV33lfNKjH2xhtYySrxll3Vpefzh7IsdW0LiyOoPmTIbiuTbADwg9L
K8E7D/Va1w3QQiLeMsYo5cW7P05D5KDWxnAVzbbbf3vpZn+gc2AcSXD1P6fld5qJclGTrWKqKQLL
P9rHeQYyRuMp8B5awYl+YAHwLf5kXy2C9pgrBbN44eqxBJqDiY4Nsz87wWv4ESDhgezzTl+nDP44
qjDFNMRlxor8HMQKB7JYcwYA6dHQQVKkNJD3K0kqj43zLZJaG51gFROLEhPLsJ1MTCzVM9B3ghZF
jaD5xf/u0agu3wXc17J0QOr9ABd8Dgs8bMsqx2pkhSUD+rAiRBk+Cd+SAzZbKQwh05PQE1Jwjfxg
k8Fex+azS084ZAgGPNxJkGvx6yQQLY/wZwqWlhPOo7ISodMLf5QKE4S0Pehop3UWBgh4mxiwDpTu
uV1UvDWknF81u7eKYK7vVPBFnHs3GtAGEYxNA9t+TlqrY7epBtP+ER8l4syT7IRBVyWIsrnoHYgu
naOarjw2Lqaw/XXW4wLjrAShquGzVawPvgUT94eD9OwRPf95bbCHRU+0yQYGzHBKeI8dLP3hteWX
TomsU35fJ6WErdLhaZN0sN+wMxiut92FGG9nOs1tmNjWK69mQASKeMU797OLZ+3vWi9gcRw2eT1o
jfLnLbPLT8Dk8eGSFbcUh3onwYUcSPQaOFCf0HWeE4EFbNuelAlUyljFMUFo+tKL03oWIlID0WdD
YeYha80LmiGpXrH4lvU7pPeAyW7cV1fcATzU+qY88WWnAOrNRHYh4okpxeMZnTTr7/nbFsfxWLrF
nUZWoW4nNL4KrsK+huUjinzANEHV4ub3F0RJZTyAiRDtXxMKUgt8+GtQXLv8qqlVY4pBCOZmVHGi
4f6EUEKr9OriK5IGb00bMVe542ulWAPfM9y1XZB2/nJIyLTLy1ogyhJKaSstU7hjqd+x3igLXooW
JoQxh8fS5rtr8pb6QvLaj8yDF8u9fHgts9cHchgOk4yqsR680U5XUYe1ZIG5DASKeCi6m6vO2dl7
qiGN9bxDphdAh7CrKiBlRnrgwpmXxopaRbNrUBey/Ky2LNRgfkiyP8XpwWGVZmGBLIP3Sem9PuXJ
qlI/LhlS2AJDGi1PqSCwLorUlztynFDgmkASzm02vWx+UmFLsXUjBeyZyQURnDWdeH/odu2XQsbx
TA+XybP0UPkqvtHiPXnOtOIKn1axDj/nopoGELOmngZmUhzaihK2eFd3Q3WHnXbmkV4Icxt1kzbT
V5d1aYgrfZjIVJUM3BwwH7U6gU9B/u+DAILGOOvEvG7YqefMlsTS0BefZBnAXTREsfbloriRaLPt
E6Nt1SCWAwuJk+u7GWuM+vTaSsmep3zT3XJwf/YQyVsWqLnxx6i4e50009Q7NLlB18EnNMK+Q6rG
Nl2RUP3yohXkHXoZPqrHGVIuJlVaaE2GwGE8Z4BszXnO3mupzHhvYqaNn545ZS/EttwPIsswBfRA
GCzXDesItevljcnIiRVDdUPZsf7Q5qBocN1bDVwtGRNnxE5ZICgWfZwFjqstn6Y6QNFvoxKiagHw
xZbZvitXZidCy/G4Rwi5KAayJRlZ2+fLldo/+tcH9VXh+YyyVXZpuAYRTJ28VtAI8FIwG6PrageB
UiR4PpPmKId8ZKzpHP4SuGq+WiMfjTOaLJ60zlmg39OCH3xe09olqLzoRECLodM7ue9nUskRbKQT
q0sH9jQXs9KaAW9wxdPYTFU82Mg70XCh4YXvmELdGkW4uIOJlZFPR8tWO2wtti3I73GxataTAQyr
hGLleAbHQcMG4R9HzrZcaRg4vU85XKnBZFCWQjt5QanfNnzmIJjjuD/rtvMLI/Y2msZOl/QV8fG6
RxlhN3YFuSx9EWQK7GUVt11RW2wmwxeYjA3a+Xh+Vh0yUMHmG1lny2BhBKXzzalX7Nwi12Fr4jIg
kv+3Bx+iEGavtWk/WbobWFN63rcm73mUiUVy1WNbMBN7VKDVi9Lnb5yPpw2IJ1jiDGkUtDMpUNvR
WXrGuWWsXPHvnBvsQzjNunMrYFTOAvdNUj9Yn6KFsmL1EYajjlEAvpLx/D7HoaDhltKwYhyaiGM9
31N3w4u1WOQn8EQ9fw7jm4ySoc73gBEEkGtGndnhTCTle15hgzp49xRB71rYtmM83t6keV6scKZw
SmmHRc/oPoV2Xphtt9S1i7DWkqLevXMmMB961KMsU9S2cUgIatevuqyoo8JJ9j6NEquyxFkg5MB+
08EfvZvZEpO2pomZAgYAk807HVlmWFiVkYk60EkSF7PSRJy6KGED7N21bzlJ6dM9qaoW2ZRhcLBx
MZ5knNHYe6MA0Lkfh0LvIAoN25Bmnyud0UDkd1Vy19wSM/41IZZyoAf/exdngTemKw3lkKaiFcza
NX9II7uDtLfq347NZmnK9m+lDYfUrsJ82Ge6H9bXiYlUf/1wIZT26Wc84s5PMZH+KYDoUsw1OqVm
hzmNmUAd3Wh9YOrzIZQyC3O6XjWMMHTsD6eRiU2rx0fzzydbgpMU97pbHWSHRUJMsaSPqrc28A/y
lA+gW6/K1Yy6LRafDTrwMPTNhirEyEmdnijZwxLMAgP+7TkCz1SJ6ddmdsYQFIahcEyA0kMxSTr2
RF9TgfuB1YQzWk/uXNaeHXWFoDZbncCBtEx/6xafgU5OjVXOG3QTlNllfjN651BAwBV+vTBrfa38
2LiGKODEyhB/MfFaIkOkbg0gvcMT75caeJHty9IMWAyCQFb1A7JXNH2v4XX1ZCGHoIKZSlc/irm+
s1UNzfFiufAPMxHUtkOWkp94J+yqCTyvVJ1d92ZvoojJhPhfZcEqyLRwx+MiEiQ9y59oVa4Syhcs
yq2cO2zdZoxUqePZwqL7k/r8dZbtiqB9iB6tRlXz6lfW+CFIHunXYE3mGmmqkEQS9WQG8M9IW2+p
zD8h4zAh9krMYHZz+fPbS45WX7ih2vQ5IEESwjyBoCUg3KJ0teyuIUDpX2JZlnHCJyTSXtkLfpm8
e18IGyqQfvAUjVHYThyu1mPYqNJQJdKqrSi50pqyH202bqO8IjQ2PMmNWF9fAm9QtYXX6WV/AMqr
6TVBx4wtm//22AHchog145l6nGpTO95V8JlQopfK/6275AT5dLKRIqlrzziDGhwBhUZaYQCLXAG9
LmaAF3amzQfj5KxkAOIf0ennaW92cc027jBgxXhtz7nq0n4bgiXXL3sz1Ut9GKH3vScYs+ViuotK
6gSQ63R9BHgZCnrmL3rDJnonVFlBoXuD6bAos2t0spM5w7LUZOXODWT8C6dFl2Qei+g0Nyy7PcnR
lJZUO6n6P4bAeS9PZD4sm8sA2z9gy7b5Qe1cYPQCFy5/GZjMsGjRkgzz6FWEfmZqG7Crah0vq6Tu
EZZbwSf6J8FLOAiRoCtP1ojW7F7j9byn0bzeyNYo+AtosNW1FZIOkl174zV6TCd+QHUOrrUky39+
2/VkmSSYpV/X07Q5N8IaU5s/VCK2li1demt0UIe4+IuKslgM+kQJ+na3tMDXH5xP79+9YI25WGF7
pasFpGo6+dh46e2ShTmzxgDApdxmcl5WSC4rIMLcmafhIzNUy6YI0jnMzUPqFvb8Rdg3gMIVTzcH
ElCNkPRw+ETf7FEctUZQ8BJiPrNOuLXfuSxHjNI9GutDp3csvG+a7wWTxIp93X4lQPuE/pV8A8Nl
9ygUGzZKanDKy6/iZRE58ux1mG2tzh9UHiQIZrd3G9mIR2z9jCkVX0Q3JA9uoyyOtRhZrdcXmFEW
6ApNyo6GpeEE6kHpQFFb1wz+uS0pWxMjYR3Xsen5N0I+BQQquHG1Hv+dEsxfDeJRszZindiJieHi
KxxMqIcktibDzG4S7Wrr+EdCMkeNM0jzFxNhiEzqzj5s9d74IxuZRtzESKKJSkiY+p1jFBR3uYdo
iffUTcphZ7/usE85pH33PAldJ29FEojvFmr/7OX+tV9evcXqSzbIo3jsqOVJSU1mkH948m1BAS2j
FUwFc53NkAHmMJcpWCkCHCukvAOOwi/yC0P8hejDg3JmYzsKBpp3xiwSoH64I0LcHR6v36Xxojk9
4CylRc+1C+/siKZHkMSVEyFZyvDrwIQ1CZ5RYNkYi5dcwrAGA/En2dbzFHwDdM11za0uTPLrQzjR
HwluuuX7NJTVA06XzVBTA3+TlhtHTGvl0bcRmLdKaW3O9B4PX6yijoXO54jAQmfg9sXLdma/1K+0
vatM8UmQla8Jwop05YjhFyZUtpdTr0a+rCJwo8Mjnx7rk/c4QQiaVYF+O3a/rIzFNjlMJpAddLsU
hTM1o8uSMPCCDJV2KqfbehRO0cdl5IuMRunjqP1X3is8+xqdvohdFwYRHeAfMSojTbPN7vQHeK2b
GkA+bj//qjY+7ndiDWLPUA+NF77iMFp4ZPzXwZLXCoIRY6dQLUdZkzm9cK3GUESY9R1vyghPHdTH
IIs5MvNuTeG8P25X+0xHFugG9Dd1mQ/PK+p219JE6gsyCPj0fOE3QtcwdO6NerOYnxk4TMIHZdOq
q9D7jvUfrguC7Qxjny/NweOEZr8EMzQvOfs5Fy43aHYBq8Y1JPo13vYfeHEIy1wZOREdg3j3R9P/
5YDvR5K9dDPAoDv8UA2M7URloeVnIK4xhkBwmEZWSUE7tiFdvFT7vnARVodq9tpYCJ4Jtwyc/NIS
Mxk+RDs3ns9FYj+2tqEZCPWBSkqsKw7vAhbj1GkSaI8/x+XZY+/QBS6hAkLJS2WL5GcDRa99oSmj
cf3kId8w9nrebNS5cKAIvEhePgpfou3/kOdARdqcUVe5PC/r8iIuiOEGGcPUueumTH2jOfcuxCjz
jNXdO/WinXIeoLW9dsVbSEeqIXeD5J9FstqqZLoJVSzPTkj8RmAln8AvnMAo0wbQ+HjTC1vcj9Yt
2h8pkRmtxxvZk2VKUJxw4ygDqa8B9iHhoO5+Cl/vsZ4xd8snj8sIfzoMOzpBfJntlMZF+2uXUuKm
vllqyQDzgSdLJX3SA1CqVPWW5fLfy9xaKdQFEuFrtrrAcXq7zmuSYXJPl+NuH5u1RIGo3r/27xKD
CM/zgrRyv4+GZueHamokEBINt++/TC/8Up4H+smyR4Z7oZFgfY5MFMQ9KYvF5A/lZvhOTzEJvQAz
2bspgae4Q3gCjmY5MHD9U4W5ma2zlol3ATFIUOdOQDVnWnEo7oC7LrR9XxkH91Pz+c6nvXQzCa/d
naCqgRnol8haZkcb1Bf1cmviC/nDwA3mMrdxrWrjOUQ4R2gwQAZ7/6wmEZWDcZTLK4/Bwi+h5xMy
8acPo2FTGx5zI5I3QWcqF+z8+NU5Lbz5f8xnF+09oMH9pJy3qXCXqm8F2kaVaCNw/3sKWmq6KHzk
+sUBUVeSMCe8lyO7YQMxn4daSzSWYBJUe2ONnu1LATNvy3FzawsaTwWenUT/GvQ36MHLVRFIXaSa
lXzXP3RVZdrX+G0eJUqNASxj+5vEq6+lzg9p8TzQRK9ZgPdUyVD4TJOvdC0y9KRBV2TDZXG3Yvk5
ucTkZ0cNIUH5RB+7uWGmUCrtzPecAxwlSdzHKYlKjUtEF+DrgOCfCUidU/Puu4WbFyLkHyN09irJ
G4KXrgl22ZL/+0vd8qipqIRzcXcLTd2jLhWWPeYslKOtctN5qK5NXZGGi1B+OZGbnr2t3CHDW0Ze
m/6elnoYXQsNDpe5JqosGr8b7f/TnCw7kr90QB/UPCMwoqYwqiJ4q6oaI3LK96U4PHb0W4dN9Nza
Cw9daECCKreXPedDvXzCPIvJaeaKtid2upDkgh7Ne2v/4Tk/WLeRWycWa+AOf91QkOA3kZGjxMEw
m5Ux4P0bIaZczMnFX0QUlIBA3Qz4kpDpCrTMOQ2ZkbnESJNiQPOL9NL7BG1McsiDqVRNNTgqsES3
JzJmFYVIF8q+Vj0G8akrVmhbOLUlxtoU6g0SsiVJeuwQzmxM0hegpk+nKCsCj1ebWYY5OVY5Da6r
wMHX8cSc3yQbq2krFVBHXJAJyud7e1ei8jVEhzwszJD/HtxNcaWJqIHQ5QpM5/CnjBQMWDMX/JhP
82DNPhmExL7iTfvqGT+uOY26lY+rxn72/EFIoobn13L4gnOIMsWVW+cF4bz1ljmbTF5N17PPXZK2
m1AUdJrxf2XIv9LV1DcmlCTTA4yDao0KhTIvYg1CHb7kK4yrqcamVwQzV2Jh0C5ua4fFNIWZ9aB+
8MPHsGWyzWxyUwJLS+LLTnuL/tR+fwOTkUHb3t7FSACLZ/h4mvjXSHOYYWQ861YctQNfRCRLR+XS
yazPLLThr1RsH0A5Pz92C+JKvOQvgWom61QLrykwInzUEhc4w2tGAmtsoLW6/InZYZEMMNYVJFaV
4ODdeWbj2oul+arg2CmTLyiWmGdyxhKyYj6J1MspmdizVT42i2yWltcyyM5CtqtbwkIoiDc4SVOu
ITjTRyvah1NNdTOZEUgc1vZQAqMx5y7jz7lEqxH7HKTZYcKZ84NiONSrjZzqlbVUh5ALLVbBbnL3
5L+y1jP0JuXrz1fzhAtSFmqkK78XdSp3Kg25Hfo3ym5YDXKSsIxWuWqmTNDWm1U5cJ40/d3brBzZ
Xy64hz4BfJEevTUYkxD2ZS6+Cmpi7ZetVsInNFw/sPPCrE9r81LgHU3XwtczEsU8JPPYYODFV/Vv
Nh4yYFgxeQ5oFNWwzvR+1JIihRvL5o72vgfJUNikHRz0G1xOh5CxXJ1dMlwFucMevIfXeSfCBX5+
SzasQovB85MFhhcCbrgrDwoPE8KbJTHYtbEC5BYQG417bjYuZAKn1QD6HW9epFkT0HRANpbK7xMJ
1DYKLIo9F/JAAsYL2iZae53SmmQvfqKcwmE0S7aeUHGnbqZgsY9w0uRUtGOm2wjroifraqRBI1Vf
ALboTpNnmJ5hUZE2o4Y99ZakQKozTyT565jvBX0qu6TZ19Wdx/xO/N+ZWu77G3bAFgwmFxdpvLWo
vhros1XfaLW1xztoascXgZYJDGpOsqcbGJvRra9erR6rCQ49wU74A/sbqVW2JtP4UgiiSXS+/UDQ
zKv5ASY+SaIImaYAAJ8/5+O8NjI6/4dqV5T3LTut93nbk2mkK2ToHxWLk4qFUEisMzSsJ9BM65bJ
77JIY7Ceau02w+hqEI08KW1FdaF3lW5wnwnn4G+EM6aGT2KjrOiEPG/8Of7SnCK3FOyVb0L/MuFb
6Hx0T4EgYc4bNhcip1kA9m5UKpSovPxkh3Inw9Bs/VztJ6XAQAqt7sh4wNjdClvNMsifrxlHeCxD
EN0fRkNvHMNr+dAh2R4G84wJO2oWij/k4hjkt8u6dqKjkh802T1meJNoVNjqT5EfNW0QyCcxbubx
/VTUTwU5kMB18+WVwoSjwHG38DUqyq91OPzScYZdR4OSOYmDsjX2e8NplVMNum1MhFcts5ue7bib
gIiEraaqynKOBv4jACtjI/y3g7hDeocRIbyFMtmY/J6g/0ByROn8cN9RV535sMU9RxITIUtd3Eul
xi+LEvZ05G3P1FgMiaKwnF9Fg3I7lSEG8tQMNcq7cyXvqoEp2GQrvDOe23P/rNwhNXT8XI1Mu2a9
UndchRZBJ32vHJ8z3fT+ma0Iu5/Vvb0A9ZC34bvlM4NQ5uprJpiBoCb+F3CxVWyazZSUBmuMcp5f
kfltM/TlSyGcUXhojwJPA6+3vXzas8PiYpnaZxo86F/UgAw6rAN4tv9muBP6zhU/Zgg3mPC9sXbQ
vCdssZ98RJYM9/OwVJaREcgEpYqb4rwdPPNWT7AMwADQ2qf2/EDKJ7SqrKiwrVhzh5bx0Matc9Hh
6saCxubTdxIlaxRIWxkHQBwVid0K8/wAktWQFURncL/LcMKPSXAGW585+GJ5DxArd7lDRkt6yr51
U9BLk3y3IVJdCK1jO/OrS1/nciMaKtLN5JSfvCEef0ajSxKIQgCVpgPukXsh5PqfJhqM20y6QV0k
VpLGIebAYks31l0tpFA0Vq2sDhDvIwCjcyIXzoIcNv+QjTUspyVI5or2/1O22I/qn9tlj+HeH0Ml
DGbzn3Qm3YWRsK55W/kjQVwvv7s2S6rNVlGBwjhj9PssYS5oD1l8CSnoCZlHA6uqQMNZ6N4TUHhu
wazPX1HhCheFktiHiEjKUkB3fI43TV96Q4scnIg63vfFwtgaA48IUd2S0BoX95h2cGuOsIlQXr/Y
JCjKT6tBVCSYcEUxoDCzPd2nXxYTcgVPfVaFxdaX5Ndaaj73WCP7VBRse85ONZDPPYBvIdf3VWM3
gR7IcbUfSdOPEAqFk3UldvyezNH9JsM+pGXsha6vuKqcmdAbGYEaRlDbpXPn50IhNE2S+AcRP267
i8+CPYDrHHyepddupq1gzYIkGGrS/q1fz/D0fScWYZg8lXCYCBZ1D2wbNuKhitBJm+Fbsm1GD6eu
zAYReLlin9lWhA27TRgUCVj/K66+IZTnbYj4MeiClbVngnKVS9kHlL5A1O6fGQfbyXbjk4tjfApU
PCPeZXE22MD2rPmq6iq5YOlfLWz97NedIA6wtKf8xNGrcfasPSV2sBB7xJejnh2bifa23aLRV0hZ
SaP0hpXH4wpTnblb5j5ZxRZwgtIaA3VZeu0Y9IFsxt3HQuANF9H3pRUFyQYZkMyqSgcyl5GrTfhO
g8L8lCio0xDk+ePwipFzKovtELF9R8OKgaFgS9hM0ZdUf197XZg3AHy9XVnyLIfsUIZbQf9FbbuE
XOinON7OST19mhN/qgpvte09ZA2S13VfG4qwX8nY5AhhWXebuLsOZ4ynG8qSJMEzxnYdLdvYzioA
w+WYpQ0lX3ZPx6x3Vwk17oMfIzu5DbaT1ZdMWUhHvE2dzFvklNA8tSV1BKcIOfbn++SLubDUcgAV
UUj8yGCCSJKIa6/UtOXs2HES7Qm50ApN4NMk7bkAdFDufik1r9NQ5CK9AvYB1ZmkBR2zcwq+3v3a
pRMJUNnpKui3hfrSgYvXRuGPwn2FQ4LY3KmqBpirBxklzb2daaHMSGiphytPYBTJIl0yHB0KGPE6
ACriGcsBr7994hOczy77EfZWPOwuaPSPCAARaWtg5F28K3QV4Cf3iWZGiNnd9PU6JRmz3e0/UfRv
gUkJtXExeiBHp8Lxtpj1Q7DigZldeA/pNPcLFLELbWpYky/XLMN0cvYJLhJQ3X84V3/nDg/mIztU
w+Sjm/nUwG2Z/qysLAABh1LkBu1gOFRY+ESHqcrpRLaaj85eW93HC/ivkgh7y2ri0dNQFJBO5icK
8LCrL4ppLebmLIouZHYCNfjOcucSTcGnE8EyW3sk1vIX9OZEwRFfS7nA5orCdEV8HiKUlJTe4alC
wGhVX0qbXYJQbDG6XCaskyUzEkEcFmK+Z6RgEIsLXqQCuay1n76Hx91b1Tai967Hurb/gbqBFWS7
ssoPpotiuP7xrXMYmuccAAV8vmpZuXdOyVSvC8YuUMO32eRPTXN0nF0wVNcDxDRlkvB8LBTwVJt9
6q6cHCxtnDzkWl48x7KjGeGgLF5hvjNHSiihJ6scnAF4bjNCQGGj5DeLyD1T5En4XFZTwO1H1RCf
sVHU+u2tc6hK3drNPxCJbLfYCru8ZLVRZ1yC5uhkPwqMTAWtE11/AIRWDlMjcCegD0qxwtOVnOv0
RfXweP1zbEu5HYhthMF9LlklurVSXyD1T2G9y3MyG9fGX187u/Q7TeqY64LIePZuUbtp5mTK5FrQ
7j4kzse0N1V8kaIU03TvLVipssnEqHf8lz2Qz8kbZmISmr6Es4InN9NsL5nDW8F/mc02N10PIt01
X4xe22MRvGtsgXhd+OwxMKKJ1OTqnOBQt+tCIXIYj5JQojf0FDUDibehINFOBRnwxScJWcY2T+SZ
5iEw7lhzjTThhXUXxNXUtly+ZfcEmfJfTIvflxolRS6iu/E0fgZMP+4iTr/aS0bF4BRPUk22UnCo
xBVKWJc2nZ+t3jB4cwsNtY1jxUxKL6YZNknf/kSTl1hlRrGw3ceVEu7U04ueUaAnNgMdVralftDN
ZHkudO9GIdZXMKZFVN4EMzTGx/yALq+KzC6KacRcalWrXaSQSbU7dJm/bgSDuRtyTirPXrHpRycP
sI+Up+x+OJFAJYaTP+F5Hc8F19oPzYdutj0a5CXND12H94XbKksAn6LdMZ74NiPYjOJ5+y0SQU5u
8jHl+Qw/xOr4BPJCPjRqUhPBJ7p/VE448f0iey67y/fYJRi6jeZCNK/ZBxy7TmTnY/JCEPzb4ej8
HVqOuHKVZOuh3MFgY1bEIWgreDsZeIebQS8m6xDfu2BXZz5/lzaw6xHn8pFT/kT+Z+Kiq2qfBC49
vfv5vBzD6RxgcJqh5PIZpxsXiPmBoOf1EtvYi9Z6WlkRv/Tj+5t8+abzznzu8nHfWkDYrD4KzRDf
cMToaWcZqppkkIY++LFRRneMomHU8hfuBL1MBR1LZfksBRgEhhJMZ72PAaWoLePB16OnDYgubqnx
d3vYcMB+gWTh9p6z7J6XI+BxYeAZJI4mvr2y8iGxsLHGGruf84TQ4mcIUxT/LuqHRTxY9BIGVvMN
1QXAL1c1HkMBKY1xHYFvZR70BYJGyTbwxoSMgHEr4G8vzoKwcPQloADElyK/kQ/mYlyBqZHk4Bf0
Wr+b7VKbMntK2BAZDGbn+APsP+ZF2wJHayBrjfmaLgP+LG3gNE1p/xLRY/A0rrefcuXCt2lbNoTQ
RuZ5+n35sYiXb2/IGRcipgo6wnFh835SxYXny+jvIpb3doMKWgnCRR9Gy1tPtBHDaBNhX9xntC74
JUw/ni1PNlHzuvoLFYq2RgXpDqpOkNCXVKspOXNoVy9DUIr62h6EXeTsfNrA+zapJ253eh3B3pZQ
fZ7s6f+i7EWCCadFE+V1sbRv0fBA+C6UgVkpo1jFPU73Q6fUNf7kYT4CebpmjqAL5J4NoFJjYEvW
qdbhrq+eK+Hybyiik+G7kamN4cSdNrTxs7hxlsTb04SndYOui9HnvCnseplirz4FYRIO4gZFgo9X
VbsRg/gAuSnlZD4kKSIY1t6UkhG1BGMcakbnYKCL0MVLLDK0zZzMfz5PGQ49v3m0xYG9z1UU02CK
aIyo7Rps0U96UxWEwOi1hIvAnpXADXBZBiFBlB4ZbLWlUw5MFCYOmZbpt8Vosp8rrlrdrcUsnqOp
gah99EVd7IDTtMv9OJZu5tmNi+TzTsoiJJ7Fs35AcVA34Fhja4vyMZEqbH0f+30sdwVBVWEo55mQ
jWLp6iaLz0UhUU47B3fdk1d3jqTk/mj5EFy+22E3ZfgTxmsb/y9HQcop4FyvRgVFLS4qxHnjmH9R
tl7JBtQ8a30ECKbIlQqGCRIynxShUkHraRg+XwfRVg3dSokU62XkmyavbUf+48XgdkFqMFXjUaPr
lOqLOWuhkR/kK5DlFFdhbbjLVZ9JvF5sciGsMmafeuzOT2pXcS1ribInXMpS39gT+zpONpgPjwc3
uT5l0tJYnlGjc/w1yoeLh3BXO8ZGg/ke60vEUiykoWOSDeeNmZUC93y5FZ61TvyYSetOh4Dlnj19
cNNNSCn9o69FZGug5IujUnMOljzJXV9gN3hTkG/tC/yPD7YRuCJyfxVfUZ6vj5lzmcegs3a3Gw7L
xYfU48BkLSJVl7cYf497aGghD9RuQ4Vz/zMe+K/qt0wifi+SpSGJa2Zpr1+M8pT+Iggl4j782b9G
AcLubpQS737bEvIYkfJ3LpgCwTbtRxa2jzjn1VMWD8icnHZNpLxixFJDitgh/gXbwdjl32noyBOq
+GK5fqmVncYOdkQ3Z18k8RNgl9cHGmoG8tYKArzGlVLbSYqDb65tpoSvCJo4oZsrXizYSEPQXgev
7NG/F33TFjK1FkB43p5JbbKlGhvSpr9ZZEqrMlGeqM4G4+oV1fcZpXLXVypHCIr9EZWbSMHYDxoX
shPDnPC990lObm52AhgousGQgsmalbs/nU0CB3ok7etvidj2GCgWwDG2kCNmj8IAJSANF9hZ+BDP
K7d5leag9nQS9K5D1bkPqumV5om4OzZF9ll7gCpqsvVsI48m/BmbWauAp4076XuT4t3E+BBps31p
bSLujf7lbU4xA+hpEZN5GKIkEg1oyL1YjFWmikySgZUF0AKs7Wj/VXd94g5rBBCMjIxnoHZQeh+Y
sSOwn3qgcCVv/pPOGVYpLrKaiNenaRFI+ifKoIf7cXqC7LC4NC44hIn14naKVAPgpYzOFABVYvUt
/4UAVIWAynxLB4/+dh/mCDjeJsr6TyEyJk/9iyexjP/qochHVHz2KDsOihp3sIQ5MiRbM0Yzv8lZ
ko1VoSkhZm3v1e6rOyGQCKzR3fGpMuWBznwPqLfxI3L5KEFr/MQFZom/5EWxS2vKsVs1eJ+00BmE
t/Z86OrxavVact2LQzCc4e3NS0T3022L/lUlsdi420BU31wx19/GsKx5U118Z2uoCfnEBORPD/Bq
GqvgKqWmmFmqcV4KjrmEIvvs+nFFOMK6r79BU/xKVdSKi879uKZTNzchJvTajnIr3Po6khluniAq
E1ImEiPqCLgt7H+d+yKaT6ycnKABmMOuc/UkbyV7wWihdSpTKZwxLnPY7Kz8MQ5qOliXQIhttAfE
wISqf8G/swuZoNcBSdQICqJD03Te5v/E0Cvh33CD5tXRBy+81miKpe0J6cPOUnOFO7Enwn34NvkR
3udzkRb0b/y84YbkdDwI7uRvFjQxbL78zAtF0TsFk3j92aH27fX5dZ598oXLZbdhec53BojSw6vQ
O4Zq6nODKRtrBhojQPu56MN/G8xk81dWX6EjZNkW3QiwfzkAwJa9By3Ha3CAgIIhxihcRtPEs9VB
8aZNgpClDVsbDszF2I6tOCSQA5C5ZnhhG2nuffVVJfIq0I7/NECeVa6s3veUNfguMqDPJnPpHCf5
S5+wlQDnX0eXSgVFmEAp5NH2tFEGFbsFADPq0aqw1I1YfXVlFP298XHYUSurFbxNTlBa+PeH2QD/
yWrdpEIVlBy8Y98l5Nr1qlKgp2E1XMA5kIlaOLyxKl1qJ0NuEFw9+MBzgKn9PHfhVgHbRQbCItQJ
GppIaKIca6MS4qaGVRaodHH7aP68h8C+WAZJLu3qdFhoX895h5PoWrPmrN5TwAsDpvEiuMIy2K4Z
kyNQ/unacQP7uES9WzQ5KdyfVBYAGWfbkpZLAlTFGvJW088aGvk09ZM/K30zmMM10deWvIFe4TeY
D/GDkKOT3Zcxx3kSMUkHSJCCyoJkBUYuRklGkdjMjfCFOAMZZpe9VDW3ziJJhvbIbPM204kue3y8
6t7k7ey5iJxqvhCsRM/6QaAWuq9HNZ9PReQ5b0PCoolaxGM7laa+iSLrou2CrabOKjFbofxaxLul
NMhA5eP+ydAL4xEff1cGKWKWOq0aPEahD0yu9BuAp6Ax0zlUVrERDwNrkKiwG3Mbl4AXPtXnclr2
IGlwc8KqzZ5p69QXIy/IxT7C/hKxrfm/r12ntSc6o74LEOfSwgm+FTfPTx1T4lOKKywqnKB0GyXV
M5ujZNuSKBXXmkkszS1gMx7NpccOQ8+Y+r4Q7NMnldmFD5rwsjlnMN9QTNjH/Hcb83VRwtg+MXsj
I6QFL+QISXrYarKAtk/288Anft1jH6eZVFMMUcOxWoH94zAR1Isxatr7bxDzCLrHMj4DgqReyeMf
Qsi8lrjrEALjWK1+y32nXc2m77GZkIagb1TPORu40F/w3euHXcA3VIN+jiSUq0XL76eW/2AY4bAI
fV02p4kEWH6Kk+xWJwIElU8ndmcoX48+GPNXKIefKeM9xrOu9c/i9aEnN0mfoi5u5MFuTDLD/TIp
+XRCDE11TvlKmZgIlj7i5CykNANZZVVgilnK25PvcSm/J81RfJvzDxb5JwZutQMr16qcweZFFALO
YT9oX297LYbg0/1xeAegsec4jM/bj1PReCw3NI074sS39cj6OlEpoYkh18suxb44CATbWHnOwZBA
x/ZXSFIftHvJoFrHoCO4M6MN4BKCCaWce65KvnfX+gZ3qRb8bfjwUpCcQLMtmS74wep3q1647IQB
p2JnZ3UFkw4EeQdg8Bo1CKU69zQhYvchcVWObawYhLGREXkL5WndGLqUCNLPJnonH1pDI4kk7BSI
Ey7uqvU62EcArmnGpK+eTAR8SwprkDCJPrX+/Zm5bWjGtxW8pFG6rG1Z97klOsKTTVxup8y2ptGg
oYjXOIEg21uVu4CW50fdUyQ+TIWolaj1CR96+9eGqHKRyfq8Pa3kRjdCP+gnBkX48PGCxtWi+PPz
+YR1SYPd75wwTaneMeSlShGLNRcsT8ubbHZrPt0QG6q5B1UPkGiVAn8v+LnQ3kHIDnv1Nqkjag1s
cERfsruqCSHX3oHbq01ypw7jQPqM38+Ohq+Uy0fmXoBl7rhNy+sTFuyHzaT55vLLRNg1Ra9x52Yl
nqpNmVQv/xFCt4MnUotMxqymm8E/Mu7ur7oQPzgwOR97N9p4ZMVf0/Zljh1PqhxXiPcFn2BQMUAi
QnYeBIrjmj326GH8M84NAI999u5PlyOIzJQBxR8FwPOuqUs1dz6sP7G232GNX7luGB8NsHKD5BA3
tgHlSzFPWfucdHI+M6r5Pbx0U80yx7arnrzqgovGAIHy6LJVIdKJKNcn9fH/D/iBB39tm3dJ6WDA
ubKwB8ehVigog0tfFEPxAlEgVW9RygPw61kxMc6Oehb4SzVNSPinynYl9enU/1b9k0mNZq3pKgGI
ByC2FfhkIZ0PbHlMrz/i89OLG4aR8Mhq46b8vZ0qpknBtFLBUuEkCa1LGYROsm4OZ3GxgTQPtCDC
QoiQZfCfBrXMJH2irnDrLlCbeeoQS9UP8rONFuHmHwUfWQZWu2amaMVob5SDjrjQk+B+aUJDroDu
BNX5vheGo2P0dxVMipuq1/zDTnoSSayFEjh2bz+WgJOOqZnuTIG+QdJ0I75fMvAmg0YOyHRmvoyi
XVSJeNMpblBWqBlBgzu6pGoozTy/I5FkHUFw+XHY3Z/M255dswEzComyu/BCKgbsvoD6kauxanZm
lRBGrrwqJvl9cTBryEoPkqdhlDittw6ntGbAii60OCMHZWrLSV+QVnzLbwepGRAs0+xUkHy7JA9R
LazchQ55VVcFJhy+QZw3qGOe2QdZCklgcq66+IqQuBkksl6jLHrc6QZMa/XTuvpejpS7QNI57vob
Ew0ztdZb4s9bSKM7G0wv//5UUuzRw6wvJjaN3zykh3P6gLAbh8FQDeQYqChdEpljQPMmBfDET2P3
GA1zmQavBGjR3/fb9gL0vhPYItPvYuwQjzZxfbrXdq6lj19hIj8d25IXcM3VeFWolF5Xy9gSGhey
KjzBNiH/7RsXb4UNK5B9PwTJMR5ulxK3YSob6/I8pv9DY3f7BQAEeVulXShaBb7Dqk1sz4x4rGz6
tLEq+laiUYlvX3UqsK0OU9BPICs3x2PGKlcz7yCWkwg152HG9EejuEWKnAH+aaNLkk6pwetQEGNi
GWqGR2AosJaTQdrhBzOcqHzjijKOGPz/69PYCt0N8LIKLlMg13TGOV0KHxnPus1TgqQ6i9qnkJKI
vGQ/W4YiX5ndZHrtXtBeuQFgH1IsK+K3sd8FnpkTBqK8NecKyywOYVIlLUg+3/YA1k0FnYmsOGDx
jAZGWVKQSrlJI0YzmD+J3mzXPoYbjE+43cyeZ9WNb4MBTjbnKne10E/LGLuDkGtcdp+szItIVy1J
Iu522HQjZ6N1ztzyBCONo+0ec6niCXGPTGMnRGMikk4ca1WK/8B5MebWujJ8me9HJ4G8H73urmCJ
NJJ/iG1TcY7r/Q5zGmsHW5j2SHxfci42XDQ4jSXghKzK1V0YlGfokXuv4TkJcuJf/IRvP/u8l7g9
PT/89AuE9LupLuDp5T6McRS78bqI+w0VH4jywABCtnvi/BQk2+KEfU5tyDElzy80DN1DX7XwEkDl
H89p65QNT9mg8CmCzi04fhqRaxn7M1mk0bEnXuaZ48a4K1O9T7RmjQQ8Iilsg5Z3VWai/x1UDG5s
u9/VmdubFt4n3PiN0hY2DAcHpx1mW+3PWkZdqGRgT8PcsK0uRS4U9+NHtDpJEIXlcq/NEeUjIq0k
5hK6Mur9sw4yLzTeKXBoM7CpVZnxYbUNwx3vcXysh6HCE4y0bWO+j5Dy0cQQBncGoODos0AWkKuc
LYwwOkt8uKiIMQGyJB145eVcamrH72gHBkDYJIVcVGlYc9EHQ/L1rTDMea+rdsd2APAFSpGsuPpt
ypwIN2uUnmwA+mcGP31ZtvgrBmf/FwLSuQpxpI9L3SUE7BT0wybf5A5gcQRAgk/mIHOvO5oB4rWT
ZsysA/0XQvYoFl3svz2eS/gBGzzZx60GGIqnuPxzqtKLk3NkZKoe/nKTnMgZsqH/kMzORVBwTe6c
mAK6gav+TdRYR4Tc5/Agc80mmcKTx/an4W7oA+AGImP6LAbTsQ0DHgBMPDPoChvpD5TKAB4Iafdb
7oL4Oim+Rh8ttTEPyRjrwuaoj9HM6frF3VunnAX3mBjrOqYjeHZ8K6FISf/VeqZMljY0/e212VKp
X4m8N9nru9WhX+LMx+xwaddrHmxWEGO2uR3cZ9+Bx8KPcQyLTaQoELqfirm1jjiE6C3Zp4p0Mxwz
Ir3dakozfyHr4O9sNFuJz50U68c9gXctF12tIHxovaZrnHf+/BkllsKZBO98sdOIx4ZBYXvvuUXB
A9VZN2uloNXZ3RmBdMmbht8tQdN7shrOY8WcWmaBGAy8fxoWVLeyzCGw7jFJai+o7pUxuHhPdRrh
plRQP1UM4tSpOEALevPWAzqmki0eQP6HvgEMmKDLPMA7ffsGuuaMSkNdA4Sifb6eU1qrZ1xHHXTg
G8rOzXoNz0Rddkv0CjqZdXlPPU85JcZFBIoAttwZFDN6iFpsMq5wGRNL00PrZNpRyaRKI7C9omUO
xW+fuwYZW2u7KvSNu/BfBy7t8/xdgtq4T9BT7unZ3IZct6yDlt+fT2Nc1aWzzIWjpVuBIGfylxdX
5pR8uzVp1uLuouUf6n6pd+oosCdkIUcN0jr5lSVil3AJ5LGZ4UVC2fGXYN+LvWbq6sTU2FpCkgpt
1cV+HvWz3BfG27vVONf4wfQ3fB263lOyJyxQeQD5uCUObsCOkmuNZ4SjFoXt7+ST2MhFYzwy2+ku
aYQxnUAfqHW5zdGD+oZ4l9ZDUkRPaaeiLA4fU1LqNIY/C4g2UUiCjyQC2wvsZJH8KnbiFI6BvAdj
MTfnHjDFMKdvvI6oDCkLZHwnrWMk/riEMhAMnG5jLv3tjMguhZb3YXxBgpUZbDJajamIZqdEn1vF
X20cd5ZVm6kxYw3kazlt1k4ZyQgGiWg0pDeLU/ZgmauphuB7zP1gbm0VgeJwQlA34Y+KFZCpwO1C
7YhCefMr6FT89AeDdboqcLE5iLc6GuwN1C6PcWmNXbJuLi0qWFMB441NK51+BYWvJpNFbhgyaePi
CMu7f/injfofaTMvvNvNb8Z97EnPHT5m6GsTJw5kg/Fbwmcnryc+TSmlfkiG7Pvrdp7QCKTKTXY0
ABzQ5fmKlugg6K/gU3qi2yUG8dsRyftrH6/Kdayw+QzfCcJiNOvIj6woOSWXfT1KT3U2RDAkJc+Q
XqNu5IxZ4w8qMmXCnYLEShQfq3n8qeUbOU5enNnj5hE22N8lpz5jfvSpmkn0HIu7C1vNFhVaK1ma
d+bZOundbezscPJIrsS+GZsxIVAhS26vGKOzFiWDLQStpZPu/AJT6836jGnDxGiABjiLsVhxOQYH
Bzc+oncoW6dORE9doWno4b35jU1PrpXOv9id1YDcFK8IQ2yI1tAKYQMm9F7bWqjNhJ4CwbAmyXQR
6Oohr8QyXJuvhZhgibek/m/gy6yiJACobPEAbUbuq7Cnk46EUDMwYqoF/pgiFcrgloUqHP/g71xh
bHP7yp4p86pqdN2atgTFvcKEUA9STo30oNEn9GQkP8o4i6nWlnMwlVkPgm7GtoLyxZIeMJwyA5U4
6GjVkx1ZnQqEBK9q/DGQpm5rpfnC+u0Q+GaBNOtP3XCSiWcDzeqNXKpNtYO0rIw8O1fMWmkPedf0
fLhz+U/o4sTXDJC/1SD/ULbh9/MizfMWrwWSblUZVQ8uKGB5BJQ3HzSzY8zlZl4SHoEBfgLnI9N0
l/Yo5JgTVmnlqPcCpGVR+5aNUCZY9M1Hp60q83xnBrfY76Wu7ObGMtFa3SmIWyjpsD/9d3Im4dnb
6SHkpxM6HLjTnpcy0Uwr653rDWWxoLvWJbt9TywcRWiXCP8Z3zcOI+eK/kAoDXKrdH5t8IOK+ELm
G59lQ1FsUU03Tbhipq8WBCppxNjuSwsGon9VgVnkTQY6EbmmYqdMoCfyuWbY/ynbkE5UlpgXoUcT
WV7zG4COzhMfyjhe1FDUFVQ3WUJsUjHgj7XZpqwrRzcobJ9D/wFF8LeJ8oKaBSVbN+509Nx0NuEi
yKKH+RzvCpl0ACu0Nup4EVj5bxEtCQ2dRe767B4PiNMTZIAAFjYQro9WSy6+iSRQdj6CwBgCY44Z
jC7sMGgRDcax1scMhVsV5bFQ8DvZXtdqz1uJFhxWPIobOIaHWgQq9cB5wU2iqzNivXKPVglWEBpx
f+o/vgnw7Xlk+GKZakZdcjIzvE4oAGsaj7Y7AHNv92cLSYdgN/FZTzSq7Jxood9874kjgUhDMckE
/jz8TmpkP+S6gTC1Y6rTz+KtQiqtbUjuPchYyAC/Jnq1ylhriB4i4YIQPGfWQRl3KH/FJXGtSYqO
CpLddd/IfwpfN0J39TFvKZfilLv5jYDlg/oYdmRnT6YG9nbcDRp+uk3kpCp3Clph0elPUOPaegdF
1x3sK9nnUYhHL5tWnYUUNp8kTinGZQzK0l73Qmo7S37vR9qIQ0aGkSNqlaP2bRK1MKEBfSoN4ykx
gsV7eXXwrvp1qT13g8NJLzSN6aYvW/FS/jpfw99N5trIrbM/w5ozO/CcNbcnJHbjq73Fi8CIZHFm
ED6uyPzQscbfczqSbKyPV87EnMNt6cejMoa78T+ainO2ExLuX2reU/+vtPjvR9/uzbqq1EUkiLW/
nBkCLcc0LwuVg+rt9Xw4FiPfuGfYJJR8DdP7Azt6bUfkwVrUgT/ox25y7NYZ3E9Aq+pE/RA9D5Gz
WLoNnZmyAGr1B8zDYNMlOQUTdr/iFTyVV/w4nYjcY8SeXFvX16fIDUPFajRTDcP6T9/a3iaZXGC0
af4xCbZz9sYr7t4X9ApYOoEL3v5kL+3i2vAGG7bXMJH3/1+psm6F1alfeB+v1K45bGxI2aUXFgQr
JIFlGtYRcGVW385yS+KfvwcgxOXerjk3j2YqcieBDx++Gh504PmW7uIbrNIcJAmhMxBc2EFpFaLW
6uN9uD6mOR+w/KwR5Gbi/gnhV5fgwoPdlpRKCcp7/9CITufmfjRD9/aHFmzh/A3nW6iZXdtvaDxP
gskj5v/6KvV3lMF7JMCa4pbPy8jMt7NPNGzw/fCZFVKvMZDG/dfhQawIi0IBD3VASV3nLhHwBp2r
6FCync8og8G3xNaSMCLpAyNFPN+lQMEZIxpIlDcp3YJBBgPEToAvR0Y+M/cwFNyiIygChuYU7JAF
pUzeRUmqMXATKSapIfbNOxY/F67HvcyUg880u7vwuTp0SsqMa5Kli6KDqQdTtB/8FTyNJcGqnh0a
XhcdYeVTb0aWWBIaahOL0wiukPSdNxJosRSOpRI60eSwU8PfFXuI/ntar0w+Ei10unQoCH9RjKfx
G1zhE/W9PgRAWlhw0lzrIXNYxjRQ/KZtgtMtjBtj+F+O+wXf6KLOmGXFPaSqowb60tcmtYOTnteI
1bz37uE42T4EAenx2BNZkRdxVragpO4/rAuS0E3qRz2E+bcvaZj+fGO31lVQJyNIKILb5gHF7FY3
yfUj+jYJ8d8XRu276pI9oDUiDksUNcfK88Cu2DOe9nelWjYOeIWcUWNL9tk8Y0xlIZWPqLJ9ypCo
3z4ku2Zu2xViySRH8yovulIUCymKHBz874ykONL+/dvyKEjDNBLYnjEvmyOGaiUCE8BIIKejnL5G
XuhNMiTPZJeN1eI2V23vfBXbK/4q/ytyQ9DhHr8zcaXNoFwAzV7c1jqowUl1oBbI0hPXZcBqNzED
2ne21NSvkMtQK7V3aWo/Ggt8hY8xI0BmURPtc6zSpxZz4k87Azuevm5vqCXrYGjOb41HITYyAcgF
0bzDNrBDpWKXv9jNe6AmEi0mk5g+G/srD8XA4aMuw4OXKmFmesSxHv6eWdbukAspMIk7NiSm3xFE
nmExXg852sGp0sKA7Z5U0julIhcrrzngmlK6BwtGBUOtrGWKNjeNQab1hggHPffKfCL9wrcsdj9v
Gdqu8VQkMlx24ydVS8R0+B5U+RIrw8ZttjZuln2kXm4xJ6FrCGj6SIQzdPiihEiLlod8nzi+z5RF
hibX1i18KS4ejok64pMx3NFk/DzsiQcjhCg4PaRd94b0gOdnZr5WCfeUetjQ5OHiFfTlqHLpjykQ
UKAL0q2D0FTGp2aFNImBt3AMxc8of5l1t0LdPLEgmBoByC/vuwvQ2kPDmQa4HBx4MLydnnVnGrE6
oQi93RvpYU5oiz7LK1AjltHbGUz/bCbZAZr3RyFLn07D+qV/S7t2wuKbiCs7aPjLgIZqV+0pdWd6
h5MElpyOwBPZkV5YWbRdxo8gJlq/SWOFHxbpI8eD+fptkWI54yO8YBCvUKOBFXUbzIpWxRBKkcSe
ZznryG4hej79eDgtxex6Nk8Oes5ZxMUhy9VX+yN8IRfkC3gaCZqNbrnCLlENX5zsOdr/ck94uzov
/6vjhZNvTq715u/xFHUm1pfYqpTfrJxTwt7k/Q4zcOTboreNZDe/YVC0jhNQhU7Q/mhIHNWx+0Sp
fYcmUN1vWBZmv2R1r1cR3bxGupO7veJ17gnHq+sdRGR8FlLeyM67+EDKLZkf748ZnHisP5KFjWQA
s7kai9giFT367Xe+l4uWKHNPriWZspPpzqGA+tBXKszSIbOlOWPhhbWo5PwGvt7WNfOQJkajEh/L
y8bJ/RCBoZSVi6LLAYpY5g5TxDr73Sf2nHV/Fk/0MMEA6EKnERQz9nvGdJSBgg0n8n+sgvsojXnq
+LcH8CrJwRZqsGejalBUHkcL2lx3AC4dd5LndJttRnKJfRfFhE7bv59jjCBWDhmDeuQlaTRzfEQG
wY0AnC+UuMc/qCj5XnfoLO1L6do6sPVlkzAePEzKzg5VOnOfUM7KV/Lz0OZ0LXbGoM2sv9cAz63R
No/PYGEt1Fvfm24NiKxaafEY535UOPyHk+44g8gyax/7RMcWQFVT2rF82H5D2Z1tZC0RCepgn6GF
Ee4RGarmIkYJyfhQsFM43p45KHDfYb2BRsSrMqVyEZtTps3VidEWzXreGSXpngVCD0tnUztiVAfp
HFct7tdmZq50/P36Gz5MEutwBRM156Zi7lyB9YWsxanWlyQH0cRK68EEY+NTuaKLiU97pywnNVAv
8p7F2nW7N3YGqeuNEd4EWpn+iGYy/STBICFAlrmr0UqAHb95/jV1zcOZ8nY7j4p9F3EtjQJaBEQA
mOOjafBCOHEKXSXHoYrThpaVw1WaR1nwNA00T/NrigwfBt/2WZj4OQ1fzTVkLJ5vkZeaDZP7UAOD
ECu90ab4PYifo4LeE03JopPfih49EPJGH0xgwfTdtaKwDE+Xq7Dy9W7FCi84NK2cO9dE/3d4LxjA
8293zxpyzK++E9f3X9ilotK9+n1Vk4S4CplllHSeRpXpSLAZJMiloxB6l0DCFDdYWQpapH9UaKuz
bo6/xc1OuZXVBGIlEVajEGjicJfNg0noOgbipUY04hU8z4tQWETQSONuJVXocC1eTyp1UvdPHY8u
1AUc2mtpLQnv8Gq5Cn2W8g+yb+5b73SRI4I9b/3sEpLS1iWFd4NZqCHGCZLOaB0jMgct/18x9nMn
kh6vcMzV30pVf5MM6vebLr1R2ZZZlj1gphMFOI230I3wWlSfXq8Wxstq6vLN9vpEAgc22sTP7QZZ
MW7GNDjTlXeiavYhRmai8h6OqCjidPHWL1h38vEpfFrsKqlwtrPgaHArweJ3vaVVgQNAjNWaYd2A
kVZ5f7ARfritWW/zwXaf/dukAAyNaTpEf5L5Rvu2zoLIMocek+Ppo/xHjjiK2xc2K1rh7eslYAId
KKCUGCK7E63gLrNRwqKXhOk4e2yhIIF2y5GZVVUO2Gkya7Ljx6/7NSEJWzztCtKfSBzD9blr/Z9m
mZ/vSE5AISyScvdkClM0MNEhzv4Hudv8/WsJu+adglt8yGoK9Bj0Ic36pzXGW40qNRLqr0ahAl6Y
MIFFGTqXDG5ycvqWqZF3OZl2FfRGvn1ZYppmKqNXIXYO3zJCL1Q4UDG5doqeRYZqTd60kAyj8Ir6
Oyhb45Xr57xDq1Jkc0XnOds8Q37tDlQHqWz3w3DXwiGIuAFzQF4+xWDPiEWWSKHJvS5i9N0gWlZo
2qupGlucPIaEHaELiajWqaacYILD4b8YoGXoNKRckN7mu5dHfXOWFY8K0+wY2qgWSDo5LxihqFG0
r8NLpy0HYsc9f56DswqfL/cFuibUE4ez0+ZGCJ2M+W3QvmyXStT1J2wmmA6IJ/S57uzj3N8/pnH0
zQrSW9xmsfwQL/q4SUbqUubJqpaD5ZdZFtObMffhByzELz7kXd0X+gk2El6TFAg1B/9gOGh9HVdT
UlXyZiH9mRejXW9DZHcyLWATSCDfKBJR2lDqQeS98S88vWp3EHXav2lxk9MEQgbmXy2BFVs84U0Q
FhuwpBJ//mmrgSxH5dLE5dzIp7nWYfzwZOtvGvbmhx0BFLPV1kf0anVQd/JHtb+8p23nK4PBydtb
yTZNwTGfHXTdRnDGa5DVCdDJEv/9aH02KYc0iz72tf7CqqfmaLq9XdP862vsFz4FYUkM51KL3FZo
Dc/E2df7eslNci9Lg6hGihyx6gbrfBX6bEXS19q6lpeuRr0fr4E9RHj/j37aIBW67ET1qmQ5WsJQ
ArYAXVC9mEOJ2Mg2jaCic8XqAcBV+2ZfLI6jnTs3xy7xeVS77w3S9UEwIKfkx7HKEe1B+79rJ58r
Ze/LtTig8uQ2wGEWeeSPbBp4qlg5nI0k2xiOHXrBaT859g9/pgdG0o9VtuYyUPzs/Ct4HR1Du/Pd
zz8C3L9ws67GUAhpkbdtQEWKWI/LqoQT0d/KKlWoRttcU5quOexGee4VvvEOwcF8owcsQeNUOsuT
BBPrH3tNsGUHFEmPABtviosvj4Coxu6cJX4LNzqzKOYUoJB3kyp0zM/7InyqTMJH02Ialan6b+RN
BfBkpGrS2FI1nchEpTrPYubmL4dfbVAq8FcZRl1cZrM/BaQRvy4VegKTuVc2lZJqYoTP2PppX9oo
kSa0+FiDcWqBPiB831m5ft+jcBAWz6HEKzAeHFUT3rNa5k7a3SQ95ygGK/t12bvCXJ0X4RGXa4c5
hCJyWvx3qShDQZDWba1VtPhQmiri5dzOBGs2i9IRb/vo8yvko4sDP7Wee9i/yQIDxmZoOnzgO2al
eJrUdvGPwYgKGHFslKzDIq8fqOvcI081kHVywkHkegKROBDmhgMkzG+UFuqhpL9YNG6sIZAw/rLA
ZxhzTrh819TJfZ6hyKDw0TNZbyCMk7vW2ywTkPFuMaaByShuk/C9T7fSTeoHVtzv9i6ACxxdvepg
ZiJEJaouESVNk3AC5cTgg4C55P/mPLWPNuYdJi+82RzdH4n5SEac3UxdrJw+5H4RnfMw7mwQfU+r
dBI4c9klwq9sf4U6rvxFkrzvekMFhu3zj9JEwZTFMUswgGy/OKIBx9tiliaLfblDU32RH7ptTSso
Y9yzhG+R9ieloXTZVz6IoZD9Puj5BasZgFDfF3AODtvDWlqUJxcretzxh3RbGBqsVIUatd7NG2GX
fqA/Zzpv+PyUvXDQ+wcHeGsg0iXcqfnr7hoop8eRZq7yJBr8Z4bCY1uMfjE2Q7bnBCTztZecWQt7
uYsPO0WEfTGS1f39rTpNKMr6J52mU9dDFyZGKnaYCF8CjVGMjJ1uUQ1A+mA+LI7BhGeweYQD+Cia
bTAxkohMiXNhQ0f8xGjTNUCHlFlTXZv1tFR6M8mAuJ2dD91Q7rma684Z65Gq8hOmXIYQcCjBwQ5n
auxlOqYGJ3cUNSZGiPvxgAUPwT1btGLwkSvmn4v5uJduL5HX/ZrrNpcMhihDg7Zh7XZfI/YXgNfh
dtMrWK4DYUv6rdqgLMOlUk3o4GXHGeqmcTkoZ6uVEKL2XLC3c63UCWfXkXqv//NpOCY/1aPX6B3x
gqwuPVF3QGmI9uaP9y1blo/H+DOZMyjPnvlY6QUNGvUV4xq1Ntt2O6ZzeQx54xvmVG8mKDgaaRlg
4tSNftU8+WRTjFUkOsXxf/osYKbFkG43L0tnHsZXVDGtqLGUie+fhB4T1TpAvaRE5IrZK3egmn3c
96clECLYCt6iFvBHMspIqcHbZCDlLEIiz7UifWEgXIT1VJtmDq+4pbFsH1qx2eREhQ/5V1L8Mh84
8e/tQg/ytHeggl2Vv2UlBKTfzQ5uuTUE5/a/UPLbxOrv5BjDRHO52t9MT9RrxAgAg3OJdJ6S1ShB
vsdAAxgR9lZyMpe1C4nP4o4Px2OOmeskmEuBK1erTxJh88OTH/Y2iBVxH80+tHXdfRp0T5zdwcoK
TefgcXePRZxSS89SMUHnWNVO226NAvIZ/ZwB9nKpZ7zwnlawP/Wvt+cbhLph0x36DbwEP4lZ0W0P
o7ZpYvznN0gDO7GmTGUW1/SAMMUqB5A8pyePYp/oqnHXdxAm06KeDCWDyMKEP9FpmkOMTFfSK0Fq
XcFXMIuSFK1P6qE9eJm7M6j/66KX7JrXBSHmlTp6zhw8SXwKUYs3mQaFQtTT3ht+ytdFzXWpnWmC
PUSAyAglYcAfK+TqhQFM1aQDylqelLFODSLmKjEtivPo3/VxeesA2uAAakRENRs4U1ZoSukdCv1l
Oenz8ah9gwwiVGFQRn4hcocR/V0BE3PrpEfThlOJ2SM5Kl4i2/CwGJXIHUTMrINJL1uQGm/TuP8/
ubjOQSfvv2SHJYbwyzZjDFTtudwdCebHcI4nX4f38iDMbiXtYZ2aw5fD1LZ1aSVK5kWEYYalxwqh
CqVuxGvfi/IQCB4U0UrDhphhq8PSLWhHISrz78JPufgF410ThTqSZdnivwDCusajz6wKrkz/O5ZP
JiwF/9jXT4nYA3RIpmcSN7vNLAyotDhyObkaYAuoXOJ1EdJU3PbSwYGVqr3qPCqq546Pw4lRV7q6
WIxYETfnOC1ZV1hI0d6dBZj0Q/OPKDQAg4LBX18v4UrZh+b4zc0tTCBMGUwALxcyMl+WwJQuejnZ
vIM4nW5UAWtHeBNp9kBdv9XU6sBOepjhZTVo2mYA9RlD6wnMmeOCcLYak5IuSjSIQSp/haHNQuki
pPUAKJx7BdiIyl45J0jI/g/Dn5/J7//zsP2dfauVrBkXXxPt2Ppy7HPelJVSHwDXxXk26wE6ehTT
1FQ9QDXawp16y0TRb3HqOQ+XphznzDw+TBP/tvro52NZB9kB38N/J89am4VtzXxfYx3XhLGYJjlp
tQV8k3fr9uKDT2Kpbh8NqkW4pvp1maU+MLaZgQAnWschPCdFFXnHo01uE5OSQj/Nbho2hw8D8tny
Yk7aDS32RFstHCtyU3GFuSKoUspQQ/gC/QBvxCFRrdNum95RFOgE0+FC1I+HhWcOI4OtIGBDKPcF
AMemJFG8KDIA+9p8EY36QTNY9NQUx7hV+n5AFSZoJ8vpdIS0pT24QFt1uIwOWeRtaiUUdW/mBPnR
hWq6dgQlF3RMzyoZW5nZ5WtQDbVx7EPxdFHcjoDhu0fjoR1+skWKyNAI+BXQzidngGGEbkgJmvke
zU/jJQlnIjXw06su/KnINQjrBTXI4yE6ySpaH1ybOlLsKQkJvkzM08J44wCyf1e5E3vD0li3OWmI
Yk5Xd10V+dAMiSVoI4Tj0BTYRAVx8zevWF1f2D1jYSFZnFplQ3/EEOuZDqR6zMXGVe2/vu5mWYTM
edI6GVHrWfyYAcQh2LJPXeTOLMMsycHfrmh5t+/FGaNv9p6lxKhzqtorTQTlihLs3YYvWtupA6ck
Yh0XxLJKBrlguuUScpUAdzjs2qKeD9MO0k9fnqCWRz6XyFJpZRQiCec96oGT11gIAzt9m9ydezV9
5FDK09ocLBDOITkmfzO66ka9OdGIAlY07OiWn2CdXEjQt9oFRmhwOHGyO/a0kgB4nalbkd2tYW6h
EF/ecd4TNyEGOF6guGkQ0G9LK5sdnnNSQqtgDD2uIh5zX7kikiNVGDNoteyLWudY9ek+Ml4HXDHx
RyT8P9TmhzD5D8+SYOwx6ltxzM9p09fhNiTecPySvDQm1epLRo1JeQi14oBLz7rxQejjV1L0Abrg
cwUHR2AVHdzSMeGdeKHJD2aRRuMEhESH9d1gVb2UbGKJv2UwYxvPJzuLKnQ30YUkRqX6px0PD3RL
sBFFzy3wS+u2LCDc65NoxlKmKRdwo3koB5uO4vvs/pS1aNzVOun80KkrIwEmjDg3YYcC8s9cxyke
kfyldKl7N5MUAT149h4aAQW3RcoqeHMbYWzwHq71xRHK5q2gT2sVBhKZDK5SIBh94c9DRhEURmNM
KVYV1VYvBXXgPJd+uK/y6FD7tWHO2mfSrDMEpCrQ5Bi/DlR4Tm6rZSVgzo/dZYgBpDd29T8DZWHf
QGeXLYU0OpOFA8jrE4Aoh1j5i7CzK1FMPZL4nmyLR6ncPCqxvMYHrajpGhorZ8k7nynwMoi7W4rH
0qXQR5ym8KWGGkMygxzbKSJ1oNOj3EW/MXrhc+haYNLzd5G25cTK+Mwae4nKdzPfQ/RSDGi454/1
r+1kO5ZODhXVBEAQTnprah2lC2MBH1rSN4UF6NoVK0tf/HBwbso96XoBoADYVJeZ9qxbM0YdXs9x
npo78RpOTn/wSVfBLbC92KLfNIr9JD8+G9B2LhaNUiarSDF8cNUX88JNc3HI/Kvcm9DEKbuaDJdi
FMowwFFmr9ZyJ3ZR3XmsJ+2DViTSeGfNLWcdb+5gdX05+FhWtarGJmxFcQk3XZIn4/u+WgG3YiH0
iKFCCOThn+niJomO1WNWK3qPiC/Wd4j21DOFR0/tFfaEueVGJ1gj0NAtE1fyPj/tY26lTdFjmacp
utKDGSLQwdtqe5RxLKTTMB+DoAF8zl4cSRa7G79aWy5+I/KuDABFOTsdYVGNbinvMM2QmLRPJfH3
A12g0OF+6vIqlVAW+yQnLxQg7rXq+6O84RHH1/5CnsO2+BeeM3RYsxVcD26bXRoB41rCV3abVBZe
yVRHhWhacr43ayVQpAaWIyVS77X33hAcwaci1jwBxw5TMQU6Wris2o7maUaO+S1ySFEmiDqWJotm
BTw9z0BCE49CZQfRt6x3MmaMxwikXcwI3sLBzvKUWQl8e+3A+J5C7ins/SRohT+M/ptAvaLI21+Q
AjmDaLBcbiHcPf+IkNRt6+vbwL7JCe9bbZ1nb8gyUbtsnTNQtJNLRXykBlYiSIg1a9T5VXoMfBFp
pVsjvGkMoTlqnB84LR8HeYBRC3lvJsfqSyRv5fX+9zXbQwHELhGVMp3BLRUh1GWug20TfVQid9Ky
CVOSoYKoVY+FyiD5xoViKrp8fFIdqjg5EylyiVPHQyW4WgkNurpiGv73PBaDJP7cqDXNz3t50lL0
gDPzXeKYAXPwyEU5EmoJe5hY7BWG0hU05cxZooibsNo15DZPtRFC26y313eHdBs73OlzPRDIdeLg
a2cNAej2i48xR6RlBCWTBHJ7EdtkjLwk9QxeUw/5gxk49i0T5Kxslbe2gqqay9DzVOswT7cfLSN0
ahgVnF6I1iNoP+yMMq6G4zWAFKmCprj5IExpw686zoDld2xC79RqifvEH2Chi7CltVRVj0s7tzXY
rv1vbqOnziS+chDStFeJPzUtSuJalZawQJlkszteuCegaL1+zmqZsfaUyog3MXurctitTgci9TSQ
8rwCwE1bV3Yt+iGZz+XdNPpF5N4KPeYdYYoXgEwZYC2aCRXzxCXxCVGF4mfxsO5hu7NuIv7rt+B6
+if6L8Hmgji3n6sNHaNglbEpn9e8XDBq85Qvehg4w5iypj5OSp8s349d9OGQDfLWcfiasl2YRqWO
aiSKO7Mj+jgi3rWsmo9wyijiI18t5cgD5ABJ5aJCTLjrNpeMUlNWD1v0kjRdUHLZfx64weY5EUk9
tVmObL9ilZmEnowO1BDxn1iOx140tD9Uic3B8UdxOBzkT0rzwpc74wZBNHH/3lO9+vi8FnJ3WjJ/
CYE1gzH/AvosBjQ0nnfDOcqmhJBF/vrcDX04Hr9GvZbgvmDlQ2ACi/rPUsMHD4fo7hY08uR2rkmx
boatzMA7lLuhipYBr8CECJUwnuNLp2BY6mSW4/LwyqliEWSjsaG6rXGSiKCdYdLPqGQVAqhq+fgY
M7U1m99q93M4nsUbaxpdlXQUVW6TzGd8SKcuee0nEBZmHHRj36uoz1kpW2uTXBu+aseLi1okMRAU
LcZmkiUCnLhumkeS/VQkDzMMmwNxQdN9pwaKRJyRU9hvjyXbYXemK27k8jZ5QBNBfpjyS96tRZlx
R0h2lvDEw56HYy3aF/HVJtuKLQvWvdgptdpmNEja9IfHbIiX007iZQatVgKJRRu9T5WswrxfgCB4
p8fuGhdAqQNEIUb9hAVbJ0A995GZ5qeHZgFBXNLH2wAGenD12XjjlNU2cpOI5DOeNw9WBx3IrDBQ
u1BselKF5XQ1rK946M0yDoe0gtRkwipGFkYXETnBqvPnbGLwHKAxfOYb/3anJqHclZU2jsB82ftU
dUN0AfBgFJZHfGy++wApPmlRfFQ9RcADg9xpk7vYXuVnjA4r4a+0jyXMusmG8UxofLadgEroW7DR
r+MltfiGEkzgFo6EyyLnZW9S7fzUlXhSJuY1TQZXjFmQ4hXRXzWZ+Y8SdS/YJLNimWeQ00cNRX6+
nkkBAzyRqQPcGv4ldi4nIqV1NWCrYBSYlUHXt7wC8Ig1L64cgM9PdAO/iT7mfZ7kOWZV4EPkwmDe
G8xkB7nfeovOK08yAUBjJMqqjodOmJ+KJHdaXxVttgAhfqrUm3kZFYSatgWH0lfn7zpB5I+e4ogN
+ykI4vPR9BeoLdzA3sO3rwamugVtZuDarB2cfUCVWbV+fjXRLV7PVAVo4MhEUIlru8XUDPAtNSLx
g/to6Gpy/wX3EMEG5LGuNX7iO7e/6iFaTZQhAt/xzNITvdq5Fn2DDOOo9iY1mgXEL3M+3ZG36Uo9
hmcE1d01Ywc2hlqAbimpwPiv+Bv8Cb8U4Y7oDCpHZL4ZD9OZd7eCc8YDkFyQBpWkINLJAQL5di40
z5z1z43mxyWtQLlt/1eX80jcv3Ng+OEvswFSLTQKi3BLurhLBBmY25kygTrhhzK02IN53/NYiPIC
c9NeKBXHGddN2g2K2DtJLk52Zq5O6uCudQ6bvpSoFZqDbh12PUHa3gmvNFmEj5PNLwqAo/b7gnm7
9E6UTz1I0XWp/O4DOSIktKbAZcYCqB0o77jmiSJjyhr0nW4HKUEvgEGELm3DGJOlOwGt+uSKgqeq
EqSCuqLNYbCA4JirG9Ursu4PypEDDBtt8Yrypwp7tT/8DKEMMjfY/EQ2tnbFqmv7rIUtO7pFqps0
QHT/9Qw6I2pEsGMWbvt2VpZS219f2G40arhRx7IfuZE2TLO4H6UsOSoDQuzRt0+zbSxepcPSaZPf
lsoQtMEDQWS21cLGdBBaP/hXfNrVY/7F350n5FxaATNtLzXt4fhwVUXEoEITSQbcCiOS/Bri8rcO
QYN76ttLyejtKrWz23gMGKsUE9QoeVVocfwBc1gdjXp3Fwruc2ChkcTZrBbvZyaFXhVrOpztZ71T
PRdmmIu+mB4JeLmSD/Ckt2Y/XZuZV6kpSd1L8/Tf45UPu3tywuwgexTAprreDZH9zkzRdii5YZE0
LCcARxrG8xQ85zvKK3yZNni2RiRlI2sNMw8Xa/JTO3wtrsp0ZKnrCVpveCz8ozMHl8Lg1vxY3FqH
0vBVuklTAdtjmCsq5ULlnhq6Qhxr0S89mrTc6xUn63HmPJ+A0c7z8GvoAs9btWx+xIL5vww6liAV
Z+RUuCF8mSw7kIPSw+4NigxYQOqUOIF60Lj4OWbpTIZFiv6A5BRLEIm2YDu5hO7Ce/+C24dG4XGK
b3NDKKi4x/b0PccjGtEe6NRwPCjskf6tEXGLWoPv35/NH0AcE79Yr/L75i/mvGNbpdg7tN1rNlSi
VNejFv7+gcxfNcxWk/rbNkZIRlvMTsTPkWK9VYVcbctSBjz8gPxj99EV/9+eo9ZlYF7P6xH24+7z
EOccXRH6VHwgftwdPyMXJhlrj0LbIu3TADHX6usN70H1kCrUpVx/08rSAjAl/g9VpC8cINQ9k4zg
TNOBfGJ5rb0P8Vrp9KmAwbzWkRsCxgA40N4ShimZmddUv84L5gnBB4EjB0qJ+cBtG07oebZBHAYZ
wh7mZiEFDfwXgZ0ijQaJuis+9wxGccg2en4Nnp3gDFSOnL7FKyf7IE2meASYhZqUVK0+7YQS1R4I
uPPMXpyPspPABH+AdrgXBCNIE7j3xb/VW8cDxCJamqR9D5knnhXRO/q2O/a2wH4mjPkf6UtHXu1S
vEvYBXIY0GashBfVPK0xst/Qxf01Np7zdWuYM37Z3B7niSMr8ZGDjQ1dNdNHsyX+cZd4+5zYekAA
1qoRTTY8iMiPfAqveIRtaIqL7nkvHYGvYwUBOIBzYcrjoHXoGZg3RbqQvvCyjlweM/X2Bw+N+TEL
Bq8OzqeiijW5csGqCfA9SNaP+B6bRuxTKpdE02uAGPQH7NChhs3sM+xyJ2G+xFQBcYhDLHZQV1ej
G/ZMHvWzDw74ndLV/jLBFXrClYaLsfELpiTFpE4yv5Iu/l++2ynfWB33dxfkCs5CNO2iPypqNCqj
0cWJcqROFw3dKR+QzajP6TzyXCVppLcSosgJ9lJlCEdSWhpg0koAbG2f9KrSvyJvX0OcJFByJ3Hh
y+Gy/+wMQErqxXlSlZup0qCEi6M23i4MU1qOm67sWkOMhHTZTTo88kWuErjhBzy0fXUrCpdZ5dCc
tLMy6D3oI1+KnCkQSoaghY4yCRr9S2ysFERxDSOeoF809ack6quXwli4m5OLcPziVc1xZKEFZNk1
4+gOYvPaCw4saIXIhAL97haAUTZcxW/mVaFvZ4WGWd7syJ639TzEddXD/PwQTX/w9BAEolqkQ25T
JYkTN5pfgMc7qxqF2BoNqPjoJxUA7Pu1Cqo0o/xkrMdZb7EVHO6Hp5EVlE+zUBKmGZbEaK+J2vIS
OxP5XLk5I35A+6qRA6BFP7nH5tIbZ73JM29V0d07dDGa/qkSU6Zg2MRnteyEnBHu2v5Rrv9KSCrX
6JU3gK+SapMs9UnBeBuB6e/3dhNnt2KKJ6twD4+F2P3DWcFhJPtnSB04pNhPsGPEklxI+JF++W33
KhGoDa4yWWa/GCrSFt3466esCKovTGjSAPyENara9yjcpJYWIKziSgqTCQWraME+RRgMrRQBcU41
dz6nH3A5ApeKZZ+JOBA9i+ixj7rHjYwYuV0Fn3kcRN0HNS1Gk+Sw7JOBeFVY8QkT3INMXxF9XBTU
2CZlqogoFE2QCO6H8EsBGvCONfCeVIvwJHdNZBoBta/CvljVfZdWwI537zK5+6nlOBWBBLBiERzt
qibivUIGh+6zNmLDiXW60C+8ZIwO1iM4h2oJ7M3B54GuzcRGIuEn8CXWM3e2brsQH2leN9TnJO3y
zSur+W3ZrJfEf5Asa5Wxy4H1/+FL9INvUVNftXwpo/Pod6ige1Tf6HxrLTtwOJ/iHXJH2fyv6bki
zWTG1465lc89BqUYuCrmgfMMhYNE/0G4x0D68LOARkY4lNi3OTEnu6vBd6AEymyca/TwiJwZASGV
2+XKFOyx0xOZ4JIR6B310szz1L0Ix+5dQFTwdwtdosvu5FBXDI+Wi4fjzO/5YgQWwSZIkM54EO5p
xQdDsdGIL3adXjs7DcSHIDhWoieKegAelHgiujqHJOBBskWpSwfWS16f/dILCnD3H57IeXXWdONn
8TmBhWQcSvxEtiFFaCdg4Q7F//M4TJbaAvAvhHHdUoMWJ1HmY6cJwfZm8fuQ/Z5QlyFbIy4a+Rg+
aEPz54paA5F9cWz1ea6w0FizeTMJnF6b4iEDu9qNvntZbO3QoRdKeP1PS+tkwDW5THJUamUEwl0h
0ihHmY/zNFXe7fU8DDAo4XGYdqN2Nyue1JKpstD2lBh4pgmELhQX6DBrjJN1D0xeRqJcmSXMfIRE
k8rUZnoRNs3pH0JCE9xRohSjSKgi8NMqizAAWiU+FI1WZLTR2MVQnbJrQelK36HfG7e7Q78bDoao
R7HsyHZrm8rCF2HQupIxErtTNqD3/tQOuheer0S/wBUlsSaTJyHK95e23KN0uDHuYf9DvccLizMl
dHF/56oV1kBBrT/5MRBv/sutiOjHIM84Kke3r4jVqzGZSg4UxVfYzsHlMi7FGOR6YKkbidwpfecL
3iGTEp4aRUwY+E9VUASQXm+9mh+RBH56n0QmBB3o0kSQgG+ONGSi2EGQPonymzKawUh3NUHm5Jsc
Qh0FtxzYsxdCTuxT1vYG1YnIWE9RHSutea5SMNDi4RVW2xmxyxKuNOMGj+Iz8dyupdozhSgJYnaa
bfCmQ7OoqNjwtN2zZlOyqEixJlRi2t2OdSteDmcI/X7go6tbMoRm43pbyuZsenomo1kOgCFurDsq
Xg6dNN4XOX3vvCJ0LTtEC/d9PhLLbUPeTA47M8IgcsxT3Ov5UgOrFtTriC4UFPklvleZBIL1nQ98
1DOk/OsYpj6kZMR77xMiD81UBOkfOuo17P70/acgXB8+FVTYG6K1zuOFMVIqSkBfbPYsuQSUmte1
2m4iE+AK83IipjJgibOZ8F5RQai8Tqrx6KGa9iauGbKmijj3g+brau3Y0vyInDvDoZddjkH5psWI
sTeXiEcfsvVVAUIir4vWJ5iTBPfJhGRK+2Xm1yyH1QEsk+36BTZZ6XJxNsVjX6+LmHgBnyrtm1RB
tLluQLTBoWmPU/y7nHN0KvkQGulxGmIMnMEVVqq6YMM22qWSyGU4JQK3GTZNQj39qa0SNFKcA6Mw
tj2rfrnG0L9oie3gJr1VR71OfSS9Rd90EwwdXDDXCGid8K5ACj6AOfWxXFCcPJm2J3Ue+bXjRNcM
w+EdlC9l0+K0KGy0PAhqvILbwxiJRbxA2vidxG+1SpjOiUkC9KxkBb1wIN/J1cBeOKdVKRzlBbG3
Tz0shsPik+vUyLmOoRuwxomDwhouun5kw1Ufr9GbLf8oFNBloN4yjsHmBv1egyOLvjPjUe+Ajfo6
YYnXs/HncyYEFCgwIyJRNS6cRAPoTsZYgX5f7cGFu4VG9BKrZplyN5lFqYm8Mquph5Q6Vc5Sifeq
0LfuGq4gpNIgI7KdhgjjnqbrYRacGpAqMyLsimj1x3n1FTxM0ylydxgyLYiBNsIuJY2m1hxCgueT
3yKkagish6Ce5XV029iLW7wUwyHhNGI2q2/rG1G5zOPYuqVOvm0j91c60Pdn2MEI2p/tz4jwmZnV
0nxrpWfwHBbOoCh30DjryMxaJGhXr3AdSyuq/pWmx3p8EjRGWULjwhvEm2HpUJ6eEwAK2hNXFLVt
JojwwY9h5cvLy7XPunlDJhObsQvk5wZYOsLKLKR5YaZ/ptTPxsOGzrGuBhtAaBAP6b3l+8zdUMtM
9fjbGu+j0etEshJFCKVAw055cZl6SGcf5GH7nIS6l+VLd5bym9VGGpJFAw9h/Njn2I9x/JjIpTwY
FtKIkbJeExW1GL3DypnYfU439VOH48/6+VzPoF2QgPwrT+cFhn/x1xFgFem8RFgPM2n48bSEIc3/
o6dAG1qsjGuN8g3CUKVyhMx2RnM19PYZ5jJb1uXv2BmPt6XsRJoCREntukFT+/PnGFBI02/9BQ0n
ef/DgD28WDItbmX+cV37JluJE+8sNaSoOa3SCun7k7j0Ai7Lo9tZ1VTCuVRDPNIZfl4bCr7Ra84h
SQJfpC/2iXCvzSGG1doWKR8RfZLFeBkgmZqIa3AJNPZ5WP7VjdB/JOZ+QqXANSBO2aoVuFD1TL8o
pmlYGhQFCDiaxNz4Xtd670k4ACGDTcanUOPgvLK4vko7yBZ3Ijbm88qVeH8R3CE3hhesfwVMv8oG
5uUQZ2R826ROexknCde5PXpbQHViF6Pnov1KyP+SHcVHbZiETZw/jQ5P43+U9bp/gNisfRgjJOy2
kfqCjLIChO5Y3dQd3aj34dR6VFHJCkvQf4oAJ8Hs3wbNxv2rpvImgthspKpYtz+l+LCMkMy3iEqg
wBPljdYQO7Hsrvhj8YOtZc7AT19nVz62uSwZkVCRuBibMognY1S4ey6IHsLO0Fj+3dy1AsjCFdYx
UKkp1DedDw4AeXZVolDjSumWvpw7eY/2+Vr0WvAV7IR+bleRPPHE5Wphbpqw8jXEQB13sQlwgIWx
0fRZGhfdvfBrOzYoc3/migUe99R/AqGvpN8SwdyfXdc8d/MujuPYGpa3q4FkQlfssvMobn7ygBmO
Fb5bcWekaoccqVY6GpAHL0DCjV1vXUtKy5jUc7JF/bpXUdqk9+zuzatCycf1sznkuwhjCpinxsdO
7mITi/yXIe8xB9begaoDdz1AxdfMnc/6h7enCuyif/jdsYYslB2WsxV7ohmmaI+TBQPuNphb46ud
Qi+groc6erBboAH4GVktP1qFW0I1pA6psvLNqI2KAFyEyuh/FBEiwuxYziKunh9CaXh8E9ncqph3
IYG8tuDEBJHNyPqcUqiLTibyOXaH77t/IBEW1OVmoh4VrMv6O7/OOJjb05fG5IU26J6Xqm92kRwa
lUlJmD2zrdDUrhxJMiZF+gzrse93Wii7F+F11qdAceRQ86MPRHCgvCg4ZL4luT8xf4GuS1EhYPex
6B36STBgTeIRe4o1L3u7riUmuhiOo6c2p4AB6VT5sqIACAPNa9ZH/2ip7QsWDgrXOnKXegeV0waF
fgKvGwITf4OddTVK6FOkFK1rbO9KhxopJn6LfI67fglzABdp0vNeFHViyL+eBz6Uu9GhYjwPjdn5
zA9PX55IVAn+CPIQiQnLn6Bg9Z0IsQYOyXZHLGcusagceWXqTOhncFX9/0xzS0BCtuMWMjEZXsmJ
0b7Fs6c43eJPuyuRe9mSXGnma8VB7CNp1ZIn7bLmV4Hb3d9PzFHmCf1OrgMkX5L+4x2i7Ompr+HV
wK/UG/yFR/dpI2uzrAgQkTPBhoNYsOxYlRYcAdChCIJ6k0WmPr0nHlEzH+7HuZZIFg4GyFz8QYmW
1g4n3m8ADa3S0uBw/dwhR20MVCkpux14uMu5aE4iHE3bQgsh6kN0GX7w+eQajD9YF1k5zEbqPpbE
44ZYpW7xkh/bjFISuPsbz6RQAotOGm+SdQjAHsj12cmY7kXHdGT9xfypnxiwvFnQ0kR+CkvcAeR2
Seh8iUi/wROD7Pl62Btnjl8Aw7NVnnGqWesO7z/ySMvHembExvjGjP/ptzxc2XE8pXVlFx15Ktvt
FvJaQIJHdjA0rIc0tLn+V8c23zQWJpBuFdDm1XVmrXcKfPQKZoMbv+OrOBVMX3T5CPKWRaJIzk8G
wPAa2HIvSJEPLVNW+ZX3YdaU5tY5V31lq9+RAFMAe+JGUxem+W201XpaDzI5QWHB+FRmTXepAZ/M
juG5qVFXaYsPPUNbscLKMd1jmVI+hOfoKI6Fn2D3NnKRbqkfJZWwBLYMwo4crIb+NjeHb/GeZ7UK
MEjlAv2R6UXQKEQVhgiZMBnEmxsNx3xi7E51/xN5o4eKXRIn2eiCfXvLmrbssfTRP9l5beg+/Z4M
SQMtq6GdyKI2UYjwAtnS/y+l2hJvgeRwtVrWVSY9Dq6y2q49oAocOa6KnFJ0xFoUqQ5TqgvXFDYz
yICxe0aO+GUkfnkAkni4bAYWUSDHASv7OisiLSbufe9KfgJURVnZFsW5lp60oLMFFBMYt+BmgY0R
5fNQpS4rmYstO47+ckcptgYS7AgglnPX7T2ZFI91XkFCfJgJG4qpzvOcQaU/Wf9KEy/HVwbUTAZj
su2xHWbS9Ykw7bO+wsktorhKW1ifN8lM8fwbYopdbzdBhzHbtoZJRt88hfbOpP6V+xk7uMChJ44V
ru6u9mJMU1LPlPdF9C63YWGsh4DorH2MHasIynAmRfxm8ffMjzQZNwC4qIVzuj3Z143uVp2qoS83
6EF0Bm3P4bT2vCTgkWF2unkj2iVD/tOqBqtToVLZx+HKk9KiGmBVob5q9QE4eFvsHoAyzVnbKO82
X+bngfnY9UZ0uuzCQzDT/o9qGvdcELMVoTr2Ghk2chkLayhB25mrOtG+gJHSJPDn7bGYYRecQNfk
xXAEgbv5Hj19hQXODd9/c0Yrib0hol2FDEmosHbifUFk9Bo9wm0lGGZx21TS/RxVFtU6aiAMyqQ4
BvoP451JqlIqpNDRY699yvpURnjeHNB4BSWttLhsbEvByNgPTtD8RT4HtPNsFha5y6Ia3LlBqDzy
CpTteHbBhzAZrCCX+n2ACbj72XYL2GfuTuVCqpUUOqUvdcR3WLHE/iHPQsXCFL4NLfihwIjcqARx
4IUKcmPzoWmKGHGO4M0e6vCc3/ahcl9jNlSGsb46JsV7m++IggpHag+k54WQd2JTHdUdRiE1wkiM
4JWyg9bvbkM1wrcuZD/O5rM7Y3x7tSRKihqtdcT9qYod7+Rh7i03XVAu7sF45TvuD8eFSap9Z/wG
rJcBrNJh4fvLJ+fQHitPzHgI1sMZ7KXf6hcgsPUz1TIqmR6DQp+LcDpOeHx+A26P1Dy5+EUIQ1PK
vGUcyPPyZ1GgUyMDGWdFytIsu4/wNF9W+ZkRsczQ+ORSxe1vHB37lCT2yhEa9DKBUZNr2CnZtAjY
G+hxDXywSCsmAJP8e+J2dFd5sE9jbELLH4e+N03cflsIBVe6yqCyg2QqsQQQqBi0evO0UM59BVzr
VachF0JCl46ftob/Q0P7r4ljkQgrJj+fQxGCnCfU+U4ODYfGJH9JZz/g1XHMlWDIfLg1Y8bn2ORb
4zhG8Wd/+CvQNMcqr4FsPTYq10S4K0jFZE73VcxCfZtN+sVQTSphC3lBeZBf3ONNJnXKapkGO2c2
ujR8w4k2UhOrogO9a1uTtRydvUxB7Daec84mtJGcd2vn2THcZwOTx4NblfcPE9aV5cGe8EDecV94
8dcc37gIUEs6wtoLZ/7W7oEqU35wZrgo1KuzUgbCTkAQlnOb2UrEMfd0Y1yyTWOWcgVWGJAsQekc
I3rIFxsPow3nDiDe+wSMCgeq/cgKav1qRGIxqQOtPEFIrbEKltGdK0+9S0wZoajOGhoBdFbJ+z5+
JjF5tsxlFtOQVWb4I7gVV0aI2aYWAPsJo+j7wj5fx2v41UA+BBFZJ1oOpOJNiQwDMFhmtNdETlZ7
as1hc8xZHpho967Ec3/QyOqMJmkqnRJjNfnTKBgW7lXFFnxVbDBs9eduWUpOhtU3HSBnoon47jnC
HBuM8NsqdGHVpIBmP/+8LLU2bV9a7NMd54Rx+EofiW/mhqOeBIADFfemVF4n0acBk9EDfS3jjJrr
HMOve+Yl3syuvBMubZ3GYhKoCbxjjVszmbDXA8WrGZcLpVAXg4i4oCspnD1v8EAquNR9Z93FhuC4
fnJ8fKSkAU5jv4Ia8wWo6XcAEqz+lNjsL6MqZgiZBWotntxcUsyrvWyhDmHr2eL81Iynl27w8lFH
UwMhdHh1igaKil7DL6oG4oQcLWot/9UsILFewmeY8tZkLDDvtgbR+6zlwYKSKDnfrGBnpwZ4MOyg
IYTRhfAmeEjcydugdObduFF+1lS2lC2e07XYntLiek1fVrMdxGNJ5bwJa3bujwD24y4abBcFSM6I
I1Y9pgk+ufX1ahr0qFSa1Pa+xPTHCZdrS6YO/oyM1s2jsEWUz5po0DuiiTBuO663eTR/9FVrOz4D
ITPq/PNS0gvWg6yvrmCx+nd5Z/hTVLyBKPnV6AeBIvK2lq7fj7s6m4EFmuRRR1QkgqVqtPFT5b72
mllkDmtJI5uLVRWVtqP2dTwZXb9jGVy6+m7LEy4rVSnMN4GK3r/sSRkZzr2VI9fCfP0vUPjf5rRs
cMfs/+NlneWnGowfmbbM/DSjqaYAPBZcpzbB3MvQP7nCrjmKyNrkM9riKJGs9vIzUg1ar/cjGdz+
BSVQQJ8SczEgcsYbb9btop7pn1kyt++kqEdjfquE0uhL7hyw0tTUlbhXBg/ys39qP6easE+Srwit
Gwec/By32G3lpHhNXsPGm3B8T6yb4Li273zhAa4NIe9ZV/NAzQT40cHBplp/L+vWqo9Y6e8k86Tx
dUF8OFZsHGyTXkFbNcb3xXj5lZ/9U5R2MF2JKNXrOkY99ObU/IYwX9cVoIkzdwglFuhNw9xXzPOx
qWyQABoOUnmNw1rEwUy9Q1jnf8RdoFYIyMIVeuLkBIHaVcZS7PBHMPoihCG5ZoU3jmruDjDpr5TU
iaot5Ep0PL9vJWuWdBgSM5ARs8B1qjTj2f8yp5ovnobKq9Z6aRZrjy2SI1Z1EHHyczUE1eSaBfaq
DdVfqOAJ9WpesAkRCEH/fAsa25V5E/cGPnLu1eOQJJa3nkTNr8UNELyPdOutdbrcRnQvnAC8qXyD
D80e25URWXsUUVlwyqCYIAE/48Z/Y4Wtu8hC+w+gWcqLshCgW0xotV75yEaDuTc+X1/BdBC72HVS
ZbrkyV0ys4fZfIaXfQ8oZnIPRtOxlq4NgqNqptwP5z/RxatdloR/THq4VqyPGBfansRFG60zcZ1d
fG6WO+GOYDeub/3gHjj2xXDHGufb2EnsuHbFpmyWI15z9S5e+O4CGcx6VbBI8sn1LpVH29tCU/r8
JkNZ6RDCEngHK4CkR4jVc4t3zeggQOq1t4PtQY24EDHwzXNMRtijfl1QYT9F5IOPiAIF4EpUzy9g
5Dn8u+g8DleANSfmLo50NPCioBG2CVjRWqm4FHBlEWfm23CLPCi8MCG3KuWucbN/yP5kbypECTXu
seGVLSxk5DIThthBiLhysJo8fv6EtnNa1pe639JrFnUlw2Z1o5UCzaYIh64/PrHHN3QpMUCHmwlW
IBDpNdUzPaROwraQugFuhWt+aTYVM6otDG0mmiFPacSFnY9GZ7XUk/gN5ItgO3lPBMN5fE3D0CWC
AhSArhPzFvwVR8nJ/STe3S2vISOUTNdNrk2egTO98pMaNM5Tn0vOQ6fZTzix6oVPT4Wx0MQi1m0m
KP5hS7CA0dYhpgWkz4oHstcYdi9inJrG9XPXtAWwmk2VM6VAWkW6kaK4jQa7zc6Pl+iAOgRU/fPT
ycAL9zUM8uvtwdxcku9AZ3PfLR4JxPe9+loELRaF+Jzbv9p/nNpLdmFMXKf4hPKbo710WLe+tL9T
V95uTbP6+rTvOWfJWRR1PedM4bemqdhT2AWQ5E9opEb0NMd6Ok1FPe7HyMF6ElWXpiCRqL1Mz2lR
WHOQFIHdhnIyMoUgX2ZTJaa2+kNS1iYY14za6BYW3wXRrT1t4Snt/ShBn0ME/RsLHyak6HoLwTsU
T3qK2n3OaAPj05TGcQ9HklDZF0AN7+4JD7AbFz4DgXzZsX9xAX6oIFkdz2hM23m+brUdTfBKHbMc
IRrsenK/KD1gvuekcm8PUhIoWDJl2VvMNieLGOOoHkeF19wPBWY1wwMdTEWdScRU8EPt/tk9jEQ2
EU97HdKAXMCsMZS8aPDSnmQ+j6Q4BwiWZEU7qO1TX2gRG/NdA1eOWXAWGPXTqEOGrVtQmfafTPg6
/B+XLGJ6lyXWeBodMMvKrS55oqfIPYCRHU3qLBcyLJe765HOjguUCIsG75pEBmF8XcFNIg7PXJ2i
SKaC6MBxXrvRX0PHXfPf4scky6liFOmWyvG1RO3SKVHFaOFGuKu79k3u4dNQ08v0AwVOU/4ph2Yr
heNMKgp9JRgHoiZC/aL++i7KKygNE7G2d630qdTWLjfc354LynwVdgkm1JvVE060cIFAcxco6Hbt
3VV4ocmW5+lFkPztX/fYSfsAfg5ou2D8VxUKF0WkRWuYv40+Sq3uxr7rRnqOtMN8cEodML3Bx/KS
J97YQ3HiTih2z9ZEmiYdp/z4odnXYSgIo88zywuMWsdBVV+mHJyZsbSxDEiKrtXU1zw+wWc08M+d
Hz6QhOQUUJC1eVS+u1k7uJP8WeU3Bdjqvn2+7nwyhyA8op3FtlBTBLWzL2RhTgpz/UOWaC2pVKaO
WGfIDYM63l+XqNXRle87TdZ41mzy7zUx0b7E0WmMRL/l+bBelYn7uza3B8j41UcMX2V8KG2LEbFY
d1Rxll2cFNTE2Qi4FbEP8O1HTGtlI1mMtRRUiRC09kCZti/AvHgc79P85ABYYcbavQ2xJym9LPPk
caALDAL8hNjsxnkVf/iBuTD2iZ3yPbJBJDTfR7+G7bKhuX1BK1Ljm2yDcI3rH6PC1PL3JntiOR/E
lZoLalFo8RHUShMQSC1wBko5LaUhb2ux1PLZ4TIckRjJJW537HWAFeBBJT6CUUlHE4pKL5jJOd48
WZftnb88WovnaLffZulcT+F8iVrqGlgYWTgGnSbgeS38j5i03I5ajJHOF07IKLRE98fxq/3R7x5c
09U4GTg8776oBbMXn7+hiUB2a4YgrIYBFLWI1q8BuLFxQ0KZ0Eoneadp2HywHT8RFlruJReo8efn
F4/aeEqVwgc5tixnakGvsKJOGRrxdq8A+OyN2FvKKgLaWRvn5wsA29+W2icJqm0JmMXGkTqZR00h
ioZ0jfsIzemmW8/ojcCBdaC1uyh168PGRrumUnuU6rK/OMPUEojOOFaV/uHE1pHBw5DKUCTQloO+
9ZRvyqXG+4f5KNKV3NMjii5y3vVbT7jZqPav2R9EZscXWpU21HWdqFHxOLPVxwKc8nKPOYh4IYSK
LcDB2gzE6V9CvYK5oI3DmLTFLTfw2/nItkYwKMprjq2ukrpMmbclEJHYXO6jBLF80aEQ8s9zfYZr
XtmgwT+5hhhrYbkG5nVnHJt4dYsOyRPubsEQWDFXADfBEhP2K4th7Gdirx0L7cKr7XIiWG1Lv3oM
eUstMp8J4beU41ACLvqJZ9AHqZb9BcuSYra28d4DfozcqR4Gak0jt2IaSWkcRH+K2kxpSG/ZuRNy
Kwvi8F8ujtGVTRdo9XjLM166BaexlxbN5+crhsVeS4JLqy1Tzxi7DuBxF/gv6YNR8HffC/6xWxrz
wIEr9FI029buKo0RlfEhN/qsZYdiXZ+Q0k4uwBDDE/qP5P0emVPO0NtkzcDds9t0zbZVVwh5Lw4r
nf2vGcg3ERaN2txt1RWbbZTHiQIyI9/olB9MMOlggisWTfPpekWVKfuwsYSupBm9RInzUqZTxp7R
f77i4ACxngbTbHR7hwgo3c5CS/9TaVukC9tLkY12s7uKUJnCaPvFRTtxuBmO2f6ET2lmdY0dFvAZ
NDFEG3gmzE9PFUv0QIqHWTVo4NdaffoAskXHFGX1ZHwPA9MoyuJiX7jrTt3kHCjhBaD44QnfTZo/
mN9X3dhnFziH5GZBv6fdg5K4WNY2bUKaF8D4wjG79GC0ZpVE4YalvAP3a9l1GYQ+doWNU0nIjgpV
1sNBua9q+T3E2Z65wXOq5atiX3mjr+0njS1Q8WXEqKbSGf6KuIaPyOaoCy3B9+a5tCKdsFeINigN
9euEBAN5PvH8IF3l3cUEw9uPZJye62+KA58rO3hue5WnX4+jAzmrdC0d4iIINJkbHX+3t3kdYbCL
LtyAOrpTk34yWD10oO62/7+BcMLKokY7AHG876oLRVnAHzwKMPVXHuGM4XJR0Y1rDU1Ln8E4tDB7
tF+GHL68kw72B+HUDqVhGLd30QQVZwv8oMUeCmy2SaIzdRK5eajGXzX9gHvJEN/i0Dd9sfUDN+g2
4Jcbxys/wQx0nuuFZiVuLr3hqqq9caHz4mZi8jz1emzVOFUjYxYaU+n1StCc3jylNSsN9o30GqYJ
ST/jCGhNKoci/vKbICdjb/gXthNYlGsF1MBPxQwONKERXIwiwzZ+Stdl4akCT5EH2Jz5nPY8enus
QbP4sTXYSehpl+2kQV0/ZyRpDKIRK8F2UfsTsy46SGrMPH++23oeaSRcLG8gl129saogyuOpYzk3
0aEaAN0FVJmIup71eSGfsQFdHrUbYbp5imSrAjUwni3ECNENBjDscYEOMrqH1ol3pbZAUlCsZyYj
BetlYfGIaE9dd6/FB0xVWie8C8HSqR90c7aD+YRkhFzo2yqRBCOIBTevn2vryi3SuE/sbrleNiJZ
Q9m/JWld9phEWjkOiR+GMEeYEVuQsqOMquaAZH8Wu08q4UFHyAEEtaG5NSH4hOviyvfXy0dm0ibc
D3gPfvalhnZP463e+tWm5nrL3ejJ60bbGLJPBvutozeSKcd9kwcARENKIkQdzw4sny4MqwRJZeXA
b2q3qPqI7aR6kIQ8O2BESLqf+q1e2OYPlQzslAs1Z1GPOQa9xFuAI+ba2BDR9la3S79Bk2Rza70d
FFT1OMoYlP1i1cqZNAFYp71kDs+iWlk3UYcInJxKyz8eX/XLZnTncc9kb0R2btwmqKEzobRQ44CO
QqiYZQ9aO02Q9WIODWw/XiobV1PEjifL1stIg2yLbJBXKblKXXiywKwCfUUDhUF57aREaTa3EAxZ
eJIA/iPKykMdAfE1zsd/rXi6oZ+dlNpjgk63RrZN50GRfA9eHPqeTItG90Gma1Pc6bbqcvas2Ort
265Vfhk5OFRI8RvuEaf6tCcSuEnL+7YxFlG+qgBsR9gVnf9Gd6IOfqEXZYiOAbYQgPesiNxeSirF
VsaPeBXWTw2h26iCyO86VB3CWBchhjuDmZQn0BPFSirHXMFsnAXE27UCpWeEszKcwAgJn9Nr8PuM
kK2wBJTIC+I2EAlUumdY/Qb9ZipECPTsv4/Nr5wQen5FJwUYDJPUrYsMy6D43VdC2OBgePzRTTVz
9njUJsL+cgAiYlay4DpsUHenkfreBg1C3KuL3nl3R1Av2wTLHjfFXkLxuogb3I2LQuLd36ob2O7I
diUPNmKMUk8gMC14M2ZnPj7xpfJMCyhjFAEjqh+/foe3jBNA54u1j58UJvrrOrtQ04mEh5WkQuOM
xVVU1Gg4myB2wNSeT+jgKWxWt3CyXoeuIpLxOEWBFJNT1pvRAcr+JwZ9rLI522ecayf/UDFfoWpS
8D/7w1EHffh27fKiFvzDDuot2C52HhTrYPSJblWGOazlsx70ai1lnUfDYSFae9bgSUZTIljNn9aA
M6AIrb1LXVTI0vKK6asn1SbRHBZbE+kdrOSwRMqAWGKZyNgiKHDDRMl6JkvIKId7rUN/lDF5wn+S
40vP/ARHAAPJ1nEQrqVQFhb/0q8OO919cDl1++wyqw/p79f/lfh6cWwurvR0zXDDH3GvwEPHWDPr
5ingBkJP3y/v1liy0DIaHV6PTxk5R859sqgUPNV1BxmSn9N7C3wpl6d3A3XTE7HSX0+f+xLyYnkO
Bo/JCLuti2cwlK2+ciBRyMyJkRdCF+glkJTKhZfOXvJYpHywPjjikC+YDSHRUVSQh1eP7AzZI4VY
FzuNkEhlRtz3OJQT2+YuEi2VTRk4EAwkW7hFjvhC4PtMbw0CmHqx27qrIzZK4q5zdd+S4Zrj426F
3WkywsiISUEt+GS7NFAWgIUmBeff2y/Gs/0QKAJHTqFJCCefWi/Zgp82/Xnm1sqtykv34lUpy0cG
dAhQDDkqVvB7f3sTX5hRcwL5kQ5F0DEVKodPqW4hPQqtioLFRdrZGFoRXpU+/x+ZXBzaExOmv7MM
vI6kP0UuUrbpN7pCcYuqEVFn+I8VNKJ0P2seLEUpL67K+q3yq3lymuJSA3TxawRhMbEtmcUGQ7vN
NgdNOr0c2ZSKRDVfoLhcR2+z1x360GpEtNHXFkHXVmuPifZ23cQGC5CpUghTg8Vmmzc4E9cYh/4W
rwbV3Hr3EhjfvZWNmLf5uBUVNMQceOFfo9nz+Iqxgj9An4eokuhCkP0CCoKBATwgabLA2HNHDor2
/nsBkz0gmEr5r+B+uxAGwg6kUFa1MxO0bwfdR325evKzIkeSSocQ6BphCQAE/+gA6uQQmN+NPpp8
JvwU/UUiWynHQTD2oau804eD06djeBy3bLgTh3Bz7kq/lzKeR4qXvRc0WEjvWq4k57fuXHkinwtE
/ZfrzQxbo9wErXpw5GMSYKFPUfxCucGMuDZiryA4dqet0WFlzzd0+a4HBM6xwXqIkHqogBmX+m6J
3HIxXUgtFAoCzwAFxIdkgGHEgtxqxMwAI/FlfWewRn4qcswqAdCbGh2pjOgkeissOFF35UrC5VoV
BVqS8Ae73vuDrfSgOW+xiO2KHY/pVUjuL/H/KPsuxrQfThDoCkhLaRRyxuYMcJRb4pY23bmeQZsx
UxE/OGrgsqm8IW/ZHx6GITHsJZyPD2++HeN6f/V3xNhHHAiKv4vMkhRf32kJvWSpYuIVUrj1u7gI
cY8yclXb8ZlBhEK++lP22v8pdG1R408E3j4s2GdQgIdH1BwNxSlpaRluT/IaMsQAdqDkp5Fy3TP2
0JahrXBHSEg9xenc2JwcVn25Z7xUzz1Whi0CgwWNtfVY4RTDkw9IXZ3gCeBTu3fycI6PjDgtX3yJ
9MnGAGgZVD1CxcgfsQvjmKGINpAp9NHem2qNJjoX5ol4HqXoJkyc2ZjFluaRvDu/rXrWzgNPJr0M
CO2WN+oN73jcKhJZMgS+FLPmUS6FLJSK64LbCgXB5+zdtr39yYjLL+RFdAqM98PXYjfe9WtPzPFw
z+KlSgQtgNc1HCylNUHd68nlIPxfR3b8PxwLoSdZ8OUSaoXkNQNjaQqLbeY/Ug/wsrNTUu2BuzWP
3Vk2uQxN3e4I6msDHY8NhEyAcAcQmby2uOd4/CHX2L20TLtBeTeO+z1VV8dfBugtBC8i6Mi5Tpca
jU53l0oaq5xQ3w8/Z4D1oVe7v0cxxFH6mDDQYXLeynOYPJAHRTXumTypRhAdQXX3/bH3GVkU6WQv
cgN3we/BL56QEwiF3aMuuwHlOh9cO5fQRR1uGIJI0IMRklwiIjCINEq9Lo51Ir8vO5rdQc7pM6ex
8mvIG0VKIxalMCEa2HBeH9eSxRzKdhVK8CpX4zkVEHSorXiWbf6kj6iFAtc1OhjQ8YssV6B8MOHn
MKfOe4+ZfVdnA6ClrsLqTwabi/+L6Pw+T2PgROYxU9v7zzllzFpyeg6uPAChn0flcqkhlFD4igXX
34ktjGu5pWrKcC4tjOkrFegcMKOplnT2EjhhmJ0hBDR94QmUaHMlqzsFEbuHDXo6GeRYlcq7GzM9
LWO4gvSpDkWnojkGbXa3YXX52JVSxg1LVFxrQhjMmsU9xa4XWEKUAQV+zmDxDTWAGD5i6xIAL2F9
jwc3bKOnKnwzX2pm+pNA8wv1kpivldzJ7D2hUyQmgJlx7ygKDfgNjkp/OXcMYWhnIQgPvK0pg6sc
1YeGS83hhhzDYwE2ff1jtRK5QEUHxxdIEm+/j0jwEwvh/8dXKDGVXNT9o+DvLF3Yi6d/OA3sDUh9
juYorvUmClbkJbjaJTWx85SwWl8ai38bTxE8olP88itAbUuHSasm+5B4DipwPriW5fa/kTmQxRdz
8yqNrOa8gQjxA46ANxDBvWVkQC1au5dYmjenjO9DWcMl6l15o4jSMiZ1NZ99SpKuO0XABntu2Z3K
a1X04BLuxbGymO8DdU9esEjpkLwFnAjIoH+QhOAq8R6NMFGLk+HpZX0FGMgjYNNOcFLRvGr3bcze
MVVj1x+LCBBl9zUMrUxvyU9pWDjHNXVPhDdA3m7UnOC0zyP19TzyT8fzPY5GVGGMY2Gzm5ADhCxN
mWJkuUeaHLnahYhqQj+oXNmzobkxzXo65w5+/sP0LxjyAow8/B88uYlwVB4jvtyQ49dbDotUy0PE
YhR2xN8GwjhpjdVD8xFbfj9J6GBL9XtrnNeFzhf4KRnrMSmktTR4a8UWAeTViEL5UdlyWm5elthw
/MbJ8O5qY6RnxDLKIAZP5elg0Br/wo+xMP5xO1qI6MqRrHxd0znqHcMauNuZwGSNU9BhVQkQDCoB
emqTtiGDrIZU3H4ZKKVY2EWnxOZG47/gN0uCRrmsKovp37Y8Kp7fpocuOraNG09vGl9LKORk5xXV
XDTujAGfIocpeH1LhIOI1+4KqhD+7SSvAu7gPx6oVp2OGAwwO1o45IpbEd2V9td2QKTzbBmVVxdH
cgbkaTYHdh/JtAFFUnRPDiw8LdrOmo/oV8QhEbCLQm2uqpqjZW4HX6as3osHxw6pHT2nzF7dFQ8K
frtXsU3ldh7r19pBTOMNtRUht1NLSsfSYnPZLjlhHYn8ef7zelYIB36roye3LxaU3fD21MU6uJAr
/efk0O8Oyxk5s3BAWNIeQ1KFRkatvSKSRFpwyT/i0wlyGbwZ9pTnKYblt4s5h0PMLlhl6DcGGnxE
2R1VfxBNws6Mv+sxMIhc5VZUsxiveOJe/9CE7aQVZns9fSKNf5YwL2AP2thj7tH5RkQ5MLa84zRV
ImrzrwpMyxk9uiT6k4q8ibcQPhyCpVjofDLan6rWLLMa38zRGi9RKhEmrSrB76tNfpKb0X8DoPgw
E+8/bfdk7vLvnTVLUIX1N3qa8n1/d0tL+SJoeEdgQZdpCxaKhJLH5y3R3peHLd5fHeMU7GSUrLTF
pJhbuqzRI6izeCfAIUfGznz3XP4DBxbI6EL3he/h+I1788VoU+VYC42jax4PshYme+RVDQwwBHsl
CeRl+BhfKvRqe5yJdtSho65iL9cReblL7yJ/C7Kdna6ZUWOeF5yPBmU8aso2Jdm0vYJ4a1Aj6RYE
vwnJal6lFVvx2SP5vTFNrNf5/YD93FykES3SBs4E6+iu7mvXK8SzkGVZD2cPbUX0VyiH8Haw3vTK
9jjTsO+iM91f3PJ0FwmOeJPj/YsmK99U5fbNraDE/hOuQOsGu82reJoXCiz0mj7XmmLRnA4nBc4Y
IdsXgJeeB/QiailUEhO1PWDHaqK2ZnF1dI4An3DLFyCIF5ELxxECSQUY+KOqHyxTkNHxDuD3I8NX
eXxiRimyFie+fl81QFlNjbtjFXH9J/VTayTJOz/zWAueJv7jGQccA6hq05HsanhmhFF8ezDcoRTj
Mjz3KfCjQ1FhTrS+xMBLG4Xfu9MZTHvZ693VTAlRuENL6kqKJuQqj636cBVfejHqg0H+3P/UheMH
D0v1FHvNJyvj6ST1YuYPtObGq+mn5eTQ8q2Rh6JN2pyaLB0eHpoz8LTE6eORciwGex/9SJSQycj8
b1sU7Q1cPTgtkXb+wif7z9Hp0tyGwiKgkjHWCDv6ciiYYzEDDb6Ekw20Sbn0Mha9bVArK76DMSrY
VeNSNan/MZOV7wqzX8u/Htdw7Gyqh5lSd1vOxzbdxO/jDEVfxClwqK6rlVNZxLWr6fb6sGxbNdxh
/zIVJORFuka1fyPYhbAz7vHXjAYiqxwBfmqL9w5R4fHIk2Zxc2wWIUeBLYTwyWCeVQeoFi5wG5f9
PiLRG4adQHT7OcA/gtOlLeBQGusBKK5IhxiKZA5Eq4vWCojX7m/p6/i2v9zZzuJB3aCpuMxNvS7c
/SoLCKWr71RLZLoxuq2XIrC0ZZBtAdzGVzzhAq+5dOsV6/6DPXtVK2s6sH616sxFU6iMu2B34Bod
nZVILaj3EgxSRiBzod+BLGlbS57U2G87UTmrlyrueVHXJidnwpSM1aBuDgsgolpqv6ZoOFGSgbgI
q6+xirLTs6GpkhhiiYaQKdBusav9Szf52xiN6wcTXidKpwO0c+inWpriZoh7l+2X3SSDGLrIMQcf
5MHeHQaYkJE4g405foxiOEaGFd3wKgow7ZRsXRQlbUDptDf5dtqJQqXdmUZXiuvuJ1q80rqyjdu5
7bWOcb9cDF/XDDnZNEBXMGXgyXFQC15zp3ihNQiqoq/7z/b+gjXANl3IRdVPWTlAYsXm1JwI32DK
Z7MdDczMzaoAlTXc1h1ihWvQoZ2sJtQwBGPeCUWrhrwQr5RR+oLElq8bS2J19R7NMhj9FLUYtqbz
MTt2ZdofrfcLcsqJByBZDLa+WSd5V8ZvirENJj63e6ICvMfI5Ni1eD/ItFJGLbibHcCPB+PVMp+D
jUXyh5rbC/RcCloqBtN1Ihfp+EXkv0Kcy1zeQWqd52nvkAvtxB6GfpaJe6Wai+DqAPliwPWhWhX2
4uBnyRvr8EfjTxYblGQHRsOyIceq0zoIyvm8j10T9oxUbiEGrpjP/PmU/x+Uuf8pb+VUjmdKFRVR
91wG9cQzTKm1km4W9S4wM+rdMsHAsbYt6blomRm/dFqL5Z8paNuiMS3SGu4uU3NxEACtO8eURNao
H1W/DNpPUtZFPsYAYQZH2RG3qf2vWcXcCN+su9TDZHBEbbZSU5G1tWa7N4jlqa3rQs2LGOh74/aW
Df3vr1X46WQHLo2wq3nZ5TMzL/IGFrP7xyzOBar9lN1g3fakS4v/v5xaZ/NrYvYDtoy/Iv0eGKgf
d5JgUplL5Jgm0lGUDvTqVRHpmNP5az4Rfy4Q6zvfCGPMfJIOZfzZX0DK646h47wxNLafIF5inQsG
QERW+D4EbDlFQaqwE5lHKaFIdGuENmnkRh4vfD8VR/BcWe6FiFguDDuqYwpN9ad61XwJ1Zm+C5Nl
1tiO0Ol5/qqX+Y81DpVvT/OhsZAV7npnSVDvt1fN/VDNVg5ltMlhVStzURdto6krPxI/i+rjaFw7
06LN9mlD0DDPjRQQbOtDJfzzl+GVP46+36VMlbyb0wLNM091Z2W/aV5Q6HHwg27RQlVo8Ds8y5f6
1Uzap5WGx4bpQvQnl5E+vl5Y+sw9+Xp3MEafKsjHNEyHvMZ31sr3SNglPBXMb6m2Z1hXQnnT0jBN
W8j7gc4XFokVa3anpqFfJMs+tZ3S6Vra2e4NeG+uls+5p8nY6KFjhnv9iOnio1zlEZIjvmCO9mkX
w4BwIOrEHn6x/wEzJAnykrMx+5krQI27yyAKXe/N9rQ+W9B7mzu0I3q1HyqKWWoo/zgDHJqNu5sf
T8DFuNzRqup0EYyAlheoJt2lEGYQfkCkJ/xFCrC/fNrz4v6f7aztijB6k3wKbPCQL7d0k3zXruIu
VBprz2E42u+qQgL035K7ZS+Vg0dvtBzkpU6OCFkgb0lQPXWjQ6bP6gceiAgUzJFr/ce/317CPqoc
N7Ay7slel9ykte0fbR2Qsxeglv8BD71qM92azeUwK0cctuncqJy9GXUmdYbfc35hsqLjwVv+SS7q
8qmqNuGOO0waITRuvBM1EB+Aqxp8eVCYuiRczjEU9J2zPsv7bF5w2+ErIi99hzDc7mLNw5CGXhQB
XtfZvv9JEvPEGJIZVf7zGPHy965OlHfyVVpfdlVCeS/LDpBxZFvUJNFzPqSWAkk/36g7wkzw4Yui
gjp+ppjJ5SoWZ9kSVrloVB711vD/RmXdXc70qpfYxqXlUa3OJ5t1Cev9dRiMKo7/E+gsdRyhM1A/
MZN0KQA8REENapXAA6KkedIlfq9Sa4HCdYx2ykv/PR5w1wOKiDjI0iLY/P/9ULYsccTsiJq+Z+e2
KawKa/N1x4HcKJ/7Wg98gB1D+fRMkkBGgoNeeftT4waY9NnZideOj9F2LSISjWWzn4ZqI7c6SVlY
LShgAR2pakfR9ZSqeLZ2g+AoeuRYxcKP78q0/tRYAfDdi5zly+31quOVqqSctfj0+kNPuw2lXpwa
b2JE6WJc7LvO5pgyJx7IMQB1bTRyfWz4I2xbLVM+1IRsHbhTVvKU0Lb9x1k7/Jgo4WxMEmnLY7Zc
MEL9DsxplpKJCrmR4l0gqoMhnJ+ASCHX54PKu34veex+mQCiAdTpqb40WbydvvK/TYJT9qgl5jY+
biS9+ZqBf65F0YWyU+87Jy2hdE5neUH+HJUvaEVqlxZwgWk7MNUNZe8gX4MWG0nXyLXJhJV/83qt
HlXUzGTJo848dYNtIX+45IwzwjWmkzPJxKt1oQxJCMG798T3xGof97AGwn6eW+RdlMEpeCIWZFWu
ah6Qn6xB9Xlu0mA2jTYNA0kb3ueQX+0dAviezrf0R8tqSu+LTNQ0Ywk6hYRJyJroFuMCYaD8+c1A
/agpnESz5KjBVyDyksGQSutdH0bV88UEDR1JewtYFtAzh1mFrZxIRGwZBnc9fQaHhsEpZP2eX+5Q
dsQH1WoWFP7/+k9YyTA0wbTakEJlIC0h577MkGQbq01ODk7I/DsW/S+GzR+dp0+RDpdFlNfkMww1
AcRuMg07zzbKTvhNMeDzTnzteaqIYjYRi40f6u1ff70Za5bhWBPLaQ9fZ3SJa836ePl0+ML8vfJQ
PJY3ZuJtGo6oo21D6AJ6KM+513hSEAP8eJPpXojAZGtVky1trAUsHwPUbB8RZ7BuMB/jb1BEi8+z
LcuRLAOlrmA/k5gj/8EADjTHTRDaoXD4IUZpOYu4HlQEZQL+PH/+sVCBpN03sjbcteV14h2jnyqZ
cvOIHDBNJEbjWyNTDWV6Ik3rEyIBrVR3B/owGqgrZ+H/x4ugPSmn7lCUWAzNNRZ6hdFfvVzTB/96
aBAevY0ZWlZoObdySMlks2P1sZxDFcEGVz39/l3VT/ZEvUJL8HjuuYRNeMfgw5q6NTQe2Qc+au5R
UPsQZElCK1ViDxkzidJ3QUz909Et+ECeQhxzFD35UTcVZ/RjO3nGRJqg1HWqtnk3vz3DBCkFupJ9
JYlooBiZzlYGy8BJCp+4tjkRKSOvvUbOHpUT2+Zj3SXW4BkVw3U8+rUDGo/UquLyYJM8d7UOvu+Y
g68bXVVz9ck0nPQdRdWmAxkELihSVCNuoT54o/MvLUwN4AGiPTdezyr6JauGay+X9SfUDfGCOrMN
HlyMynqRTawAigxFBku3qX0L6aPEkgeTW0RYJFrn/x737P4JSTy+cckyQR3Sr998CttM/d6sXxCQ
Ru4+aDw9tjMRTmCVdFdo5gvQ4yFLPAIZsfDUQlJpGYOoKopJi5LlA+dGsooB/Z67EVjjD/+JUg3c
5Jpt555b3yL5aBLoDrJv0T1A4/w0xnUhVDPHPGWeIetl0yDgD2mbz6qeQbmYk3Rd1QvI/9r+3gNy
B1qiQ+K8ka4eA48wn6pPe08+LTsaVAi99inMU/iocdug3NAhFY42Ih5HTnvi/X7W/mIPW7jCbRHQ
2KyLXystnTPtm91y6ymk66mWiAXbe933wfQeJf8j3YyQtw+J47l1tlgXBkdPP7E65tL8PhMX5wz0
17IkWzOwq47OeQ/psb6pdYBlgbxpfNVUtUFIwkXiQd1OIJELIEy1EiwPOcYDcXP5OuWp44A/54Ha
3GFZF3eVHnEq6CNQNrEmkfS4gdlkIXDGsGq2nD3ypgPi1GrgQ8gpAMxDm4ZvKd67Vr7rVQzqAxZl
0IQ+ZTYIXxbGviWuebd6Tx1i687oMe6tmhjsD9eLEF98JCqvuXHTtLlcgS0BxpTVQipFWQG88Rau
RlJZGE7+07z0ZWAbEUnpylw8Kp9C/5FimJqz2fW93o60r3w1uq3wsjF15Yx4pMzRaRgPkqY9CFLv
TCGxdKPiHkGH7DBJBUstQa1/u1MF9J/6ISBKmSmtEmf8Hut5vRGFMvp90bzvcqd7XlDHcFgNapH6
LbrzoQ1IuA9rrmW2TtkK03TcWND7JQA0pp84CVjb2S2sdV8RRCzaOMqDdc0wMJJrxpb0nlIUi38W
wMr8BH6Zafm7LiGcCykdQ/7cTn4ydJvMg9V2DgYv+pjs5j3zRwMit7hJQ3Y951hVBtOG86E8h0fi
ZiJthOWOzreM+XBteybZSl6NcWO91p+xrT4kQ0ZT1RZ1qXY7Vj6chHPqfBgF/nyit7fu50EKJg+Z
A8LpHx94UPdF66xYntzazgDD1Y/51cOrQmm8uRA3OTf2T+7QCTxgvFCwz0/Hb1fdoDa14aUJB51I
YMenpGJ2vO36lk4ZUJJNsjAz5WAuvH/hY1s8m9tjwOyofeto1Mww4MucETdo9k1J8wSWQz/eE4jl
9qslPAsRKYEOcsx07KHPdOAeJdWR8dxOu2JqEa3PYOCiLrU8fS2FmXMG74erx83m6Whd5+0qtpGB
RTkN4YMx9KFhoTjTl4mQD56Fhr1irz61xtpf4q/ThTYL9JzvO284FXojqoFhT4f7wK3KJWi7Ve8u
zqbJMsTzRACy8Trk1phv3I3VuiHN1YDksZoGGBdOZ/OW6pTO1uIPaTiDRvayU5smXk0xG21u96Mb
DP8acUCaCKWr0JG+d+prDQqzCqKlufZloWBGJ9zpG1lIAiQjIaB1ShXfLEGrnj1OwTNJ9Si6dbi4
n7DgfgM97dbdpgmrOOFc1fBBDJkzXek2Yey19/2mirBpW3TVzBmujbT+HaHVkS66LuZy0OUeg7xN
d8qoZD81OIdTAOtUnoCdae7cYJnnLz8rOr0yGh/C/zQ7LdJyFF9T4WyPloxb45wPLIeMh2Ln3bKn
ub+t1WcmqPPrsr1ulIbjLMMajGRbyqpkMGlsW8G+M4M6mpqb0z+pHhM+QveMKvIZYVuXp2gdt9qh
CyFQTRalTCDTHoERv1ucM96f8SRVeXGYd46tVGNKFaPzgMicDgovwaqWfrpVc9hTJXq/2mrsKZQr
FvzxuXtfxEGhO9uAzO6KWy28nkhfDk9FP/JwqEKDGflD7JQ1QCwn9BW0R6uT8fgqW5TbngrZ6fNG
xMBoH+WAVMJyJywnYwPEDS2b5xmGhJ/K0jrNPWCDftZd6dqRXN2gtGCyzJQekKSx60jdlJZ8KASu
AfAy6OkAkfU8I5G9hgmTVrVU93531Q5CJLyVb1bey5vJ/7hGBeXAb7M4Xu8QXqGZLMH70go1t1ag
xBSjc7L6cShM0KtO6XFdzOPl6MIJPHWN+Cu8kroxrUKZUHunJBd/aXgiq7Dse3261L3cm+/V9fzv
WQ+il2mXjBP6h719+ASta4pdwOZ278DjcQoM/aX+Fneg98nCXzE1CMTg6KhgpxSkD3m5KAmeDs/K
9pHiofU8coo0b/XSlbNqJyG3ppLX+OIrPjpAIbUyB2C8GnutF9Q7sds+RqpEiP3IJD9v+btmGFVa
cPxDoOA3ctPwCpizZJ9aXYHp+/7/qKakMSqd7MKErYOLDHrMSuWrd+Q2nUuIUdimr49REVxvZWk0
Gxqrr5EcC3/x/zJKPCYykHcYM8bx5cEwlY61OZRk2+hz8KxW6lRzZbTUWyB0YdTpNpW+qJgS8+lV
5wE4BixahGatp57i/HpXSXcj91wPKHujdQN0qmUE7CiL14YaaiFmuHQZDBpmXF/Qo5Gu2kZC2yy3
QR7l/Z7ILW4og/D2MiQaaFRpdLYAluuknuj2ZuvsZmmTlqj+6M69SoBOCkVQnqFH510+T4jxar3h
bfsqcWBjlEOdaNKIGZXy6r55w0DuQVidpu+sir+KAmJPeAIUMtDaJxgPMRBSw1GbrfBeq6R0Tij4
NEjYp2NEbUfspyIguLArfsb8/r2t023IndDpKu3g/yhl3o8QdtbJfObCkkbrev73WX7KLJM5n0pw
pBppmRhuEeMJ8tpKE3LjO6hTptWW7DL6p9enmperCGrN7dIJFfTgX3/aD2cnaRIO2g1785KPVFGd
lO2N7oyIoJSqxiG4a0lMzA3PR+fek7k841FCJwBTP3yGiLxuP6UpEDMEcw6vGmzpmxIcWL+C7iV2
5wxUSFw83gnFYZ5Eo+m3jPTPjbsx04vw7WeBBtbHU7v9dJI4cvD0+tSqY5e1HSMdUNf7UKPzFnSA
5x9SdrHWOPCdxE9PM3gnipDwETlNJGaL/vbS71HqqYMuEX1gr90vzur+ATb6fk+F/s4x8eSxyDL+
aaYjmYHMPP7T8l4PCkx+VN75T5SwTNLtO2IyswN8v3nxJeyl3cUvVbj7gsxE15NxEuDomKX9jIWe
WS+F5lLGClPahFgwP3mgJZM1jc9BuMV1JWEYUnuUyKMGQY6sg/aJylj8VUbymwBQKpNk2HxVTldt
jrw5M3GhiBEd4uvx8h5pQJUQmpoAR9VjR0CJfs8WyfVAx+sDBZ96okoQtizhzGWgkLj7bXoXtGII
Bww6R8t+jH7C3mewh7ixCWmr03aFszviRE1gl3HGlzZTT639KpoDkFUC7g+NgW8RsOUHrNmB0tah
R951pegN5kvmwBqr+JbkQFFOpm+yFU2lIaz2wjHYkEDxKl2vZbq4J+8T09+Xuyqs0znoxm+N3GaT
8MMkK7/5qTc8Oup0DR6txB6Ywq3wTvl/ARETESVY8CO/zOpHxZ6N+7MzYDNJpoHQNu+Tvgjc2rIY
P5Erc34BqW93A8+bYiXRvWzrAopuMO3XOQH5MCcoxVuKmuOSNRiQwnqGAZSEk+8I3TSBoR7nmtsy
2ajF2gQbojVi+FbTm+7+6zZ7IHSp3i+t9vGQVc7T85lk4V/Mtm5c3uKYAOpG3oAloEavUKon4MNc
rSe0vgbWcZTtHGsNqnTl6sWJuszlVEvkgm6gacNnlRuSCJj7VT898jgkDFW4XUfyr966oqUJ5sP2
dM4gimQKEIYgEs2ARknwZjQ46h2b/wsDF+jRJbK/d4XZsCQWs1tXtZaRi/ARxY7fHUT0wg6BgNcN
NfltYptKCxc6TE+GKcYO340FzYII0N9hNBC5mosCM6IgdYVUnJYOtsbjCnJMARMUQvpe9Q6zW8+r
HDk/k8qGRuKuUK26XrsIFHWuho4ybixrmkk80VKfYee8IqdZhkiL1S4G/mbYT06ISncILkqwY7CY
ENgNC9utTgl88tkzph9BkXMcCmgKyPqnUgTnNQLDn7R+Y6a92HGu4KQYpKM+oCufq8WBpG3uoYGZ
RATrRN25ZRWK3pa5PFEhVoyRUbKnrGmM2K/irxUF2O9cGNVrTmnaofEGDzSe3unw6xrlkBT4SOzH
vk0/TliLaF+HMuSsWg0jmoz/heGdcbgQJQOgTHM8j4ONIuZk5KaQeRFLNK4equdq/6q7IPXS+2YU
0HTyFu9tn965KDTVndb6cRgOWEdC1L+wU4HfZVjLu+4IJ4Z54hJvj1kOy/YPmoZeASS0PiQCCaix
prHN/rZUCPDMfzK7xn2pOZFhwdWE3XwAvcHBpqW5OrJvvxTHK6C+zdg9lxKcavUpGKG8fjTvs+ma
uQSn63sr4CoObXE1VghpCt4EZq8OgjwtdAAEqUizQw/zP4ZPVFGurkheyYlxLuxl4k3yCCcXXwbP
YQy/b+EeL1yRpIZAEqlo/qdsFIjFGNQePmNLdB8cLXP8/KG8fA1iMnP+O/WtzU0IwLXCvk1i7MQT
eSZDUlcOfsct3bA1pUDmfVdGzwIy35i3JFKxKcJ1vAepsWFMIxp2Rgol/yN+xKWhqtlP5OzAXXYw
Tyf9GOrmnhdIz2jdJmCEOf4tdYwnnA5nhkdKPQV0tGbRs4GZ/yN5Cy7Bx6Pa7c6eu9fxiLK9NXxo
P9Gw/ogDXKm2KdJRwlcfnzh5JN5SXhGz6v2irvPmImbJop1jgh7sMea494QZGt+eKieViXrh/+vr
ysdVwUcD7kGgdg0/sHrqnUItL9nymXTGoAmuRfiKRm2uRyGJvk4j9HF/sU8BxA6nqTK6JhuD4XkJ
+r4Zs4MglWCP5WY1teCQYBXOzKDQItfMXY0qdtU7kxjtYa9ESNretWzL4dfBXKR8F4vd4C3//08P
Dx/zmz4zvwe34MNuJCuWaYGjGU/nqIqPrLyilsofMDm4DO55l5h8Ej1T2KIjbo3gRTT7i6y1A13r
Q+DBqfk4YUvzFZENzqJI9TJOzgX8727uZg4jxyE0KAwGi2j2Mxn6fVL+tewjp7rSSOUVM2iXuNfu
iKWDW1jNagqZXw9SufW2kjiV+x6+hWH3iJ5ZEWS1z+1WW4W49YRcWTpMo+Tp89GwLK6W1KT4OAoA
NR7H46NgNUip+dGTO8YgjoR5MwHfUdmSdqOc/bcyAthMcmOy+XUj7gZBYnWDL6qD0gNhxqwRzpqB
mvS8kuCGIjD3bOIfw+eG5qiYaxf/sMBz6GFdLyFuCp7C0xpa+8XE55iDy/TcMgegwbj/xW1lACZX
bqZewd1MDZKVq9oS4fYOQ15OlhW3aQJ6UWQnKMUisKtQuMOgtCW7HHSnJvDu8VOX4Q7HPmhHdXQn
eDpbfN6rSv2DtgKlYqhqeijE6qV8w1V7ZtypoM+n+PRgQtWaZJAx2hftyFSZx/9v5SNFxY78OAN3
SIbWyK3uTI0eECDAZPNH0Sna8fQ5lrSImW/DnFrizaRpUxp84OpaM9iMDV4QqYyYxLDTlFxBPdC6
mlcJHsn+nUKnDMA5dfA2sZcslyKUqUTOh0Vvd5kavWRsYMElGuVYPiRgbLGXbx3vzG20Jz+ga257
lawUdNN2QDb25yJwPc5E47dTaVGlbqpZD/8JadC7XE740BI4X9ftPWE9Jo31xuh3AFi13XCyDrkl
gWtsMm2AcFl1AsBROYdhFuORRWbFdmGEK+giAc1FnnMfFNs1zcgPkLOenITLUxBDioi0iYjHtTHg
j+ElUySaNyGvW7r5SReVViQpsGed7GmiSVbdo9WMFnGGH1JtIYJtdq4rXBTCBKnsDCHRWagn5B6R
DIPKznkCmMkqXbiFysqyxEGI/tAZKf/3PEyeCvnJhHK2LevNxnoZIFeqmdf1AGLIR9ZxIy0boE/e
3DfxPMlz+56MNTUZipT3l9neKoGlp4AS/5q9+BXvVo33W9/g7oh0tlaJ7t4Nhy674kV1I1l+fEqw
iZINuIy1L9ynrfyNsuI/R77hwaC1Nx6grUXrRK7V+S4gJJJfoJL18lM0TaACdSrTTxqIoThlFUBk
iBn/yMoj+BsbUI9LoRDvg5hiZj+mz4YuY96JXYW1um6WGiG2CAezPXvilv6ArdGK+ogQQczeC/LZ
UTgpWBGT/YVNIsWvEUyRauvCB4P/E1GdQoF+4IEVbfuXTRHu3PKgXDOoqHgs92EbDgMrdrB/SDnz
igyB6ZsrAkFKb2EV0P6fWTH5l/bvKL7zDj7tkp7C+prAz6Ysgt+HKnf7yHQGRBVOp1u2e1+2gd4c
ktaYJwy0nybHQaUH0r0tirDUvNdQ5zJgEv9540/P3t+Xlo6+0rd3uXr7GyqA55MXGUMviVJDWrUi
Goh8AR+uqOYXo2t+yQdTGMZi114f3OyGSwuOgq6hcrLQwFiSnxyQhFML6WnCggisK92rGd7QotAv
UPo1oRA9cNQroqnj5xqSRKOassPySpLcMOKd3AbvuYcFjTpTcGADuhwAP+oVmTyhCJWxSOg3qIsn
GopVhk1TG2hOB3nDAg94qJrqaQoElDmuFJZsAwYfTEJUh3ZgSyRefWZSxQz00ePh2nysF2wJwB+i
w6jYy3/jeIQeZLE/pyVv4p31Oqy6kaYSyhCsJR9WKX6PPG14aBbxjFFkqanZ2b0w8moVjR8uZ5qU
yuk3QoV4PyYHSF5TB5B6HXZ6XGINttdtgvDk6EhBWhCM4m0bHBVw+M1QvbOC6P/PfU/KYGC4C3HH
++fxxtI6beC8dLlbg7MWfJdUpMH8qLqZ5psf96KnrU+y6csPvahN5zKPVufMYUhQ6U3fl3/z8/PN
uThl0XjMrWD9X6RYvEaKZoFhTX3kA5CluRDPQCwg0lTgTwFTVW1GlaoKO7ZWNRAOcmogdo/DaEGn
mY5i3R5fq7gSnEwn9+X3Ygp7KD1OLIFFBC3M65bS/nhXCXG4m1vxyk8Dm7WZT6fXDi8HuA0GedlN
v5yjldyoOg5fU25KB6XyR47U39ANOs3bhsnFtjg7gdqR9e5dds7ZTwqq/W8Z4CkzmEqv04DArfL9
nt7k71R/qeRuA2evuAswgLXbIAR7AhOAOGe6hXjkzjrPuu5s3yOw8yL2l+a51xJQSnJpMywUhtJq
cgoBPZ9eP8BMFHMKBiKLnu4+BEH48KvMi5389dTUaFa1FM5Pqj5x/xn9XkcNPwfQ/dl1kQGYpUF7
RpDNcozXSaT3vrdTDbLweJztDLzSG8QYDlFQT2KnjU3XFfl+ai1m8+/SZKGyDVM2rYeV08CSMXeD
BS+8XLwMo9MQZunT6sfqNsBWcBHZw2cO+/pJoPAemWbhacdrJYAdu+erwJq13pfFj73484fvJIvC
j0sQAxESoX2l/h59TNF/dItx8WXl/Wo60AqFVcMuPr/IxfO1WFZGumkK7CX+GzH2GJomd5ykPYvf
TDpq1yp+JEaxw6QaX/j2LkBcmJ8yihAPxEe4lt+0ojb4czzuWwk99868+WcOTsZ8cqDCo+LDsT47
EuLbbejPWrn4y0di8GwP7aVcwKt/O3aLgKcQDoDDUXGr+xza6LbVoSQA2Zz7uytENSdenybDaOqc
LJKXZso31TJYtLfUuscUbh4kvNGFLbhA6hQT0vTPT8wYNNjSXPMa+5/OpauO/qQahcJxa3e9RHi2
cmicK7npm02WiSltlD242YDYCRxkK8cUx5iFTINgPQy/7hqz0pzjzcWsjL+ssXVvPF+AyhPInty1
PHZwREQfu37jEMuQF7WWdYfMWIb67Uy/Z9V5HMf0lDVMODpZMwLgOFR4FQ88+avAdPYlbVRWUsb1
IwqQS1nGCNaEPIEGmO+vr5Q1XxTxWqCp/rRON3LDz2GXUd9he3p6QrI1yAf/+LlvLwVHmbdmZDUz
fb+wYdc039DpKfcO1CJJgYUG4qzYnmWkoHQStmEBE+s9JY0iziXbBEC8Y1F+bVvBfrbfn3kZcRve
W6cw/TZoQpLKRK5T0l8kJB7/lq/6iLHCtrgBfrOUSom1bVrElcjy3AoOsC3s+spYXKySviMuW+6K
lT0O3NsPZS/WnvI4KrhbrsQGZifayb2SLKXLglTWw0MlAGt0cJDNFZ+b79GUU0FhCMJlvW4hhUSs
WSASz5h0AONbmPcLOJ7i5p4NUo5EhesuX6ADfFP4TgQ/UyqCxMh6x1g+ucjkQy/YdBSrMRgj3N8m
PXWm2n89HNdhUeOzIjQDpebxFGOzZPPBcUo6+QblDRFmSdDb6bPoWRrJwVBtJCs2b8FqOcyZS69v
3ETzCWrl2QQenvxxmwudZ8gBEoo0HAvFOxD976eAC8mheu0y/184vHPGPdHWS3mVpAURM6j5JgpJ
eUiMt802MgMeUMyKwhOqtKHfUa6r5yNih718kbGOXsPwPXkL7UGc7TtU8SX5EefBRdiaMvaBmSv2
ZaNylNb4HWQO1J0BlMf4J15r0prUUcZKW9cyorTOs4igD6KKm5mulDc2bXYy8GCvwADRx8w6y59Y
h+IudVqBVAmdQhVdSPvsM+f3kYiIVu099OHblu2H8MJb2T/D7d4cK62y3sDwWyXfnaNl0s51Xqgj
vBy45uxk/OxF/DNWwHSJCeRr0t+B0IAO3mtcTO/PlLY6yZqqFgR8/OiMLaQQSnbQrvQC6MYKOWuW
GUn8DItXUgJdvE5A+li0JeJFRloGnmYWmB7uMbjiLJeBSQzhTAUu4YYFzt/P1ZCA6anFb1YWe74G
0DFguaRYxWbs/NuY2mMFwd3XC1P0CDv5DzkP0lU4RwWzBqG+oRh3SM+25c3Q2JKzUes3BuDmwvlV
LDC9AEC9hnc8xXuTT5ZcJ7uI402AiqcxO09iQLBafvaBQdAfSlLumSR25orcXyAmHrWLX6u54GgB
d3MlJebmyf+HuUOupyhmNwL3+E/cIiswUHS5vpgW91KmYDOVAbUOV+0pkN2vY5SC7I5j0OSqFIuA
OPTpt0m1e9Ag4eBZltKrI4vwItaWiPvDFy0BgC6FZodgznv3B/dwGdx4Y6u6GWVVLrE0L/c3dMu/
QL5DN45aJX4A/aAyNlo1ANSCkk6dWZFHrw+NtuG/NdMVkCK62bQwnZBNWZnq6UV+7bAecWIh3VH4
MPX2GGu8qEK9QUgqqW0oxxwYTeUjeKcc6gMiIAbTD/SJb+mYtiFUgJ17w0jvZfU92aEwwHiDIJDk
CeWkOEsQYYW7XRPNcR8cARaIXa2w1bUEo5PEfYtLHzoTJSrE15oX2X7PeverzGPldh1NWvk8Hn/w
NeWPoJ38MLBdNagVfUhm7zPe52UI/ymBrwtqXZ1FiMtVZs1i6lTqm1w7COzlKD1nyyfTRZDcf9Ep
Rvn+pJiDEJD26bBc517LOGA5LleJQkwAqhuHCgWTvIIw8R79izsFZNxP4VpGXwK7YVhPQCCCbqTp
4p8e4IRoHPU9XILipc6E+zJm63qB8hEKjPGrEZ1BUEIak5bTPxEYQ9EC6lh9MfEhag76VY1/nH4r
OC/Tvoa/jXDP9QN9qLny/vKM688uYpBH2YQrZ29QF/Ut4RLisoiRXkKtjOw/Jb1CC7vojRV7bf/E
veKiaMMhXBokmT80sWK+x25DknwTHc5cpe9qKoIBcrsuzAtU31fNm5nLdNf1Ipv+URig7a9oupuB
iTXu6JGWwtftB+KywEj9AVpmcngvB5CckCYPTyRpZu3qXVZYtnlYhBuAfHL45+QsWzCr+V1Akqpz
FAdcuR0RT68ezoczZt3OEJI9CZSfkGyfWWYrJr80JA646xzesJq9JXvHZL37mzgGxAZXmp+Mtgcz
qOH6Nf60wLTyJM6euCGkPWIg8LqQVfC1ZJKsOTjHn9MHdQFTR99G6ClV07SAzPKCf4NIC4kr/r0f
gRueea92lpq9d/b31ZWzliXYa1yCjVaRtNykGc3zvCEqveQy3rZBXeU2IxP97d2FKthdmcXxv7a2
xXs5DdpbKbcs2SF41X91w0TIoishDLKpYtsXwMa9kvqpGW7eBqgc9y2sF9qdFZdxLRAbDLIGMUwW
4t6SUPojXQ+cPZHAGp4RQDqAujO3Z9UztBo1TyZDCunMwLNBFfVlu9YklqRawQwVrXJycPaeZK8M
o0MZr16fzbMCtPPfNSL56V8EaqNC8Y3PnyH7BkKso0+4BYnve7BTS7ghutB3TOT52P7d+DS5ULo7
C/kRWFoS9v/YthPkysOdFyteW6CVU/aQzSl2nbKuIGs5rxYUF9+saGyuk5ZDuNsn7d/zU0kA3z6g
/BkXlmZCZqnREre3lj1mixl+YiA8ggdSjqAFBh9GzeRGCeVSRX6g9Rqf8jVhZVwAajQu8cmUl1a7
qM2s5WfZ3nQXScBAIp/GWQmxbnXssK7t7R15rps+vlAZ+W97AjE97XJaCIxpmKpA4DMitDkPrnKo
2/SFMgq53yAzgVcgW5KGh0vQDFbKDIwdTVAa96rkiscHPEpR8gDUz6LhsEX/P5jREEQUK6thpe6J
3a5rFntnR4LY7wNU1w+RfWS90pYPq6DihyY+nl+YITr+L8W09lVjV8qELlB78jJ8olMQVyzPvbQl
YITuXByyBKmx+/O6cuDJ4rbuHs28n+DA6dDc2xjcWuKxek58LfW6UYHzE+gqxP6zeXgi+WlWjCUa
yTCtuuoDsf1lPkOIqAy/8RhO755dGFKmoE4QQ6ma7f1kP+zwbDWo70Bc2Yzm65rn4Buw08Q2QGVM
5QnALRDI0kL1tdwt7UNgC+J9lav9s6zjdqDftXPgd+u4D2xFAIkuQpLFh86jcbcEPG9nuqoanOus
Paf15pTp9N33mF/hXBBtYHAyZu7Bay9uQwzSJziupxhmbMzWllZT8tZriBDgU3t7Ee95ej0Z+cwu
RFLYHbmXwma6nhBRjeFIWsEF2uioEUGaSSR5nvIpOMnPRxn94iFQS96QacqcxKEr9d+5qFAP+qrB
+EM2gH6kE4CN7Tju7T0unCszfjvk3WocY2HqxC267MB1jAZX9F28i/o6ERLLAbZ31hYWr4oQ0Ym3
rRpsFXmg5LEP29PCQknlj2Umg2/ulm53Q9wPd3nXJ1ZGw5Nw35NdUPMwR6V1X7qBm9+e5gF43CNF
ArYdO6nnraQ/yk9igJBBwrjv9xUQLW7+DIZzr64X+9tcphaW/UhPYgjJIo5C69qELKU9Amb1EuI9
ZVR1shSth+Q5xiULuGmpGzVaekvzU23S3RtTb7/gp1RGlGXKhR9m4fWUQ8al91Kz57IEf3ubwMu3
VyHX7Jp0u0JfkLiMZD8DRmu0BiWC3TuXAFPIZutU/xiE/FbP1Ox5xbYXnbTLrjwTAGkusYGWQldm
6lB2QGbAMF7ZgKB2IFsZ7aJIpkAOwR+DQF+K7wVzVc168YWmyk4IEYCA6MMtZJgcnks4lFNG2yy9
HdLfZA6i8urgTDUVjsILpd6+ASXhhd07qPMD4Tvsl96FDejMqDSdMDtUyuL/B3nVLhYlpBDGKewk
qhVFhFcHb75UuRz605RzJjIAepcMZnFwmQgbknbFZi3U/4dTfkFdBeIc4575tkebVKu1oOtWH+Wq
xS+6Hposu8+Pp7FuY34VauucJ/iaDmHmKviu6jHAmOlOnyZM4Zd7vqs9yxZkh87BkZu3K0ZIBqh/
9VIHr09/ys1L8Dyv/gKbz2oWpdPU3pZcDZUSVi61gpgQo/lKbtZCGNOgCtNq2Zq52hxT1kjZx0An
uBebAe8RVDY3PEGF0QmLRlEMxR2/Uc98SAT+ZX5rNwlJHRBN3G84RyuqXXTE4bjOsrLEVwBmwT24
YYFKP/r8v60poSHUKee3OuMKlSy8JYtB+cmn9LBceW55bZ21BfeFRgOK4wt3VcGOEaj+2c+NuWMp
l8dhqJcSw7dlnTA5BDUBA9z63fz9vhS+fKfaP5xcJ/s5ffnMbLLctxd8BFSU95M0vK3ktD+iN4O6
9q5EB91/CnbNeNvoxnhDLLx0wTZmsodga1M4uYsmw9A63maVQbVZPCh1/K/eJYW+4V7Bcm0oTekX
rqhjiMPIKVAKmARF7JUwoPs1D4c1qCXaSySgK0T/byLqAWwr1IX/0KrDtg08p/4eaYbVvOvHkzTN
6lg0x2Lv1GEXPqrIl1+so5BQK3t6hgkoTmVIAGMgpFwhGKDfa8lzoGsPxuyYuZw4MZUniee6Kdg+
Egp6GWpLtIp5M1NVEHYm/DC43zkhaAgiTtM8pgfncVspPdXKLeEohz1qT+NZvGoFxcQbFzc7cvuO
65p+XOTio/RH1GBMExAGCgTx1TjJOCY3VEYz3zFkHwJsWssF7HDP+ABfRBstFzKm76Y9dljpABYi
di0K1OsbfOzooI0gMT0cN4F49g6FDq6xFhGNbf62Dz5Waruj0yyKq7YhlUJPXAQYBDR1HTkVHceY
jok1ZUKZzL9VPma8Pt7Bxw9lWkh21yp6SG0bMGoxzh+7BYMsKAqD6PZmd2Ry9n28amLuj0z36t+e
CrkcII8B6tBSzxNih6o+PX40ergzPMxLRYhqhuhP56blkxO58t5obo8Cp9MljIiIRBHyPbmWXjc9
Rv/idsRN97oi20JdYrWToLoh0qmNx/bO7AbB+Yp+6zUErPW1+xFU+2N6uenk6Xtz/IXfTo4jcHUk
IUebDgzZCXYjvkQmJKpYs2yr9L1Y4641v4pSZg85mmvMN6OXOP4U22BiXYth7USmJWRJ6mECzVbJ
jOAAPRufp/KTRHIgNemx8LZUg8EizEmSMRoLsFWq+TBFgEDucc5oQJGiPfpA/Teo0Ot2BUCVge4+
6R7BRY6wy/bVEKI7FHJ3lcBjIZhsV4T9QP3gOgxVUtRcjDSiievRdB+1FrkTZqFws2AnAgPT/Wx2
zLE86aRxP8zzhVdT4vtEKK+EyXfKDoJXezMv1xa8x78JN72YEgAlhfDn20qX198yAGCrezYJGOvn
HrsNG1OZwtZO+9I/UYFqAwlc+/swyRqyCd4zKyDvT0vpGd8Yu3B+iMT/UmR0qXWo+H61pxuzUaE6
YQEtzquJeRdNSqeWuJ3cbt9H6dBVIm9h312/xHwXW5DCyY1Rxb4bT/ryeDzVFIi0nJVQyxMoSi5J
RXIFXEzX2uwiUAL+nN3dHsm3qnkGLCLUFym6qrfpQvbJZLwRGd+cB7EGPRsi2ib3nv6heUXJjcIj
ftb4QjVKX2cnHT1Ge3jLBimMCoA9ZVmQr/gU6zPqAIueNU+elOpzRuIiJpTFTAQyLCF5+iF8bobn
9uWYs5c8n/YuPVrkucePnInHn70HGYnZmNi/k04lDkzNpD0U+5VpGxdedQ0cXQGB2N6gEgVfm/Bx
55OhRLrJmaVYJTgrTlDx6lmeV4wQuZf8WZINbRr0YGJHO4QjNxxOnofaXfmn/dn53SNSmweH0Nvc
ahPSj6O+KjnSKzvrW3FY12E0tgFfuy1H1crhWhdlkVoQIsJP+/2BxAxQrUIRBSdp0x9coJQTJhzU
CFlkBvaZchPAScCE1t/YFVY4Z6bwLP78Ccqs0CpKrjJXZSfX7ftHgWB/jzrQQngBr54uR2WdkK3H
aCbcDzJn/KKrRjrNGjlY6tfa7NBWvkhGAT3hY2Jm0FsW5jNkeP5JCsUOb1xNUl+Ubsf0d0ZdW2dq
n2RDMt7ciB8eU21p7ZgG1wp+Zu9xVqA6Ihsr5RWIYUukQY3C2TdXMhU7wmJLjXHYL0lkdbnHDYxl
bYg4JWHevewrLHqk+GwYsAZDGhf5zRveBSSPSJRoOlV0rMPiPVzUm0hXdPkNUjlTM98K5cYLK3sh
CRjmWqoXPyUS4UeVyAHKOhXaI4+GXPt3yj8Kj+1lJQdr8uak4Dq0i7YD8+pKDrgNwDJRaX8+aq7R
mr7r28UTWoiXxfgyb8EVcsDWVLvi52HoQkI4G25Am1LJDWrKDghJhDmUhPLpn076+vMFV9qjZl+u
Eb2xRNLNi+IdTyqbq6AV7QuwY8OaAdasyRemmlcMwQL0CF+3df0mp9nQDcQjBger2rok93vD8EX2
s7jz0otxriQ7bV+rD9DeElgmxAWFa84OrWMFnhIadg8xrrJjuzfCj+KkpxHaxhMl+6hg6y4K9L9W
To7v/FQ9VK4o0/wp9q7/M6JQUm4TsC+h9QmTSoqnhPuA0bxY3LESV50JMx8YhBKjCrfXOmdL3oqD
ScDgXDpocGYu9inyBvK5ScMd6p87T+5yNWfRILkyyHk4HMSq1s19+AXmIbUYiWlxvHBQDCciITDL
UXHlPFxO8L4Ww/oDeQ80ds4tHEs4tIW1ByfS5YPRabEdnh9jt8wMU/VifyNPklQBXw5S91hv9P4B
8IBfvR+vavBeINdYOXyZNXlB7XF4ogonsWxyr/zKyH1spYngA0GGRoL3KCOqWtZ4CkqDdXFYLck+
JbmOMmYD5JSItsSCCad3DtQAhJDUXgAw6UurT2t845cjC4kaYdx4xvCIbnFX8kiZ9oRbQ7iCLs7Z
MvwyHodNIEGUvHveanW5D9A8fWISrTh9IP+knrsozFaxlpCg01sHznxZjggNteqUNt08AhfhZSo0
bDpNeYiJJr8SlZfqU30fDWPv6m3zYGQnjsVxnYjlH+/QBMVrEgnq6HYrNrR1lUHu0oqvUdxTx3a2
1UWHAB3EISihupQztOgrP0Ri1t/RveSSIjOVWLB1VcDCX2iYd5sV/yb8gwClTR1sc4D+HbWtJ9Vk
i+rAPxFG52mgXHnwyTqpREaRPK+iMHeCsi3c2IUfIdo0gn+U7oALD9CP4wbiWg50ET7fa1hSLYi3
730OUeNMo0qBZeKLBYmYCxHujTnmXl0pbD35yD0S9Z5LRzK9rGth4kL5cQRAX2X6ACDwH+XbvMbx
BX8LrjhipScxWFkZgTtG+uiD3WNLDRnr3/sUCv53m495JeVxecPXl2NQcQB3041QAS5cJ6dLcSVl
NUQomYHTfP6/4272vrWe4qZlEV5xMjbEmjDjrkzbPP0E2BdywayX29KRXSBbJFlcKiSIwC2KrXsd
OWkIaer0jBiKbMpb/7IGpjXM6Vwxyq6Mw/7J/yMG6CN0rnOz3L8A85nMQk0kebigMtsS/4pPgi/C
p11nBraTRSQPGmuj/KqmzMtRMNz1VsUJwQyHemPgOA7nyv2x9f3WAOEeJX4U+JLmFHbN4Xrua4RP
dLM7mdQ9i6ii2APwag4i/iWJR9avLy68wjou32hQs1cA/b5Vz1HTJzaspOmxZAdROcS7Z7vTX8z3
t8BRpkLFdrU0f14wdjLBe+lmnR8a/Gytef+DkMDyV7VTRlA7blXd7bhkR2tKLQvgYkxZDDOicls4
3t7+1PEWLAbFASTBTGH3lyUbLyqL16ZpJq424rTqeWDey+xwUkiczX/TyGuihaWhr4HzX7LYZwWS
RkyAVZJUptzwru+d+Jz9Lo3rTtzwuRVfJWOlKWjLS2939YWgOj9rqkCj06Q2S7OFcW58HNy5LUdX
xbxax2ZQEsXqcoxDDv7EkM3oYLotk/dsEUiDpVnE0d6bmb3xD+85BOYxyGDoxAeDuJ/DPLVAG7XQ
yJHqsuFxom6weVAUZGF24tF2jAZesnMB1rY4IM3Yt2bHU1Gm4tcdA3nyxmnpRSofcUAf9VrEUfMm
4ioDt5pO2p0eEyMRzn/coZ5bfOF4hwRqujE+UrvsIYzYnRrVvZRbMg16hevJWuaRVXrilgtaygyC
AGZNkoDepPWVK/68OOo/mmLPQJHgkY67II4GA3QEHUyp12ur11nXZPuvG0SCRF0QSi0jEGBYvUkW
9v5ZAzZwyBdwDZ7LNu633CM7vhPXl3JT2z6pYRFbJLnF0AeFv38DVEs1khG/r1oYYBcx4Ssm1vfH
D9GyHbDsZne3wokzuAA8SOpCDD0jaBTR9NeYSuKI2jj0X4Xc+2aKXlBcPAzXiImp5I5lJQZ7b8lq
McKN7tbHIaYF3JmSgsvm//ipSNtU9ij8bzUdcXf9zhuEtvvY4/k9DjPAGujbrtC7PuJ8vp2PRsPk
UsxLSr4Enanv3ies3TJg1jCdIxZUkRpf/dhCiMdtf+q9q9QTSZDyXV3x36lkIbJzYFtxIjrSG6Op
ooxc9CPK1iAIfqXluT8FYWOnVynj3kBnHAK0aDxVFG/kT5IUZxWWYJ/BaNy9h42QP46+j45tAYyQ
8ch9p/NluOBaiokP5sJyDsUnv/gMSKpe2QaD2wodsiFKCkITJ7qQiFFxdQLWwUT0vmE5QjQZQeai
CTtv4P5AWZTsPXnoGYfdZJYrEg44xcmen8mxySEhb11Khn8+JC/bExcmIUD0hqjB2XCcWTvkkhQc
cX2uksvXc69XztLxHuHA8q6QjGP8qAWLWBZfOaS3joysaSJxDij/NxHmy2ftcCfugHTm9uYQuFfE
uAuyrroVG6Fm0w5Eg1oG6INOMxdYm+8Sshnkg2EjP0ksQ3VG9JP6QQf2+Emw/kmLgX5u4d1AbCuE
B12xi3Zv8c6EmyA41aOuTBc7fEgr3ftNrJL4KPVFvYcI8aTJuGMERHUIXLRbJgLzwi89C9uU7AVj
sHhSHIweRG45ByTuM9bdx0WbgY82AFZjsz1OGra/t7w+JvBkXZBENWpcSO5fT1k3D6qOxtOGeLk7
4fN6UV67vfyi8giQk0E1aquwrthS+A9/XDoLjN0BHi/zNST5aoODXIcyQWXOruUPE0dEFH0P4pPF
cnhsTDVoQaLx92RZvWVaaXU4QBOikQjhKyrlr8MZ27LFQw4NTXuGgl6Hc9f/1WOchfMNB26dYHJ0
ZUPIKB4vcOCd36pLFfUe8LxdM2XJXG8d2ATPUCICbCSUfVWPIDdR15zW7ajYUFJ5M2YUrEYndf/j
H/40ruZ5K70BNmRtXBrkQXBwHR0j6nOvdTUJ6MGaFhvWBwkoj/CTg4EdBngxdhjVySBSCZeVxSnZ
yJ/1T4lcU4pk8L2FNvO1D+ZNbaOf8HLGNCN+GAgbV6U0Hb0z/SKBlG8IvSKFhiRIWsDGM2TgSa/B
beRHskY4Qg23op0BxfFTwHAaNS2qG6j0j1IqV8vQ3z+IQWRV8Crb3jR/8lRpNC7y24JIsPAO/2WN
UZ98y1lJkWc0cSmyawfO2VARq+YDCDJQ3IaQm5cQJcNrYJ5i2puGKCwvWkEXBDTXY+HrjZFvM7E3
oWNvfTQTgqY0J4MLbJy8lvUq5ZVOCJxOF42uEBCYTFndpDmWHnjU0ESEdrCwpYPmLTKCRIminThz
l/5wJkHaXzAfg+cF7qz+DI0emmlo+MeOXzrYH7Rlv/pN/P9uW0BfQ1hxNynDMW/921Zymc+8tihu
DpcZhpjPWroOyMPotlRD4HwBZe0hg3fto5cRKJfGBReLL6rFMTOZyX4jDvzmacsqTeQfQiM2kUwZ
XlDJ72QMviobF8RAfGoxOXIYvK8ELY9LUTP+LTBIyv/a+3iJph1ZIHRLnGkylEdHxrJMUlWKrhIn
IULbmqXhWXBBKPQ8TdhxMH3rt2Mgm3WQrqhxEuTBT2mpiKxjaxnA0byHPf4J5/k22xFE0W6eTxxR
Y395w26IgCXvgnzGdo9aMi41fUFa5USDSHdwOhL/cM3LQ19+k2545AJrtAXZilOSxqyCPDJJgGYc
UasRH7RFmZDPbYigHCl0tBb35hCzPzMmCiC2qneofuSBIUgiUZ2PFC+DWnpb9+iYZj8yk4+PIEYQ
eqJH1KBT0XFhF75hit/QB4791Il0WI0q6hqJ+DipTXmllbP+wrRsS/dHEJiQdLISQwxqJKe72Wd1
zKMXRnBktfpBUIs+qIyvDeM+av9oQ7Uwz/Y731tvQ3OnzVqjlUL2SNL/TDaYBfSuRRKAFjmp9Q0U
rPEtRVi6bp2+rHyGLMOWHRbDLjL5wjOU1CdHpKvZ0tup88wDdJAvaRPlKuUYm5MgvOnrW3r6Hr9T
IfqhyrYjjAlpyLicUvlXaiCZDl8bm/9zT/UmlJeUowVvcqj8zaZhKCfK1llGazLWP3NuD2uvaMcy
g3iwwLCuaS0OGgevx1gNWtKRenrrblj0m9wCVS3OvMH7wB1el7vECqWnBE5MPfubA9y8vLomTE+u
sE9yxPxRHJHCeFtXlgVqM4XH0pbzWWHmON+z7RxhJ/r4240gTJqgLbekvS6mPYvAOVqMvsSJkDrG
eUgoe+Da9FFekaJAhrw7aIb9MtNEPexkTqV9Iut/GVDCJSLqbIAUPSG20A7ffmIkSPEkJz0Es1A+
oDYiy7FLPrkHYOdKUDUZbOkbfMlTOKqMvKqOdYNXng34P0MS1h2dpj1r4ZfKqLmcLiSJ4kmouxSz
pByUD0kupwL7KaBgNGxPCa2+d0/+9+E3taAQAJ0uTjNdhfFb0Brm6ZGS+YdQbZl0JHevOLfAF51r
7qUMjYFcmMCW6abtYmZWNuvjYFlFCAjNqVz8I1J+516tbzyi3nw4htG4gAftl2wNPsqbcpz6uhBd
Q21xHwW+z5FonktiTyrBueaFVZnPVlbQbDtgg1fUMlNvqDpj02p/PzraWqWviwi57hlbm8E7/tym
/+G8BEKvTRe0mszZAAPhSwhNEPxdn6HqW/0VN5rpJ/RmSNYfT1QMw0xW2Dn6gHZ19anKL0iD7s3/
yeegKYkjwG1/fnpSH9eSHbq4D2qJIkgqPutQvrY/3P+4SUS8KERvZxQezVdTqaju85t8EyujgZUK
+zHUihxfrroFchbG4DazKCFeWtHTMsPvEaTqLb9ib9+npiIo5D5iAbTtXgHNeHXa6Ip4jDQRnQtQ
3gp/gGT1dPcbfyXyhg2Al+l50/FP/Pb4oJNGNy8fhZv5c15LKzHo9BlTDvp3m+T0Ifp9kqEUemvE
rxUl1fO6dep9QBMQXJcuJU8UF35qlJ15cAVQZbmopjCwGBGZBykNKB1cVM/XUZ18CITEufmDaLxQ
obJogl+fztWFYwjtT+7SH1VOvtevksasUeTcypKQCR9EXMHZlLj9LI9TP5xEx7598khdylRl6q/F
imuXwrt3Gdu66bL8ve3Gse060L9/EBQGMR/hBb2KzSB+eUMosStIZQYoPddf1u36jKUX80iZxIm/
rQl92/2+xEWD1laWh0cNahe8ZEekt+mGWjYjLlu6R3JZ7rgsde66VIbyFL25EqpcSgzsIJw1sryc
i8+mlBzU9uZYFIxGL+klTpIv8fMcCccI2XiLn1shlMUNZXSG/vhtovy4axKhlHtPAW6J9REnqK2w
8HMCoexCg1LFVZIbN+lfmsvFdnWTf/V37ZbKGxcGHjRjVgd+XAUiS4ysMYG0KXhmKe/p3eGHzFf3
2/5gwiIlJNeFQNN6dJtkzu3dgpgrlNhTm5YZfLlImNWAc87AUJtqTQr1Uu6Hkt8ZS13lV/TsITye
WM9dUdbFnJoQHC3ChiUPYqMoqYQekezMaR0nldxIAxqRiEzJw+82QEDVyjFwxsDYF9P7sgtDuWLj
rOBY7+u7tDP1uZmHZLOKt5PckwFSBn2opC9xDG6I1IHNcLPHmtSsS87x4u2yXZicHQeGns8SQhaJ
/WOfN+Nsf+nRzifpDlVI3h9mlN0WKhgwj+84cFl3jyh8BrwCOO47O43eq5zTw8GgzfSUyc1bBlWA
44IOI1RWp3ORr1SKjGPGtwwdGPJ9V/gXNDJ9HbNXI3f+qWiRBupGbtOZ6B9pH+WCG0wKOvhzOJrf
ohzhnbZNrWIujGGuhHsnIHVLeivvRkIDgOKR0vfP3+RBGXH3L5oT5JcgzfuV/xWgtYrUCvj0YduQ
ep86ebmxXT5+lK8UWMbRkKQyKiaLyOmVVN5L2RNFcjO8Dd7t+toZYLpTXKCHUbP5FpZt3Za2sPoU
KKvUsa7/cfZdZ57J/6mX5HQ5YVoqM95e9KvUBf5f7VtiLqGiT5EpesRzdvla2nADZBCZ02uix7Sx
4GiETXC93RWpe5C3p6FtO3KRrDtdyhkINuqxLQ06fDjOl6T/YzcJdEwoSaD/C9RRXZZrm0lZ3GbJ
1IZyAWs1qLSvWjK2kc11a4cD9y71BLcTa5knNx0OeySwV+2doxZFZuB/nq6XEPwG6OjB47ZMK4zs
0ziOIYyME5Ch+EUhPUUHDLLpXuYvOEDPTgOYFPfBksrz4LatQTR8AW+WUEfIVnaBM9HN0i6Nh/FQ
+YTvIVaggV4hlSdvkLXhARsOVCMir8/s2NFN0dK1o6oHPB91KHkt4/zNHosbGkOhdfrwlFrDhs2H
QGXw7N3T2GkYjLq4ApdpbwQ/hd2w86LQbmtab0l1bD9iE3Gy6wI1C9uvL+iZPXte+/xBeSKIX4K5
iiKd5FEfC8XYAJ1NdJfiNQ7Xsoni323A82u3/XiDSQIlUlhnIMVOV+FlQf9+rJ4MoxyWPFvxoNKY
2yGxG6gbiNcg2DiviyzOyqAE+gNcYpau3SXx/X2FbP9nsa54UVNYZ8bCQwQRQOknKcLKF2kKGRbg
5PsA8vJc7LUkw3bOAIe6lT/ITwJrXNzmZjBj0qzc4OlR9Ex40DqIAG6V0PdLrYxY4balvoT8yjgy
/+veCncaoNOGrVavWyDtNMRiik5qO/INIzSmknLx/NscWI1WMbVIu5bRWrJXXiNs3X4fpLbmAITw
p4tX5+U748GLXyjEOyB8IIpLviLQRjMtfPyb4A3no00ateSss4GpqOJG06fpXjzpL6/MPIpp96UI
4/lbMlBeA9HhS6VLfHntgvh+tT4kD075Uu8Y1ojaK1W6CN/vml2rqVWK1ioCYO8bNljof0uQ4kXW
LvApFTNctUlkAL89e/Labnvs/r/3nkTjH1M6m5dcBM3DOgJnNxzu9EdTgoFZZmFHj+oYU9rtIFR3
WxsWuSKePEaQdTg3HIT7kuAcOm0tWz3xXUPUwAcpvEktjlv+BwrmVtACVgIMYYrH9/mU0jxkP2iS
+qtcznZQ5RMTUdv8dsjS+Hqx2aXx/DSuXVbmT91YUyuspts7+bqR40NyEZvwXJGrChH32tlzgO/p
RUtAEbHUBO1dxD5Xy0YStzdIhs6Oo8hRZ88E92FdblGANzs538dTBbe42xqDGFkbaus9pMWPdmIC
651hwABJPg9Tnmoupqf6poQW8Wiyp64VtSIwXLoW52Glo6ESdev7ybzoxKMmcWXCkSwTtuq5wvzH
riN7eVkTPaDvVbLO/KmUft1eTP0LyPclUOF0F3m0AFGRaM/m8ATtWwot6hX7IHtztGjyqVHMp3Fw
jWPU53EYaRltRhTKBcLWPyBFrTLSwbYtVVKzYDQEwi2kPgzMp3HZO6b2WlNk7+Voph4Ra5SMKoby
x0sayKj9XOJCmssiifYKtytThJ2ChS8oOvNUcZjmV1cyMWMeHgUhgE/X0UlHoWWL5pytfheJcwAa
i2B3sVI7IK7aRTVvIxYxogXnYYgfNI0CjH7neXBJxmontu1Umjmanf8+40p7ypRLG4SyIqStP6iS
4SKD4rjzj3JIVPali4OJvpNwAmi3oh4syhtdh+KCmo8tL4j1gkAOAZuB8ZVnhy5R61ugJegpmztL
wPFQoEwtz7z5gODqdpI8EPdefm7wOjqRJS8qjwPnzrTGLKSRK+/t4fjUaouM5r9yxoqa3UzaUy4B
2WBZrmvGRR766wRYYGeQhIjnmOgKkdwmEGiA6PZzxtYERkMK/c6JcpW9ltH7V1RIX29S/Vm1CFRM
AZUhMJPKI5X6mfgrrkmryeZOwRbqezG5Y+FHAyo14ufcD3Io6LVK4NuYZ5kDviXu0VLEkIU9r68z
oDhJA9vp19TidAC6AfoU54Y8jzKwkQeF98QG4HMQoB4SKi1Pb+VQclcQ1hOZfG+70Rk6KfYUO2/2
zdVEm+IRinFYiFBYvJU4/UnfseQbKbQCP2wS+M2hn0I+/80OZFiU9Zd6xRBKT2mlUjYywn5YgrpF
X5Y5Fau0UpMD1NAOrHi66z6FoAPUnInk/eh3LkxYfIiGVAWQ1x8+IDJVPvA3IqC3/Mi0SkaAF3nP
H7JTev2tIsTBvU7Q4yHgfMW6K8sn2X017p132iRsShE/+JI/wx6XFC51y6inJbvzvCODZMcgCPHp
rdqrCtRgNTk/xtQ8H0+IIAdke6WKu7ZjAiHkEo0KfV4vVwRb2ymvOnhksI6vcGil+I9ogxtwEb8s
3cvlB3VH6pmrj4lJDryFGSzf7tIS4UpiHBNavMwjNs2VAuk01WpyV2vcdZs+OX18pUj8i+y0Pgyy
V5pfMXaDFtqrCOl0S0GB8gcYx0inS4rAM44wYcXypFb5eL+FQRATshi8TPAdqeXZtCsZBKV/yamZ
3gsL6EFjLALBLCZUwxwrMzqi+amXyXLHUnKLmbrCEmmKfd0WeTDiLWa7R1YYGmEuTHt7qtLhe2pt
0VDi47gp7h51jC5Lq31QYN5FPoDBZqMCNw87WZv3sZK+Bct3cfxFBgvdXAdVLLeRvCoPpWZyqsHa
dDvDfJ13Xtz2UkQ+spmcljtZbUAVujONIGdyeyPCZ2QV6K1OY4uvT9C5biQ0Mj7y2O6O8UNzr6tU
d7+xthpD9da5LuX6CNMXgwfI/sPvwXJvM1bfRJqhXvC7I/BexoOuhnNHm7lIwDJCBaAQ1s1+uHJ5
t3V1YU8OCR9ERaBbfJeF+S9UQ0xKIAHA1Ab9siiO7CCo+FXQUhfOM3H+MYTKxi97kdkBAvSwzimS
V351dc2WkxNVqu7iXgCWU7jsHPMLL1yLXnFJBZOsvjkhN57Eskk535PH0EItybJlr1qpyXbefSQn
P+vHo6C8zPXRho/BTD576KqDBvX5rQ338PiSvLCIG/qhxeLyT7K8kECJ8orOYkG5IMa+pIeBO8pk
FZDhsaLB4+iNOAOP2ugaRsHQYxc7nV43zWZSIzK4Bi1J4T/L+HiEcFoGugxDjlYu0roglCHZZkzq
7spTzpjt0Zs9/KvINSJKtS+HjTgAw8Tzhq8SYABJsV4VM0o9zLaZ5AQDZQQUojotHm6vVsvqg2Zs
O+b2Pujp/anny3gNYCYIZXKjMJt5meZPA/n3QiYL822IKnZ2YPJIb6UD6AGwHgy12LQBZ2BpdOdp
Z0ok7hW9uTvMRl2nu7ZkJjpTbR2RIdgjJlOg/evpNGQHjtMfhcFGHgj25R07YJjBxXyRWaVb8lD4
FNeLhxPwgOYUIIC0qPLqvjijnFLwB4BXW7c3vJ74WBBM+gLCH2vnaEZvMVP0o9ZVYEHLcFsiGSNB
XSbH4VGwzM2oC1VSa+Epby0ZGWyMjN8m4E19S+Oi0VInNErqWoVq0vRJXEzn+rY7Dx5Gu38X3+/J
4+vfLG32/QxyZNZiNqj7KrSpTx0EaIJiSEEg/588yt5FNDlvDSlUcygnIgh9QqKvhQSsIHDaAQRW
wBeuOltiM9F1FZfWB6xqadrwtEHpIG+uA8E/JTkkbNVcb0vOT/ogrkTquXZr9QrISn0wKPU/5Agt
ChDJShx6hoj25MoEUBLLODWJgP+w1k3uJv7xl9l1Q7qgw9cmos1YkLMG7dWpmC1A5VCNuZM9yIZp
adONdQF99tF4d6WPTbma/o7Gdj5tpICybqjGu9R61inSmVGcD3+JjjCJVnkcwBewl0LR1W5g7XBy
hYr90jDZuEbHO1DeTcqeTapWSI4qpB6Y3YRK8t12qGDGYTBf6syfSvUrJQWWtBv54JgXiwVHACFb
g7sfuybteJhqsjkFpkZ8WO+oHZSU4lWFGnpM9ik0FNWKWq08xtylaO6Oi0vcADZK3BBrypWCMqlN
HZEcUQHfqG/23nMtOm08Q9U2SgmvHhQnXgjaWwwg3+BJSZ6YTV/LkFuQVmDqvRT5sMnzOIgGdgzi
qo/owRif1jdeO7XV9ztDTle4aSZAC3wJd46vqYONdJIziyvadUQBDJze4m2EDNrqEzxrV4oBjGFk
SGIG4F/46LEUk5P7nToJ3vS6/TqSLXJ2mydTCDqbp2Xc4f6fgg0VOncaCmec5jWEj0wV/lR+9eMg
OQXKmEj3P9oWbw/0E2tmhhL0EcENeuotIUVkR1uCv33RJ7++u4vbLZdeCCCDQdg+rST+s81czFg/
R4i0ujCt6EpmEkcTGHFRNqMY6dTjA5qweSS/M16zutB3UZcLZWF/JP3BRFhNn7K5he82irZFTJAg
hZN4BQ8pmMIbGmJwEQBxpdqzXeMuEpSeoR6PUUm2NHS5GyPQQOAKBz2BqYP+vBwgRAtwlnYVMNmt
3ga2d7xXnj5vx2ZzLk1mTVSWaB8kNJB7DR/y4qb92EH5BBED+a43xL8TRbqhOB63U2hsduMjZGsJ
shIuwhSeUq+B3YnpXjLovg+u+uGq2S56oSfzNqGO87R6wKPFCC1/joWWEqNVONpv74Ck5JAWaSXW
RYb4M9IQ1IFHiOv1ns2GYDuRAHcoRkIeyU/0a6I82GIHCZqXJ4lm2Ny073opwfDr6Nj1cxAiYKmz
4GEkKpPlR3p6cnBZSas3iH3Q8IsNdU7tQhU0aT2hsfyfsbTLoBTehujiadUCOFS0Y1UT48+EW4pT
odgs5HSd20Fn/SH3IJO/F4gAXB03qOo8C9NZLJLSj3zpaSBmuEKacHup1rBQLDKSjxFUPx6OO/x7
JRWoCCA4xoo0vhWogrtlmFI9eSGFkokOUaqQ6cH2ChbVfEdh724D/VZvRLLOXjF1mZZs95/SMo8c
8Tbqr5Q1YG3JBINFysqHdh2sAe7X4AMjmHcvCugT3H3ysuRC2zrp1bX/Te0pm+5khwgPfQrg+Auc
CLcpkIEcWyIND1qrQ2WHDJL3D/n4EEy9RHfF5oA4hHznbu5eIdBErS9xtt32Kk2OQ2s+HeNtusm8
6srmE7g6z3asiQbutNOTvn6gSrpIcXK6/0QSnhw91P9vxkit46SkeBmyASMwXezDJDnGOyjSC4qA
SyvECNropiebFSjBD4n/YbOgHF6YG5nm3R09pXK37GYTrBa8U8f5lKn6S1Ubs1q4a8aT8/xYPz50
44bhUiQd3/5/goWEx7M3KxzxB25TaRK6qg7oHIbwBYHBGonhWoXxuwWrWY047s6QuyEqmDpSHI+F
HyUQUFJhnWOilcKzZBLciSRp1Hpuh9eRMT7EFjxmtyaR8VgO2M8OUVr9DcJENe2jiRSe4pLypISt
+wBRroA/Ltqm7HrFbTYR4cFQV4nGtaIbHRi881SUcHH2tLROV3YqNDCpZTIe+Zu/JrqI+U91KdJB
RrSyCWCAzYo37L9NQD4tRALFZpdw4tiwbqJme53OE7LDOBVemCYmj2RIWWRuVZrkcQyaoXzGmYxf
ZqKILxxl63xRKhOQkgmRr5VXootyA1M+J0Z/4LJTQCRfCN2mxlYHnSPv8W1jrYeVAsGzVx2c+R6z
CLGAMdsdGL6+CQvLdt9H2fO586fp4JH9Xchns1vkkpL2hSZW99Qe5y3a+dDyfjXAISGIKrUarpPu
wY/m6FWMgDFR9w9wMrbJWNEyyp+I9G2WQ+vDWwJUd/rIB9Qa94zULqEmjeQhN/gGpULwITMtvOKk
W1+EI+3UeGQVY15N3ivhqv6/zGQGYXxwFXVY3QoEcq0SfcoLE4Bx8OMqtFS7tHp23fboTwFI7+GK
Dp8AHliF7WY3CNYFVJyyO/ZfJUdDk3pXGoXtNpCvjaXT7BquWyS2JslX+YfkJN6ux7AOwNgcJMON
lyFRlGlgNDrOzJMyomIRD3uPdZ3ihhQ+TTv/AMgdRoEyuoYV0Am/cCgtEKGaYXYhtZ3PJAmV8glp
KlWQ43a+6vxK1OoXhZJ37+UVHHXAo8tSflOvd69LDaco8nhRBeeLI4yRyDsQyboaOsI4fz0kA73X
+Xk9jhB6GIDJYZE37QPOZAsdXrN9b91rO+wg6rJxZqitwxuKRDSox8tw5BaUJpSQ8LYqf0peQ9Kq
/Hv0YyaUTjvmo4aC0Alzn3US5mdSkjk9ky74kQIusmf7IfCuUqfSsdEj00ggCuMupxtiNxmXTKcf
gGF7dbiDNKKv1xqvz8psf1pg/ICSt6E5y85dttfxhkB4ZYHl2qHo282Z0qZEIFMsRfV9rhEVZzEL
gid+JpiKfJPY259fbAS8tL8aA8HcwncGyagJRqNs27EZFwyjan1dkW52ijfEXJf51TZXWN+oKHMD
FzS2wykyXL9GiQ3Da6psabWZ5kUhne4Y+reV2r246DCAoX+M/yOvl/8m/3Tn6jiIBQ26Rau/bdhI
zSiI/pCuCdyUcW2AP9iErlt5ExqWoONeAbBMrvYmAAFfg78kAdHzlANukBDAB+txmI6lFiBnqTWN
WqxwXliXK9Qtau4QBmqCDlE1YFTqH1a7VjLcYzJ+TktkR4OBww1rFZj6zDL+l63gLk/mCE7HetMZ
kfBNUNi+oHz/0cpYxu5GVo5Omp+Cv9juvUyYwNkMwjEBGsLt+3wfNS0xI243tsHb+05f77NpKP0H
0iHUWdsPhSdsqidmL+bRHuNkNkTKSUOybrL9EjdP7CjyUNnsPSO2vhcfgC6IPge4Ww5aC6LjJB+O
Am91Pv6yyC+LNrfSQP700YM797waXYGQ3Kt0k/2v4Uz5LI6S8KFh72j7/ZqZymSAlOK1RzJWKVYB
X6jU3axKMlliFxuWUJTq7nGJhu6A4sZa0p06oErnSCxsSJ9AXKIbw/nPd/pjcBdTNA5moyxqCtp5
+0pXl5JDuKZdhiGoBtAcXt1m+sE4z6DAWJ6BbR6Fo2mUyN9NmxcVTcELGLgsD4yNX98uy4BcpyCm
4iUN1c1BzbEagVIrz3ahO1rckxuWjnTGkDqvYYbX0nG4mGoL0B8H/0yDMfjs7Yr51KTdFlhY0Pwz
siAZYNqK4tv6hUX33eQOjHCfmoYuOpSWN0myDNf8BQbNpsb2O5RK68lKYaKKUU8dnqZSX0aA0veJ
/u0yE99mFeK8E5Sg6ICvhJ7kaPr4htFASP3AJxYv8c4rDUyH3O2DR6IMC8MtI9tNB4uH/RqHlv+u
qS0eSV2k1LIfzylXnWToNOlCTuV81SOcKBruYCZBw1MKeVEGGXE4PetkOv8npdDmz0xQbmXxcEhb
X6nBVgkNV4V26WLRIyiA0XAB4T8t31n6MzvlSApy4u3w8jz4kZQo2PsVTgM8u6HmanV58sTLWHUq
ibN6cOF6jTCLKiF1/QjapZkeUmLySp9l2tL+usNgtuFr7y9yIVZx0JMYGOVG/LUDscdbXIMY4dES
xSqH6lpSCKDzKJmC6x56/kGbuZVhXEMxXGvMxLNS1SNgPGD99xQZ9vj4+Cl2aUkv/ZXThMTeX6wL
LALQZ7LRT0bsgPDWnPSu44qGEaQep+tEaFJVfyX1PR00yqADXRrZbGUcR08g8M9EbiI6qNXDwPzu
ORC21EIykpzIanFJSwB2l3GI7h550v68xMKzvw1b2wwuj/uSAARivyidn2LP0BQmruruWVijN0ur
iyhHa/z3GIJbH6urqYagLp14ZF0v+Zxhol9SFRTndur9R4fk788LAiAVY2hft+VHMIIFAnfWq0XX
4UZLgu9942cdlPzWZzvz9YO4/TMwQBmwpKRjGU0E6w2OjHKCFaDqDVosr6oIaSvn5NT1mswy6d+x
KrVaQcq3/XzKAaRhNABloAyQsiZqEbz8kkp6PC3QB7lCTwk9kBkZCBJryUnY5oqR2YZPkEFsVfpP
HIGf2myPcbfKHmRCViDFVCI0fuoHD27Qm11skqCzpKMY1BGoXNmrKSrIzHu+Z/ohq6leAzsJkh+E
3TlwyuTHl8K1fvZOchfvV84QxmdCriYepJh7AyctN+HcULPFMn44TVKKZCEx9QtDj+H9PSXs1N8B
MB1ts0fL6Q0ZNJiShlYgnsJsjtNoHyvpP2+kvNbVEfKTBBHMW72mPij/uxnPoirebaizEyvaM5gg
cay/SAej4iUANRHhOrIjJfHFxibmgMzovMvu4SsjIfyyvirs1tbdyepEFHdCr4jhtbxhXX+4j0l/
ayryrF4SuANnFv8XFvKMq3DNTLo8gui/rhhmcpIkDpE0GGI1OBZxw2Rxxqxv23QKV93g4bvZKSUB
/52R8iwscHT3QrHQtWcdus9AM/tZZW/B/JVMpbtrsalrdFzwaQgAivUN2Q/wGQhMdvnPMfy66zlS
K86T6b6044O9Z3AK9Pws3EW8GwH34OUojYGbgWknp0cQwz3t0VB1r3cxKOyEBOSzI+oSrNEsY34G
PjPnh3I0nXDUZ4qD9dLocMMcNXoGUGvuQbpO5XsqWWp/TXTuWQ/GzWuXQgMU9xhc9wwCn7wkigtd
eiPHQ5M8N9J0MntT4T1XBw4aLsp0ffS61u31IHQeVnFG8xcXMUkAdfDpqkirEbboruVs2snKyLZd
5JdAw93uHHkftUqeJAPF7c9jDVJUwsoZ4nOz2lEmNnCktHnSSOmhhfVNkaghTNwsULulz8FXiUwi
0WZUBB8WmRPc0tH+YAaRatQehFpXu+o/1VseoSxnQ0aIzHxl3htyx6K7t1OkSnEdhAp/Bo5o1OD/
SQI/LiaDrhnnJpoi6NGtG1NSgCXRXjNrpacmLvdF5h3JcCIyHT8tgMHH2Bw7sUE5BV23Spc4UOrO
hUMOsEbOPP1yWF6lr1hTCCjW5ocavs10sWaQeggy0K334Kc9Urt5xTsBAoRMMN839UnFFQGyzEH4
bJZaPtzClNBTeD+Osw2MkzvRgA7RnHhbX+jPsRj8RpSwERKJxzzdCzvzmlhCuYsktqjJwyhrTgpo
MAob607p1WwiKZ8dQNwhvsW2ov+CWFdfvWltWbdiM6IKXzIvHXdMGeRZ3NXgAyXnlm6UKwSsUz5K
m4R0u/bF5UrDdqNcAoAd1XSKU30IZPhxTqWBrp4BmFXffT89tCQ7Yl0Yn41c1y326ikc9m0Ycwox
Auawqf1IjZyUuO2yPrpCQpmfa9y/tC2+HCoIYB3mBVg6J7HkDyqkwpUcG0LKVutl15FTVCXvKMoF
N5Z4AaVntOD7nKtFgfhWOEWQ0BP/XsF1W07wuUcwheZPoBXtCDcIY72X5ZlmiwS5f/ceW4XK1GTm
KKQikUEB8PEqL4anito7428fIsAtimGG4mtIDtHkOWpEFLmtO76C4uoqBDpdX1PHbwibPaQrn8C9
aqVcwbCeHDiFsSCQ4lm774BnoVQvWUA352LUag9FJmIDgMWcH4SED8XS+qRAVbOb0g9ZFCJwNICM
ieILs9zrcKy6X6h/bPJ0LxewZKi79Pf3Q5v549WDhsMiEpDD2x9w56K7HYZKcdaWnY2Io6mxafYP
ULk6m24UVSx5M1QOK5DKrg2w3AZKdz2toNTFC2ACfnCFPtUwrBXADLN08rbzp77UFaVZu2dTzHEf
A7cKtu2uU74jNoXNmWaf8so4SSAIyjAGnlwwpWTSPvrxH7/KqsccS07zWlYP2QnGis8dkGY46g1L
oPDP0N5pJnVh615hA64T3Gn2OzjxrEQOcrYkDTSCTT6FxdkMB/mnoBCAo29j6cIgwL37L5i9PHoE
FOI2WuU9KCYQdp5WTb9GcupGLEmVVDeIE75iTtRdnwy7fCAsqwp5TyOuFtPdo70ZxRlLYAjo9ctn
1ab4wzdURE7dbpW72g5RYqmXFNTq3AtdDXBvaZXJdcwhqU3uerkzzWxvKqJ2O7z3uM6YtDUHexid
Zs/tqZn7w7gIv7UOu+TkzMMqPjiDTNAcJMkJmEc2czq68oZTKpDi+vHaiP1s/LDoROTgGhtSVoqw
sMCFPMmAI+6uAM+feR+5HQSamO4gyt2UW8Seu39hXQe5wC2byopcT54unkaICu8SX1EDF6pXLGcK
VH18xTvGMiBWnKcmzEqel8ARyQKqKmbF1PGdlCQ4GCZxUESFa4t9h8U+vcQd7s5k5V1LRBBaPzY5
o3y4+W+OBfopSxGx00P7l+CugpdPFUUosyg8UG3qYrM3adkqtMCcE0jQXYhAkTxTxnHuBxjfZU9o
k6h3cabqhkknQEAVtJ/qj4LVZbPezD8FL6lPtFGcYFVWCozrP2iBq7TWDaPju2JhrFVEk4F6tlC/
6MmoZC8t2xtyRwouunHiJGf6rf2QkpQA56xch/PU5hFRR1HCul16CyUE+cNx6MsZXTzZ/RkbxHQ0
JaSPQi1YqCzPq7dh/namOOZDGhQyR0G9UEDsipNqHn+BChoZi5dOJuZ+92hSCqahiB9lA7JWpO9m
l7UuXKAnxQiXuozzbQmdOSQ2BZd8pGL8FdskDzPnjhkxn0/HHzWtuf8KDqMc0F62k8ezidESfJD8
VR1NWXfDVyInNyKOewdyp+3jkMibGcA419SAfiq2mo91MsATCf/yCNCk2kwW/sMrnoUxLL0i+UyS
8uGl3mftgKbBaEIM99q9SVU1Bs1RJowgaI4psrcypSdGVMHWfC8lFMCc1Fnrdm9eV+ExsJRElCxr
tio76MfPIDdgbfZLvBmHzOxTTwFYNeqDSJ4uN0wHiTG50NShfHFGLT605vGuJ3iU+drmzU0IUvmm
9qISMcxrKgRjgKuPjyIxwx7DmdaPwoAVzAN6GNY/RDWmcFXk0JJromAOTYdw0Vwlb+KM32EZOwKp
Q5DofqVllsj6C5w+rK2kUG3q6MbeL6LijXUSwYc1tRg4CStUH/X35siAQYr5NQ7vSuZ6rmfw0ROe
yEyEKVngR4tgOxJkqL2CAbqt7xArvJKWWntCI0pimsxHaGgxKR/MGFj56P/Hcs0j6utJkh9l5z5o
0zvtXTzetQ+ng4/Wx6BuUYFb8GclTrW935Ry9TSrJnflMFARgJMGzGDiGIzct1yPADF0RHjc7vil
BEQBi+hkwjdH6/o6spaB1ewnVrtH3QiBZxKznhO28r0AxlBR90YOinNnCePhuwLFB5UYx3m68Hwz
hNny0zQyL6Vj3L08d9ePTOvdduyFKpVZcfvJaqqPgQh2cNM2wWxRxJByPbuNL7QOh8waHzC2t9mg
18psngRw5Z8mVV/ZyJrIqmO4U0DKvZnF0RyiumxugW95fTs+EkW0ov270eIKLmyeCN6f0/+QEq1I
enXNDLgmC9whbBlNLbQ2PUsVD/Dm2mgj1k6i/0HNdPuUQMFSBiLSXXQDca6VuiV83UkUej10t0dD
FVOFvNvuOuR3YVYUGA17HUaOiA+OkShc5r44Uv8JN2J+I+k3n7khJSX5HtyMEiPNxFA8C/PCducy
cNBo6v1PS1NkuWsxAlOwwdbw1SOk0U68zKOV89Mw3XyrpeA0c8VbduYxm9fR3SmQqgC87d6YYCgY
q6QTnpkVooe1Ka2k1QryS2/PPJBb9B6ag2brQdglAFQb5sjQ8UAz4GK7DgVtmKKMD6YX0yyq+LdW
PoGXre44eb+jUf5AMylgSQPvyAZ23a02vQ8n8eD/ThxwGVQfll8hMau8jwGLWPqUvYQHG+01RycN
otciIljkfj+CNhwQpsaAVOEZyVISXAVIczww6Ra6tgQjGydkwjhR/Q4vaW1TqTySmT6N3ub3nI/Q
S0d0g65XG9pgI2SJt0trEo1NyXlMqm609EMXHlr8AHiniWCj9UlOTiveyCM4GuWzEr5XQ+xCibKh
goZRDoCy3k4uiQ2gsSNGkMZQbDLxnfPIrlGEGvhze7Z/yne/34H5tLIleUShi1H6sOTtK4ioZsaO
xYtbLFwzYO5t5dQ/6ov1gW0Bg+NXSX1MKKoqIxOmgtO2aore7HBsfdkEYOG3nW3nnu84yJDiIJfh
tdcvoKtz0YfDU+RGQO1QR3BIcLxeOvpzSVGtjKLx1YvNoj5mmFC15yDQkX5ufAc1bWaqnCzbFUHn
IHSzmg/R5+guIdvjb11vR0SIf9Yb+IUOn4hh8NIKWTVoVCioC0DNA9ckxkkuMpEWA5b06ex4pUWE
HC0mOFRb/SUrZMheZ1ERoeUXt1/UjwHx/r9eddYQttbnYZAEgWtdjmwN17wLEDwutiM/nCe3hyZw
Xk4+qYs20s2QCBcm2IfHWnCogo9TU4wCyGDujk4aYgzZP4HBQhq9q97g26H6422DBPxvQOIm/WWq
D8AMgKVcLAkfoLZQ65s7EN+Wydnf+4bAHmjT944BHscJVRjr5+kX/4gbA9o2mEvA/7I3m18iBl9E
7twIlw1D7iwcYYPtXOjQCl2OWPOCwo46rcwjMB1VwP/itEDolXOgKzR6Fkk9cuSgfgAa8ryKMqmS
oiBVHB4vSDYU5GsXAqve3lM2suNTxlto68aovy5qpViwMpMja/CGK8pgFt8ol+Vd3V8igV8tLjvB
aQfzXbjPKy5h8Z7iYMHXG7qjWc8nNNQs5d+tWSByoTh31u8z6L6PPmJ90rVoWaO1/vRuF7ozqEX8
czdqvjKqKvUs831i5QSZiwSd1qvC27QOcMB9gh2Z/0u9VKE9hh9xV2C28FoGdRUwmPaX/tHzw7ct
z8G+OYpdtPdy2Ie+G0OKw9S5+QH+89oMluyJ+Zq1UGds30lsD5sB2nMHgj+MCEKfVj4LGQmZPrJG
JpVPJU6FZFzCcIXig7dPyCEyVhV1a1k0sNpta5BuNM57o5Epkfkj4Mcv29ykqL6yiNCI0hfcl1QJ
IbcWPngvq7xjB5XgdUqnsU+5dPzFeoNb0nUFA1t/BX+KCMK3Oeim4ltvwgzzjMYlFxlj+QSlqusM
Ffb4JFoGFZqSrrvFFDYzDgAD9RvdnGAhkRsyzLzHR2aw/Yh0IeT3kRIAtM4o6fPvX3qCW8GxcK0P
furoJcfDZyY4mWGRDk67Iovi7F2stTvWrNey6SIoH0knCH374lLo3pKL3orIEk/oMZObdes/Oqd7
2uiayfEGAglkZRODyfuns/1ZwhTx2FtCSmvuCDLP74KskJV/V/lUY/HTNfZgfdcZvYdRLsSAN0oG
A3gWtZk/tESMm/oWGGjn4dgFeYPyVHomiSNparBEE5dPyJsmMuAb8XhT04ggbKEHPZwTfb72QS9B
nWEXb4+woQEgS22yQLoFuySzLmSaeQuTripooHBG8fbwMrbn5jDQu2iepd4M1czO8KIC5Z5X+Igi
yrxuL3rvPeQKSMBYCGOEtEnqqW1YXHG6RU2sv2sOBUOq+jdJCUdILViQ+SWcZWnWIwb2Jk9vbPSt
MnDHpQu6WDRf28DHyFQaWSmqye7StPyjhgqSZALKyoZb1gpJmmtC91zmWaVSqJNWrcKgjqzLlpoZ
JgSKPmuLfMIhKpoomcAYuwEDJtIGx16geL+/0Ymkjk8TaxOVMGDc9yjrTNDRKMw4p0YLOzsZELcJ
plh82UDQ8gvKVqOTHz1diOhY3Mne3Z7YAL138tvqgTMgE1kVwMJkx5OcMERSJakgQo79Myf0STww
ZLdDpHI8kSYigxjhlHRgUa3JTCfLyLVm8MfkOWvxDQQkQqm39eQzor2mNR0IMCN0Dq0rdMEFIxrx
ThWuOVLjdRlysjxyJfJJ9Tbm9MzCaciCDNPGRiLIc08isygmcy5sVwNLPPgMsjHvxB0ze+UEuZuD
Nj/CP1QzuauecZJZk2UNsoOsGTbb+ZWak8Jwyr4oSezpgZ2CTVpZmwSBQTDtiDxqsQEsTDtbAJcx
UqL9izSmhdL3zsoexvnmzW/egVI4B+SEBmLIf9fUUXeCmPbmxENv0KRwyiAToUKjPdEe8w7kJGi1
B05mOtOoBW7TcVTM7GyGNINjwHbi+v5h6VA7huRCrqLnlPVu/JFCyuh3b+MIx2m3eTFlIsUd++sr
cqu0c7F89BP+mosYzkFNx+hcYktrJQiwpqkGWmFMwWG2dVCc3eClgRJYPIMQM+wrryvnvtcA95M2
X3bItPKwKhh/ZZc6V5+AcrGzllN5htXvLr49wImmu8iT51mmZ9TZiVtTu3aWfZHE+lLJPl863xEa
uXew1wxYHjTVVGg5XYj5HPHbwlFJcgFjPFRSt1BGNO01tvxHkvrYoDA9Sa03jMwptJTRodqezbyp
PRF3kDoFkTozAh6D8iqNv8sCC0gNZkrf7+eXyAXyH0e+DMLV5NoxSd3ARnamWFSZDswCAYOLqTlO
pVsyyyGkLQkK0mLk65oNuQ/fdlzFDzI+ZPRxmHwcs5Dqm4sq/wDr65kn1k5g87tzVDeM2trigTOz
cDlaqVbz7V8HBsVaSuPRXDJK/5lv8Cov72K9uhNrtuFUi330aqksBirurvLT35ZELZosAC+p+obv
3P/PPgXoFMBcyOHwEPnHofB5XTXYfyt+Gf+mSy4oCbWMO28TKjkz+ZJZfkqvoyr9NzEVJ6lwYxY0
X2mqfK3WmtlLQLjpeL3chi0i1yrnlpwANo3SSjUUojEbjPBzyy32cqXJmxaBhdzZ1DRThcZW11rp
DuTpQa/Aet0EyFkocy3vbaJRaUKLHgWS08JyROGHGNqIhdWawhuZwvR3ky5ToMhePuMzXAHrBirK
XXsxyqEntze1jfIKfRDiz3zPpNGySKbipv/nr3VEEtFXEE6Pe5LsQMUaby8yrR1gcy3lRL/y2aLF
fbOt3Sdtp5j9SNmm1zqwejct+NWq7IkTBD7qCOnKQGFbYQWhAH8MlMWJRISF1kyTL5UtP4DfEUzR
lghVmWnLs7WYPJDK8VssPeo2go9sn8FNMUd+UAMPXOML96pE7cFRjVuHeYAgUlr1pOTRXzseRr9y
g05298CzI3xOAWgcavEDl79hjHra3G48dMN3c60PE/21PWCPNea4SEOS8Y3NnwlLDSAXRL/67vPH
cBKullYtQXnDMB4xdMEXmh8Xzv8oC3PhF9p7VcaWmFYY5S8UbFEaVesH6NHk3r0skcZPO4zntG7T
Y0iG5KhinjBD3qxABcB9Ww48Eir4ZfJ7BuilwZnbjdeSk/mSDWNgoD+BY+I9BzIyuMY235hDQYCJ
Rpe4bh/y3aBF/yLLwUMnSPdUqlcX80Qu9254yDRpICb3Jpqo+Kejq1PYTQAwSMDTViIVH2S8f3nM
+04w+nXio3WfSsKSJLw905hj+QpA7W846oVahqKXWW+zW2vnPv3V7L+4gFi4VoKVhFfG7p3XetXi
JA/Oy7toN63bIfuf7qWEVsScpEsF6Ic76UlqXo2NyUwRcAabicaxu/rHdOMSK6aAPizt+iHfedy+
OVBcg5TGctgfClXCVIWq4qETRWj11EIRx4eUUz+FCAucYEaii/HwsjhpZfnaNBZfJWqE/ThGSaua
EpxkOtLXrKftxXy0cIhJcR3Rd8fKmIeJ/4+kbk8GzvhUg6JtvMjnSz+a87MFls4AwIfKzHdZpRLl
lmlmPBD4cUp5tGC6fRZH5O6HrABdnvAdVcVzUdmwYfih6Xyudn2yiZfJSsnxQ99AduwXflVUyRyt
1tEX/vzMshy/VEohP7jEVm5esIv2DfI+aa6UN+6ZCxqanH8HfoULA8Jkk3uNOB+gW8iM7t4lhG7W
EGrem79CMtoM2BCXmx6VLDdmpkeszlEnENBIAeSBqxfjYQ++taLl7m1Mjt0MobwYmrJIWaaKbens
ucojcjy3029qWWDiYbH0CfMtD7NgUZZLbPL8UyJPaUNhE1v6WqsSND4PN5PAKkV9sGw8tWe0q9Gh
RtGhSfNj5N+0zTyCGOXz1xCtm7KvMzJDBq1COtVsJt2Z1pH/18viifjTy3iTKb5URfNIpv1HLcGT
shy4JMYvY7n5ZniMexiO35MT/p5LhJJCAybZblvI9FLngiH19R5rAUjNUOcvvfI4ZngUCvLMQrCL
aKps5kO9Xu0rdBjmmZMjYAkDM9rq0+4nRTRIzxGwGs5Pyc0zCqlh1KMa09gxtZLJv3drcOSalvOY
u+gwl49mYmKd+4/xdR3rgODy51ahBXI6SkdQTrAiKuhnNppZlPOs4AOI4YF5cTI9qoiYVQx/o7I0
DVUyRb+AiU1MngsISswj8/nIvTpx6RswTtc2m7+6a4axPRafYrDtf1Yt9tR5uDFmbuTvqeKRJOO8
BmQenrdwZtEMpAvGHZ57tAm2HapYILwnZo+skShuU2RXP8LC2qtfJN2tGaGar2O5loJiERcH8nvi
PnwD57A2zlfzcdqB0LjyBXhpQIQZnR2oNzeDG4fx5CWJwb5nfA2baGrx0ggcotiRb9CjqQIxtvEX
7rmh8S9G7wl+4RJ9UPGBP+GXNwWQ+kR8Ra3Hgm7iHkAmL9WZ+8gSyLWHNWj1uUJ4WyXsE5w6SRsh
iyo8kEWkW01h4rDPh8arFVvdib+8+141I3JBqJDOQVXaeh2s2qiKc9eOvbEGCviAtEqqJfS8nCps
fxiqYhZD8slrAAzwPj9CaWueVy/coKrjLiNvVUzn9KYiMvR0Clx6PdrV3TjYYSnbShRKJvfjjkhF
tzSNPGrT4kIitE70uOiN87VRKLLlH0l4JFFXXKhewEUFzRqcTlhSqDjcFsZNsOaUnqr4pyxLidUm
bLeRdq9GbdyX7El5FilLAbiPtAUDJ1Jka+xUd2AVVUh66tEe5a/3+pEFNfWm+Sl2xa7dcPo5jT4o
/4ycp4HrkNV/mkkOfY6vSs3Bj2Tm0KkUdg1F3SCDKBJ7mBL8cRZWks3JKZDTmtG78SziWDC8DjSp
drnlQFc4OegDTvz0M387gR8AyrxapHCe9S/g/NZex7w/TyfdcjcmQViP8q3QPjINGJrAu0uUXDwX
ISqPF83vDDYaCclGcGauHF36LsG/ki2QCZzNVZ2gXlZRJazYkNRwSJwvnWyoixcOpmzQpHNKL+P6
Pe72xiT03H+R4VJ+aN9WeSotO44VjLAkFEKFlFXaqgfUL5p10kiMQrYXkYPD6qZmykOs/BBOmIdy
UpuWKu3WWdzvqin8cUkgzpCz9oNnQwG0n4UnNtsdD1zNCGsJCR0CHL4idtQIE4EJhHEg2Pd9Bg55
akclYAuF4aeiROqNmdg3ToxpRU6/MBamqb2/xdkmgHaJLXZ6kK2TXHtpaa/C4VdlXVdNsCTgKm9j
GtGg3UldN9uS6CJPQ6N6rzjd1hNJ+bWEqBzwSI+SDDfetThftpZ+2QaxGNAG2EQJoy+559ndh2Pt
zvaeo7wbAXzV0UJ9OtbZWRyEr7XJs7Nnsi3JyB68NRLydmNlb0qrRBiu7YvbTsTP6GaKwrdgeEiA
TwgdrUeSU6DaGQhijU/JD7lBIfTznVgrXsUIsE8xeot9up0ES0xccCd714aJkwxfheMXOjoL38FM
KVVpDReL30YeQAIoxaHIrLaQEmSC2MQYpywK8/fZx40xXKgY4Qdtx0JmxOLWs529kqy+BpvpTrlI
9ZlEkYhVLCrG+DT+VZanxszpXKs7fWalbD/N04O1cReJRYjdd8CrukFdwZREPFdZwH4kh52EG/6X
bpoFVOjOasrAjybjISAkqteUNUWvl4nkQ47mZHoVF1xLhdDsd5d8k49ss3QmT3vFjnljb0cQWn2a
UDq20swsuZqokRwtHpF5vCqY7NlYtZeLIbacc6nwmAn75p92K3lGcqFBLoh3FJsd4NhpcIlaEaGY
y6IWCJatABUeAg6ioyA8RuAsAdYiv4nEizBFkO/Xq1afkJApAyPAjbZfpUNrGRHKAXvg169GnMRw
MQbVcUnurS3HRXnyo7r5M2LL9FxzVtg48Q5qb7HsF2/JuAh6wkHb6+xNmD9KMRJI3v5in2UABmjk
KuYygt14zRgthjxuUmVHRcACXUO5CYliUv0M8dLJ7oS06OYeoZjm39Y/DK3WB1NGRnqjTE6XOFWx
Cf29WnWv+V7/hzXSqfmb/VV5W5PLtDS83at4gr4/wHC/PcgHmPBD2IDeMaxJfY8eiQVCuekEAwEo
rys0E6vUWlv7JMW+nOEVCjtAbXGquqDrEgIDVAmkEOAvnVgQLiVejuNbdkOSG0z3KQJB2IvVVTZ7
UXxg7devcGGrYnJqH7I4QSIKFuyUtFP8M7hHMB4/tyaC3XpqVF3iSd/kW5qYUvyMTBNCBwadLKao
hw6Jlo0xylsPB+pwqxNDRu1bnHmo9HGEeSYbYS+elFGpNbw+ozHpjAnZ6f0wNpKl/RDPrMXfgm+n
FPIUSADbXWqRFk8yqY20RFJOwhSCRpUILNsBZ++eKYiVkvMZboVC3sPE1tHxpAjpTDhLVydabmUs
3fWm+MNlIKtU2LHXtY3eMLdYJ4nzdkzPnzHF37IJGjuGIMV4HB6nkrriPB4R2YVOsTsjTpWrWVC0
q+rmfh2ikmK13fNJFY6uewI+EkSrRBKvTtj6Ty9gAiJF5Jn/BUwfNq8HQp2Ng59aYTtt0oyIO8fC
dIOhSsYFlPHR0e0sAz3CPfS4muc3nQ6Csui3PDZZXcrOKbS+saM4o25XJybq0X9wUI0tZMYIy5lS
tTrA5BbfvMBzkSqfIPnn14wam5G3WzbWK4DM1oJO59ihY5yV+QAD+lfCp7RpDO/uEiTEWNKrrldP
R7GT6OflkcrMk9mRUg9RQL8p2O36XfjeBBlSIbkLxKQ6PHdTj19/nr29DaqCNEhhrGC0LbyPCTGW
Bz8ThIxPO4aEeVuNw5xDpDe3o9/im/NugOfaKSM1ghC3GjbM/7HqMBmYYCknJA2xx9hVwln/jEsX
U9R8xz4vGurjwOOjLEPCvPKUWlMvR6WtV3seu4pNfMusl6kDmJ9sG+HkJvSa4jiSWNhG1Uq4Ovlc
ge0+9Ngn1X3Q0jICjgzFxg26vwkTC1oZPEa1ZN85+91yszz4gPiOiMYkZiUmISTYAyL9SFLJnxue
dDIwldB1ke1pByGThtOE85okNdXkaWYSqoNjYZdIXRQS/yqI5KKv/A4hSh1ac9zuoJTpIuziV3z3
6RouBBlN5CcE9/McQ4XGUkIT8SDT8gRGCS3rTle7Sm7fc6TZWsHyyOQDwFCff2o6tHvxI29Stq5+
AeO+Xm0JlnwxnnxkoT3vW8NQJkIXmNJY/iPxGZITVrTjTdDVa28KZ1L3fCfbNFOB1pWHlJTDth/+
eGNwWySHtdzYEtWP2vBjHI4hTpFRkb/RCDyKZUjyCWI6U7itJYnEIME6wnyisAp94cEp0NC18yzK
6tVIfc655hc9ItQyt8Kw8rqFEwM8W5VED9zeoNFe+snky5k/OkViOK8L5pcOBYRrJi9Zlp+ShuoV
on4QCXuWKTADA1FkTJRnLrvx04fh2lG7sT3QRludUSgtTKd381SvfJeI5qiI1x7fa1MeZBoFdehj
JAvMaZydztZELO2NXslYSJXF/o3ZaXvRVF2MBRTdgTt2eH28TtM86B6+VX0kTPD9llNNohTlwzZk
+hg7oHARP7fLVSu1zPtJCpLFl5YYVXAEEm+FDlpXS+ksEqOuwY9BOWi78oYDW3v9dgDfhPxhRDqX
nXA2jCNlHgktPD7rsxjqSVq+K2qe7IJNuVo7ePI0przZ6YHZcby5PiXs7ty9AIa4U8ZyBm6AiLyy
MDf88Q13CUTI1hWRRSJPtqFPJBGDp+cpgIsfpXfC0wVR6gQeBp5tWIcdULQ5NzR0fLvADKwCg9DS
gMByaxddGQSIb4p79ZJ5tgEsAg/59sLR1cAV3F1A+pN/vs2GMygLmr1Sk8+TXTtdSj9Jxfukt3hY
wHealDX8r189Lq+TNuBhpVt6LWIvc1naG/3zaJWID8GQ089C44NkVWxUKdAydmbpRvZDrYJz9/3H
+lQPpZDa+yzeY4758Rja5HbZEEB93EWIBZHBSfQBrvvuCJKsOvQJ24ZWSAJBHOxcqj7oqQBR+VBR
g+CY5nYmQfCJk/YhwVhzNIpLYqbMNvutZ1lOD5dcomvVZ6uSV4cojKfiws3JcUylxiTRHDbeY2Uu
Y9TFcOOFRRx3THBem5J/ofnEBwiR1P7rzksqAOeN+EFNpZ8iRmvy4PtDuZIRK5Q3PbRAjUpQbEJE
Zj12+eM41WGO7ylmD3dFXx6Lr5iKLn85/ONJ415Gdv8kQEyDMfg+vJAZrSPgRMft6G7AqsrCe17q
N0CKgwRdRU2UsrObisjbJPoAPtPYVdR3I0SQnsMXN6bo+ywQu8VQMLexDiAGz0AaH9gpZyRAHylL
C/Bv73QAOmzjH0Jhbcnq18qRGEBG0PO1KmMggurQuqNBHHGVnLK0hFzc0z9R6bMu6S6Y3HnWpdrL
8M6ym1qtsObeabsvmNc6FGpaKeKEJMWbzWRVu+kTZexSViyNyvEnOVT+8X8xEhkqdgBMSIi7SHgi
ieY+3IUVxeii/JQfhNIci6uJ8L1NQ9qlE3Hqb4AwaMGv0xzHbNdiBbLsV5GRPIgcqovUhDiEh+oo
8OQ4hMeEoe0UY5cx3pjQspUXzHx2HrPmp+e6ay+iLDstrT5kLabCkGK8skgo5K0XZrDXDcq8PlF/
Xl1PRIVzEFOMC+yxMGFHVwM5wsqWnqxnjrV8+IBDA8T5yyWYDI8xiCNfXGXE3NwnJo8rBciD5zMe
O9p29FSNlyGoRu6pYOY2HMSLm/XIngKAQlpdhjCE08a/6AsQElHTYG7BRA5fOvlT+Wws+nuQffyg
XoJEW/jEMs4p9fQ0m9eiSHYOhjT1UxNOyTRWVrd74D0hFT6A2Q4p15aLCkIc8i/21meilIdhgONE
O60mt2c1LwJZbY5BOaA41a2wuODG4A8gQc75MnD2KNt83IuAqg5eIdaU3nFH0nCOD2GKasCSKKh/
2UxyJ335XUi3qjfJ5ias5v1VXM2plj3yo62EgzPdGbp39WRP++j42Brxc5DR/ClTbmSEKEUrZplP
dPiEChY9ND+Z3te1zATgVjnSfSc46NBQ1MAY0itWQKDimmAlLxQTOd6Sssnwl7un3+SzNL+V6uBA
MihyH46HHUizAE/kEefPQIoBVFrL7vKCknHRBk4Mj11tLSF9QJLiHEotP67mtulMtRbM+9Q9dEga
oaa2Hl2D5MLFAyOs6Xst6qVlq4AYqLk+ETldiScs/Pv+D63I+LsT3cMYUO7lnvUK8tkq7w6osxzH
Fslu4MGg04DECdXP8U4+TtX9MxC/CYtgNEOg4HLuwTBvgMl9UZ/22xxZkD98pUx+2enUthXiz2Ba
AFHVjfh6n4fVpRxZQRZ7obvdznTDTAC46OPzePNviw0I6mypIdOn8D0kXQN48l5xb95O1OYOcdkN
SuFqtKzjuV1cdfjMF9NdQfGF1HlJwWJ77ttU8w0tVsBGaC9ZHAodd3Mr5rFDtlRw0f190hLxTykb
lGG+WFKTYdJ+d4OmBSv05skFzE6scXbPl8xZuS0E1QTgzNZiCmcTJW2LLLPTnz5NMaTN3UEDbbMt
7PhbQy4Kj7vthaJJlJtg4uR+2RTT8witicbu8ovtBb67fovIvwlsJXuwpCKhpuIPbYwtrQkvFsro
HyY3pVqAVWS5DxxzAs45J9jFro3xiah4vxErSbbhL9kjQESyX1Yj2yvmMv79iPc75u4eAo+Rawv8
4754/CeshIOjD6uyJ2ye3GsmMkOnBfve53FAsgDYmC2pU2SIGGW1Clsg1OAIBEZDc+8RKdvL7OzQ
Sem6/uY9j8xqkyai2Zw18chZ3U7yPF1nNv+0ha9JJNRtxDAU0OWuchygx0s97oLnPV4eYhFU6LEB
MxKnAst11QhEMtZcrIyOQ7Cr/5QbAOnCC3OyJNrwyOQGNQzWsu5PQtMKl2hCkrrGBWS94bICgeYI
1IG8QSXDeNFL3hSKOnZbLlhhNHssnWKlffxEyu1K7b8ipGDvzO1C4vnfbx1htlOc3Ri2SkCWChJX
JgoEUQoy3jncNyUZMrJ2/mPiCxFBuslIEmHl44Pp79wg7MXHpdRkQej2HPP46OLbh77Vcvvdx6DR
/bLCuTeBAZJSZQ299r3LB5Ja4i+nbObMqkQkYtGhnavWeBc1IsXH1y8/ZsJ1x3+cHEzw1ZfjPS1C
n3aABtA4i2kiwgSM+8Q2tcZqO1VVysPjXGYh4yQbqO2tXddPpo1IqOp367gMgCut+VX3Xgwsmvvz
GyQBuBz1zEt9JYy0AjUukMycyiR+vN8sHMXTuxsWmA9tT+YEvZQjfvKvQibG4s6dNAFrd+K97A6b
d3YlUk2V9U4wJMZE1mjt2NjRcPFfNcBVptttVnsUlAGB8b/lFqn9Uyu7LPIv+alVd55/GRyQHg7S
oIY7K4xPq7+q7ah1I28OfGRoQ+2RLK40P8TdNkxTrPLsHiwyyiaIIfYV/4n9knzquJnaiAv2oLTY
1S4G09TWjOQcKKOxzFULK4rVD8NjnNwUs3Sio6FjLo7Wypa62GzDoNHBMt7Vw1AJZEPY1/7Z6vEu
lmhNAdmt0whbUJW6zV+7afWe8QqG4fl/2WX2QPtlCoQceZt/WTmuStcWFz031eLDQYePARpC9Fkt
mu5c1fp/bfaY/hqqtuZTJZjmcRwvq+WP1Q+RH/07PD4gT34sAI1qT0IPtc9o9ixobDG1/khfsZhN
TosGxIaJYw9G4YTft/2KZ5fFuwi+4PXlp2g/HVM4NTJtSJm8jjCLmv9XXUwxs0TXRSd9waV68jCg
rTH+nraXZw7NX4OTLNLE2m7+VEN7+71knzzlMZRuuDvR6qm/R6bo/MRcPihfTzFc7pUbLNkU8mie
aOOH6f8rN7IfyjWeZu/SiawpGIhG5jiYc7UZLfU0a0jq6SwGWvpDwsMaMx9GXRo/uRmXpg/MFSv0
unk2/X/ZVbOJYDjjogQ8QduqpzJaQ+vXFCmGNsuxiTEXCRWbVn4B29bC9yw011yWG+ib7kTKbKWm
LPCdPlS8D8wF+yi7v5jEgHos1eSbJX4HUzrG4DVf0+pH4EFfW50eofHr1uHhIpi5mELD9SDQh7pK
yGiXHEC5kLp6LYZIZE2v8l6qob21TBNbiD2sDXGxVUxd+YbnAte40nD8DkRpvZeUG2m61LxLduFR
Kv2CXBwOcQHsQwA3aY7hEjRK+/DmhdU3xiEhfZ2Pwn3OQLUm4EQiRvpAyi+AaLPiPADJLnpRZ6yY
uH9rlaCm1ztb5h1f2eLGNeEQCw1mxh+W1Y9+BRreVajwOEn6nniGI52kI5s/Ju/waLzbJvj3l5fC
zRmw2ZKSEmWmuPya8WqNKaKhcJxIk8yz9xKwK5ScORR9sAKKb6rjz1y7ByRhlQKkOG6P5kC+ydGj
6HWhU3C29jBn3ugSEKdaUX9GD+/qa3aasbJR+Cs0Xqc39VT6VZkVT+BVxGPOLyvv7qRBPgEGp+MM
zBB+DZz9KEPRcjQThPBw/PNwditJArzTFe+rax+c5mYCoBXT7uVyR7yIkGnlakcbzvPHc6yUZGn6
w8rm/fff1Wol9RusmtOLU/qJEGcI7r6o4ugOOWvxUF212eiLGHGfUaUPFEaQrS3UNKbR7cs62t/E
PsIuvNF2FV6NyuVqFo5XcnKU7ZF3w+I6by2zNj+8i/Okr/Ie3o1w6KSpzrqO9CIso/kY5w6o7yKW
ZaBSgoGEQ57Lqq5X+Y0veJy9ybkx9obsBryyazUicYKjjWLHEOpVKgugmTk6n2vV5OA/WKan0HG7
DHDLgRmND+JNvluIqaTP72/1TGm5+SOT00tCtfhibeTNNIQJgNfbCA9uZ/jYuDi0Z9Q2lHdq3Va8
qSw6er067cNqqGtqmDTF1nVnnXkPBmirzBwuGJQ3639GmPblkPc0f+BGHdykhtHwhcAMShMzxKWt
UiId3/dbbM1T06e+jsIkLFQO6w4VsUzqjm/7MMx13Pmmr13HPD4HFnH97qkYo9MxO6ewfsuTuJqS
n6Um5nYMzpRdRq+mRPslIfzD/0KUUM+WXd1ZTBc30bZwNlKceFdd9viBnqausHyvBynNYR3veBBn
zzcGQ+VqfqQ0wFhFtlReY7hUbUJ1vP8wlF9Kd8fmrWuLWaQsvOZeZ2Ct8sG4LDqPvGHfh0JEjgx+
mlVRlhomJB80B8+VnKzWX44Ij9RhxVklczaaWoLYoRBlHJv4es2CB6JGe0wpn/K3uLcC+e1sprnX
qNaV5nC80FWUmEwyj2hR0m23Okup7Ix/40sfrxUv034mGAGNBCzCvH8iClyjI1mB3Fmtep2YODfC
omaXD9lU+roRv4CldtvOuVTITtAR+tIKrXPmzMRLd4TQeypEWi0lHKtgDIEsjH3ddnZ6xe7wBiLu
69PMWGbCckkw9ntHItzT41gKCmEFBbUcL+4QzKwec0JUWaZ3/y16GgnGuWpVbANRzPAWqsHmjj7O
xbWtvdk599138o4xnUCoz023d8WwvdN67IrwbktkrvuXQty20Av2/pjZaftaARFFUD5Y7ZRlQuYc
KziGzLnXhP1XozfTC4tR7QMQDbtj0Sg1nAtgjJNB7azeZpWiurUM+p7crbr1DEk6/CIjfrHjU1ef
o4lE8B6rvep+o+0FPO9qiXM9Fbr68/HYCVcC8FX9HYYPhOolT3AKtr8f9i21dVZ2Lbp4zJV6D+PJ
04NYk43zYeMMisPNkEABbXCzGlqrTUcyHMl7y9asjrgePmTIemC+GbN5RGj5lo3viCXRJrt6uwLs
2qYZENnZOyeUV3BhrwLQlSHC6+1NDsUTJLwG5b4C+ELoQu+Y6lopHmTdnnPiG9hYcqwEIMURAKRT
xnhXmepNL9EPCbjFqUxLVEFcfo17tU64XbrGNKWP/zdZO28SUBV2H2tYNGtU9sDhv5YT+ChV9RL6
uoHBUvC3B2yYR9/q6bCujefIxXo5ChvctW7ccIaUjQyEdrekWpB4xJ2oHh4BPZiT0xB0rcxJuqJh
ZeZCuXCW/eEihHC2XGuQpgJFYH6S56VgpR4E78l5oLEtBPjdsiEB4hpW2Mh0art0BQiOYOOgXWEb
6m1h0gUSBy+jWmr8Gcp+uznZwvCz0f+1YhrluVaJ3ElssrUnHCKaNKC41qB48gtuLeBL1UuqCDRL
EFabhxWSnwdmIwZhuBKQfhX+GYs6WBntac0QiXjWup+xrYEGV6ydHte4mmT2kRqyu85S6Rjo0G8n
DmlpE3wu9o6RDkrAMP2o2LUUviVl97qrTENF+UKVQt7EyABKUtmYfNMDNLoB2jlDWManf4Vi3/Dp
0H/rx7E0oomQbYlIlPR1mJOj64Ti4LOxGEeJOqLvo+LXlUq1NSXGDVWGZFld92/b3p8pPeH05xfy
N3jei+GixAMK/k+TvpJkAbz7YlJQxoUxEMBAPAiZ4NMI7Q/nG+cX9PnMKtX+vJSuAZ6AsqRs8z6G
5mc232m4YqeOfcwGSmyxJpJJQvgVSKu8ARqD/yRTHaedwYJc/rtBxKNaSJbc5L9R0xFs08FWnMgi
QzKWUHlxIGrs7+qdm5NLYKtTKY9ExYffL36b+EYmFVPidi8KaupgDpLUPhLGRnnH0sf50AVog6QS
Wa3YlOnt2X8gfKFlIgH9yVPZN1E6/D9Nhs1nGcprpqgKX04sLADigJWf64UqsEyhaWPyKQRmAAzA
4CIh7xcuVhPdXNftxIwbrRu/+5+4nVP4qCFoNixIspee+/BwlnakcbQAnJ1ODTufjGSjIF62/xaG
8V4kKrVzPRpaLnpFQi8OH2Q7gmiL/83cAZlTwRURdIQ1JT+XOiGlLjUApy2JovrFpXPfJNok0Dtt
8TiQiB6ow07IVuUNH4Bt/U4N4gddBld+eFIvCkixNvsTdAlcCo0XICUNLmvX8ZQg9ORLt6yCRrfW
DVpMv7E6irYFMJX02fEutcIPY6KTIkpDN0MuzQEUOiS9BDInEOQwDfCMVOyig1q0Tdi3pRcM90e1
mPTBAxtynpU9dFN678nX5QuxyiWoAltu22kwA7gUdtrJs6dqD0qZlb1gS+Osxp/D/8RER4asWHGW
sWXB0jMfj3HOS9aCa6Snm56lqhliKzDZZeLBLWIZcE3c84/Ianw6o/kg3dZXpZuGDFVfi+D/pPt7
0drLaAWf2U0mSaz9MdFLfZg386tCiZNIDoxXwl6y5tL5I7S0HpJwPFGLHnHk9DHoqZFcJAzJk7nf
m5+9lKscj8r7RrjARs7Xrl74lWJix/h/uOOMNx+H/LeFlEoQap8irdS3P9mqEhdVAkmhhKDvdhQ+
JFqik3XGd97GFJ7MPNXyCd7WpISlGAyq4OPas+bj+yTOvE0u1X03yfL5BrYB7A85nDOFuSvW1eG8
kDY6qnUn/KnVRIgGkS7Wd886VbwEDCnC1Tc1VuSfH+mdnE6DlU5tdXCSrF5cTU4u4blr9yFXdksr
UNHgCNeGORGE2NJSmx73onsuHE8xispfZASiQM2yz6ElbRsgSbDgVqK6dKriJoV1k11K+laAqGDN
bWcumOpIjpuU2vDlSBFGPX1ZMLERltks1s3jwTaEBJwT1ddA1eEMibIDvL9lvEXMX3sSos3zhL9Z
C9zHkyrVBrubmUUL5gcqIT7lj0gqob2OIt1/YYn65jnXeqAROG5ir3q3iLNzgAM8IsWWyGsD5YSE
IRPQmmz7/PXyF+hj7G7WwwbAOP4xQwXGEfENimu7uub3kV/pggzTdBkbR+7naGmIiOYMDduG+Tga
gvu1OZaehbLWaRctXI3WNsnhloqJIy9HMLoHFkLkwdxKWfQ+B+FaHRhzRV+bwmuyoNNcqkwXlJ39
5c7ZhfJqRcT83q+N1sq2Fg6h2QiWRLo/IbmBkd7ND+hcUVweaqr4JCwRzk98vLR5wX3whFdsMdIr
FZXlK1QxU0m68iiYw4onZzsbD55bfUuGlKqUlc5TUjsG4acxcpmsw1TIfCif5PEAu2dH1qiAppxJ
65x1c839ZGYA3xoKvhRRGsGLWueXpf4JV13mL4NNDqGWLJ4q2hhduXltmp2GSGVDz6QkLg7T/1Aq
/Tq8PPD8KSkaqhJtrDYiB+9/jOa0nB1LxBJ65/FktTgKOOSIDi5S/+IfsArfni+LVEc4KFUFR+lc
vRNKK0sGQo2AslrQFhLSvd0BciujNZCCufgvUAR7cJ+Aop47Vwl2Hebly8zz37DzWwbVKdcAAOuH
YAQTuMSjfQFCi1J6+SoM+Xv60GFen4VAwcSUOsbxI76eW7vYQkyg8c7wKX5e5tpxRPgwP+1aWnNm
jIz9944OG5WQ+9SjePX8nBGWsWwbXLRMvixc/NS6hHoO7yYyOcooxSyYvX3r0vqGZsXf8wBLUL0D
J6+X5UlW+OqsugA28Sfg5Os3Hw/01kiYlvTgU26tZme2hXW6dpb3YzaeCIThfg+gqw1NfDX0eO01
qBvmtuZ+QXHx3LD8XWIAYQqEQSEsumJqxRaJHGdN5cHccfvwjM3KBg5tgc2+h13RInxtGqtCUnou
BY12LoDQBRuEOHAzlHIWd3J8+IAFtwJDqQhpFWeXswWLss1bFW0QuIINtQ4cc/tiqCPH2hkUqGI9
4oO/fCNkOc/flqQMaD8Ia2Yh0ZwS7A8HAAT2zkJ9rJVTJHYCqNv4MJultqFXDxUvukmUM70bdbOY
HPRTtT50thAg4bYdrkBl4sVDwdqaVocyeU/XXZElIQ4UnsiwpG4sV4b+Jc8tfkHQ/hpgJ2TyXl4W
ccn42DVkpd1NpJLVuScoyW3M+BbzYEPXWO4bKDpxGZvuj0UygfMhqCNzMscn85Lgzbbto6DlvhHR
03ckDV0s7zhlu8DInab6i5azbUsUlvwjayTK+eM+gWTgPCS5k4Oi6RAPEzW1MBGGnZ0OEDZwGoZF
Ft+pdIY8Rh6E+SBPnlIn7eVj0K0iejuQgNv92aF7xPOo2T08uX1LPuyeiQz8aIM4mRApYnQlpkPn
iREiUZClHOmGsQzUBVEpCKKMrDbhzFvvoUUO6sNcLAgfRfxShOi7WQjOAvQfrXpnNGSOQBuQiLoG
oVfg9h16XR2e+6Ue9FqHuyJGx4IIzuSvZBLt3QPJnYc27EkkH+ShKhM4t9DqzbqJKBKlclCgSeMB
+1mKtGkxSXrukkvqizb8+b8OepNXEiU3c1uZWh2RshgOiVq03TlurI+C9mlDhiUUrxlfGs9W2l/H
4eFyq30RtzCUKQc7P4UHUCAJkEh4w74kIsvWm2UOEsEdCFFDAhFW2WoxFppr6LSZNzWKM7URc+DB
SBZ+957VV3G05u1+Q1RBcMj3p7bJ859xAZCYQf31cDvfSJ7xtCVzfQ7//RIWyFtfqYXfVd7pNgOV
ZJ/c49TcfJBlhEjdbgJ3Y8b2lkMaS1LI+QO/Pyj+e3tbQxgu7GUIbVUULFGiqDcsyFP+44Fj9Z4p
nFfgnjhzTDy0dcxoFCuMGoixzi5Zb4uo/HtX/DLJsuIPRWM72l9zTrArwoCI3Sqc7BxsmHcvTPjx
EHeiU2/3HjXOSCUuS6vh6TsF6ZgDw6LFkF+y/9OsVPsqXTKd1KGAlYqKm7zg1IWoCeTV3Zfm0wHF
XOjGHfm0WNogDFM4q2s+8GfXpZ0kLzx1a8Uaiiu827wpeEfIAeZN2UUZ2OkNLbzZMZZO3dbVmB1Q
R6/awfmiZTzw01ZrVl1cGh4crrsK+j5jA7/ti/86id1uP1UJa2oBwiViLlvWxmFY/jNwx8efnF+a
Nxec1H/qH7UGXIBjBcAo00UwPZC8ADo2YX/y1eiZ35p+yJZ5oYJeahx7PzSCP+nI0+rak6Ykxsa9
ibOyzQJxDhS4Rsl8QNUnVavfDbDBg2Mw039/aUVi1JqR+amaCNDtbwlUCOeaF131nm0X2feDfXlC
3BNcj9PO4w23iCtA7ckF4IfvSqrlRPkHBWsUMeTxvFWEDi9L5TaV7yg0FrSADkjfOdEJ1dV2kI7O
yY0lPjQF6a/duQMI/FQ50jmJpvFgK6NCjvsazd4XlaOsq67ctI4cLLRrQVFgJzz20E5fO+Z1hKXX
fZ/KsvW9mNe0mJAuTwszjQIXMG54P46d17o2d2RM7nV2El5xZgN19jbKg2OcJJnR8ncO5SosClGJ
rBAdU3de8g7FReUFhnOfBCz4kq0ufDYMQxXJ1mZ+/uigcBZ8W28Nhd9fExd+nnrdiH7kn2uDesFc
LwmDJ9zsukRGExO5LhlBqmZTZMSIZmY1xUymu2oXl6qBPN2sJMT61BUI7FPS9gYkmPSvb/yavKJd
avptkjSZiQzDJOnHGanWzfTkoQNGV1y4tjJUWAt92pE6JcSPYFFZ863Huq3o1DxRYgLf4Ke6pzK0
958GiCDU6bcVu/c/ia1O4xKqNKLtPAeR7wDOkS6y+wI3FPtmolSRDiD13DbV9R9GwyTuXfbQwtrL
ukxLlDDxN+9JxY+jdEAhUVo4dmGayuQQyfIl2Snrdmn3tr71AaO+xaIKARK1O+5PlaLRet0EXNn7
OzjORC+b4eT3/lEYE6+GFTZnM173PzwhA0Zu8i8dgFSZc8UFKHDOKuo0/jpCDxKM5SuUN+fgrv12
x5mLVMBXsnAmsaWJQXq8MkVGzTm8q2tx3p85kBv8u8IeulfUomuqjoT2Pi+CxhugpxyKOnFQl9Gr
unlzm/RLqLG7pAJ0K60tZNEo9hEsDXOZ/v+hMNL3RYPnZ96PVp9TS8rLx2Ua3TloOpPN/aYhKbR1
zMTUmcW+OpvOvHwVvFtDwvJhZM+kGc3yx7ok3HEUa252etWn8VpUX0R3wih00BkpbruKm6JYxvcY
BjhN6grAUwpsiwPG0oIfsLDRNl7w2FSyUXNKBss7i1VlYBIafEvYCcaeeRgZS3h+qAgkrXdl8lV0
aP/PxyFqUW1FNinrgo2QrkXlLpEcvuHuNEjBmHBJ9npugvs9DGjCjLZ6wx+1VR2CY+4FZEwulBBb
A0Te9qPsE8A7F65cHj85vnhrNLDVp6pmWlmFFZ3hnshZGA3itZTJOAxlZ6BW+hpX63xnY/kJhbyz
0rXJtC4AG58wDz7Xr2HSEMumsA3XPmhU1BmNoxf8UUmt2Rv3pvK5f+6j1VrwEEbLBgMihH/KI1gE
T6/TFbXCaFo2EyUBqV5I9kBbfoOz0YvXIrsTg/LU233Ep7Za5uQFStNMB/pMkMpwxHWisUw1T47a
MJTXSJDuheljfNBFXK21eQeUy3PN7iLirY/2FbyhCaRCBSCSB35OvICIBHkfTvzPnlHkFutXv2+/
MCBPtntP1gcmZdBEgj13LdrAwnme/QiOpR6Y/MU2Oy3WJ0WE+9hiqqNa0Jky5NoPDqpbgWh9fsFR
pm/swxBsqFsLnaMyA0q0bI3YKhqWiGU1N0zH5G1MJOUKBFUM64APSmG9PyWMhlooqfWKnK4cAaa1
O72tMjJG0F3buNkCmCq6RrottMZ0sotUn80gKJHd3nElRmjO2INKf9+vsnznkg7APh4qBM3/hKVE
lUKh3AHue89rIeQWlMf9s5tEID9dNEsAoY1P8IR2ymlFX5OejXxE5M7RTF1DLCMbz27oC2yfFWIX
ARJrrsfFgRwBpKsSEIakW6UnaUXrY+rzK/983xFNhEXCnv/Tr3vGJdJkewh9fP3YbYq+4HOjkHD7
5f8l6QOX44kaXVRPGdM6TKoHWB1ZD7Pa/+lKqaW4dygchWvCgH0jZUQLFJZfZnSyGENydfWHvib2
g05knDOZnYSleHJnQthEFdXu3WHHk5T+HK5fj26ZPTTkSmkQZ7XkNmrX8FCDF4H1cRTkEXr+OThd
fId361XGAmFiHLzELqFHGT0jE9NRPjJCHn+li8DkNKItciBthUc/Nb07FJdJLHjHie/yaZ8DUbys
GZ8RbCByGxLuadift2QW4ds3gPlY9xKY+2Ov54Rc+ryyp0/tTsP1Zv+fGVlQEGsQAqXpmfZUoyt3
HYt67w4604SoY52N5HxKqAKbt/HRO3a9OagDK+uRVeNJy0OI+IBpGeE8HRSgPbbv+Yl7NCW26v7j
ePS5wzAiLYdOlIqa+ZRiX4aqVxvXdnFq9uBPNErievPKOmleiCs1SbAE+r+icanakV0NMs/bXTnI
38uHQIvFB4zXg1hR/jOcPzd7aRiE2I6ORYhrCdjSvl1Nsh6/r/yqMarQpsmATiMlJegsFFa2/8G4
+HGHxQ9BpxyUTQEVi5s3qKEWgUfBaM0NFE0A9jKfx9t2wSbFxx5haTdtw2ul95gQxiU34ZBIGDsq
A2nYvJuRlZlwbAanQg39OuGfP6/pfwi8tQDKKruDzMdjjka74PlBCXecWAcKz36XZeR5tOdqEO3i
BpueBnE/egxJGbuZb59YhpwCwtx028IJ+RGTZHzVprP9TelzeP11JkwBCiy9eNqjH9pLJ/Dz7UFa
6Ny/uz3PyKRKkHOeY1jtXqvCrcpfOT6H50NDCxRhSITfpUy9Rc+TirohqDD7lTclTw0O9YFwZMuX
1NLwDQHc/j1R9zXOvxavAmqC3wStse6tpjHzmfpbFAhlJmYF0kHQbaDha1bCuEVnzHvx2Sw2sVpU
QeakJk9d6RxKNm3e6qLAdgIGpurfNSYsUIqwSMsgzhIvxwpJJOr6gC748A3ocpDEcVpD+xIiWhds
n57RPj723A9jZLx8gYRhXyJaNoWfnv30NWm2a5/CN8u6qYM0Qome2brwiSk4xJC2tN3qXpit7TZr
qBOr+ng470/egKQVp1GICd35mEnjZb1mqccAsrkuo3+/RMGCjVVqVyzW/4tcIyKcykGc6iQ2zgxC
ZUTV9VahqkoQ+C8PfHQ4Pitg72/YIAeqxHXOexvkhwaSkY8UWEgaOes3mMV/vmsO3DizvwsPsZeB
QTA5Gd/z4jvUPC1sRK4t+G1Lh2J3f58S05O2J34AtNWNclyGCkr7lSjoqx80bGTfQ2tf0zwMRPZk
MeK5EhGEiQJfLGEjWCInuoylPkXujMxFQdkrqg9vODUaj2FsHS+1VkB5tyr4WKJwvOW9MJ7Ofq0o
AVdbl48x7fYsBEFwJVEQqBhuAGzPM5iO1Nt4W2qvtN94+NGKHR814EUCY7OVPCvnQIHmvPJPziWm
r2ncMZOGAA8WYBff31FlxyHhEeWhLFwTUf4jzN3+3ljr49+GoPIx6OT6XNyJwEwid22U9UqV0NGK
gerF6jml4sP4K/GbWPyonELZ5rrUQIC3oUwje187HzNsKOoQQ4O5fwu3N/KUhDrbQeDSsmcWeKXU
qpp1bne3gixNrEtWJg/jAuQFIt6qyL/CREQU9wyZtNM3X7hqBXXzgLn37rd4hX9Cl6BC0+aVoZRU
k7dH54WYpFO9r+Oyjz0DIrorDPpxs20w/D/DZgygB199cHTwr0bXwi7XLwB1LzrtvXOA9QurmNNg
lJjvlZ79IEJuC7ieaxxR5qwnYSFgrdSldd9Rz/LB/MwdCtHSftOUHTzId3u3dMaJ1AvNpYrOiDVv
Q0CB17HhXClVWxMLDT3vel6nQjMh7rsYdm7j89ZVVMUWIe9qA/lkXcwya/4Yb9ZqsA6YID+A0m5w
a2NCPpbI03s0zsE0/+GkCJuoDRKkGFjcANerPmWWh1DARLy0o+m4ab8Iw+s+KuUarj+WsDQu/+fa
MbGY1hjhw25x3nXOiX2jP2cYpP/LIlPmDRvu4Ap2luku5zYmkZ/ZhpdNmcUQTu8gZvhmP7SOxGX8
5PYznxfJ+YYYIrW6fkOv4xYvzm/WrF6ZgVA/5C996D2FloP+jkVAMSUzEH2pgmhMJXaRdwfx0qfQ
l1M+7Dc7wVMuSz++BkU2jhkqSFe/H6bXgHDkuqpT8u9/wbgTGlSMcNbw1+wa7SCKK2AktqV/oWs4
i/C93zzbQr57OY7DuX08Gqe98ZaEgesUBpy3Iud7nLDGyeVXuD4jrQDHjhAe1z08j4jmZEZA93/F
OOouR9WQqklweGZNBAkVtWFNhe2JWfMkDYhkfnJkhnVmZejETAKUKJGZ6gLkx+JL3VCOf0AsCGks
GwPr+gIBS6FFWp3ugRAkj2rPiKS94+hTo++apcU2pzoc9bifJwfTpGiMCKR5+skoEH7Ido8q3wTb
ujtjUEKdgu0rcio7OK1b8hy/wEikyZWTbwzfXWubVF1Gd9smSlhrIjuY/UgLm+/gt/hQrAUwMmQ5
yW59dNHnYgJ/duruYfstuWhhA3ipfL2KLOs49uE6igsBp6EDPCJKG9OAw8GJElFuG97qO3HUUUFp
vTie4yF+qMCNaO4pzQfwhZHWa5TbpcTJFoA57tf0Wtwnjy6xLJPRIAOY1ua2yQ6Kkfq4THAEGG5u
FVMgH+mAjGWLBpVn1/3FxC5dkOtoUT2TCngnf9L3PtQB5EUNSnbR1ZHPTrdtdWrrqnHx4IExXynm
zUCkhFcfIuwMcN+1oTacFE/hj5cHQd54HJKzspDIctlydDGolpZ9RcyWBu+IJuLWX6w6ahv8WSeW
8FTpzR2fysZdv25l628wOcMI9wZDvwDux2bphNqRRsXI4eXytu2PlCd7gXDK4vP2quldoYQOn5Rs
Y+YuxGCh0XtgolaY7bQQVWW286pDJQ/KfU7MPESIknP3+wqseSWAKFDYnWDVor1P/PA76U0WhrcZ
Wj39n3ESSm5qJ7DG7gdlHBxD9oA/JyHIHzZsrTy2GfOpDASCRGy9WSRj7z6+N1xHgQ6INdOaCjtn
gU+z6ozXejYKVvBenFkb6EvArsfbwcyqYP49R1TV8h/F57RSfOWuVOCIJqzSV0cbsjpl+eLCTPag
Qo9VEUMjQNSnz1f4CYfFScNP7G+bQs8oCOVm9Y8hmPQ6zQEnJ3Rled5eHSOuYmeNOWy8JXkY0/6Z
kC3NZEL3fDVYNI693/mOdoqHSl0OTAHlStHUKzztVPNdLPEhdTtFCzpreJE0xQGHECSJfD2AyjyS
1M2pYdY5R+/FE/krR0MY/TSjC0U9aD528CVfMFZJAHl8tuqoF29brbGOku3CaRA6N2FT9eC9FVDR
MCkLqzSMmbdRbNQQgx1WJBlzBekpPGNaKn73WoxrH5zc9UoHsndqNFHhujrr3Mx0e3FgzkoDR1zL
PRMwXA1Xpn/fqZSTionJyfOrCvBJZj8W8v8+glGTxFUNHyDbqWNPXOlXqdjaS95RKZU0e/haNg3c
pzLT2MAecYMrlfZdy9YmiBTlc/sKG622gx0j6sZO+JlN//m7HW5UPCzULzqVsJcZ1qzXIqkoM6J1
XwXmu81vxaxpy3IkaBEO0cpfKGPDhVc8JX+TBGnBwAT11lW+6gQCPanp9CLWHs4t0dPs8ttvsGE1
BNXZC1sogEF+dQdt7TqOQv2QXO2bX1GKZ8zbZR+gAORJkabZ5NEpLM40jR2/XRSTBYhKvS8F7Er6
Bm1f0whACEmyYve/cmhp2x6W0C7sBwd0Kf9uWvgNyCjql1RFf6QwML/vpJoCum0clF8BMc6SJ8wa
sEsTlraOengxFmguVKv/xVBfZeDgo9s8LaQfU4kF0PTN4mrPF4muLlNtP1+EI+w3wmGGbEyUdZAy
avs97CSn4o6NZ4gVm9jydsZs6A/LUpob7q2/QOYbnz/vDzFEpBsf+OcO/fjGq2HxIGpvx3UCmBLb
gZ1jiFYZQPUfuBHP/iNDIGUFtUtTwMNQArYVSm973xjDG+UG1zV12B4InFDJnCauGDYwwZy2krsb
fRcxxiFofnI4rbDuTDct3WCWqelgPajbB2p4iyIlcke5sxYs5SkD9r5CT5BtZFyu85oYpFX4reE0
Zu8Z61k4TP5LP4p4ok0fa27/xn4Ap8V1GUvXZ49F35pVRt8+vItLeSOlkkW4FNWsQ06//ce/w4IQ
mMDuuWdKSkmQcBS/vqABgoztUC5WfdDY+7Omregbt4GMMPMgE1T+FrHKXZxVpOcZv9h22Cw4yu+c
ZiocKu89vmtS7fLiNrKT9XQtELMmORTLIhfC47znWy6jUVVSkECXVSwg8Gs8r08w1tpRNZr9/G//
uDtUOjNPwYK1qyyYxcaqqBWJCutcLcJFZTPbHJ9C/GYRNTRkz6H7qJ9V55mv8k2OAjQX7zmi+JLi
ypQFp5PptR209GYjuQ9XZOyyil8hT3WLEDwMonl0VqcgpFNPIGprK7iw/GK5CEg7CC9HpRyoz4EU
VlZXLOxR49TOrmgu/MkHROQvjW4XO3WxOeOxTC4yIPyw94AGBXVncUhPuLMTCMdjCmO3pn9hzRqD
Odq9z6KTc2A/huXEXQjx36kdiWff0GcbX1klfw98+sKvaMBV1E32VPIDc6MqiKZXz6oZcP6lEC5U
keQscpJrW2zU8hATva3wLDd2YRakYHGE3f9h9EhoLQQR6uCQFqJuZ7UqDjZrk1FM8XxOqNBb/hbR
OmmHEjVU7Zd3+gQmhBz4XkWJHvCa7QwtlPVPvy46i8UymDQSPYrmlF47M8MN0EBMLYEDEa7l3xWs
QpTlgOeuAA1XdKkMqQfJlVzoqV/ow+GuH57vETmDeuutccU6rdY4+EyEHDbHNlZdK06k1mJa+g9S
wfuQWYIXMhjmEUP5zJ2UchdeRX1ouC17Xdwu90CG+zRDHQ0nIH0aVoQM+Y8VTt5eFXiurFAYehoo
laoADYysk+2e/dyjM0vjKZxbfwjU4CJvYY813qC9VfXcPn6IKWUPutkTRExQwByPhV95FfpI0DmR
j6jTvUTcdkgKaGi0TEvi+W/bmdadaJ0pgG2O6p9UHjJXdJe+VhpXHCVucrWouSYkDvjmdJ/Oz38J
WnCe8ot3f8PmWl1zAYhDV97KqhBqmvIZi26mL3cKMn+HZORXsGpMkH4jteI8sCz5qE2NSba3VTbS
3X3BueiZOXXpVosmbov79fAK2I6p92DsA1M/vkALry+ssAZ+3vzdT1g6WDAOTpRnS5g0b7mUYu3R
zOPAddHUcD48qlqk8Q4cI/WWzngmtVx8vOSCaDDl2apJRcWSQ0dcrGXa96UEzXiqdHCAT/6xIYLo
JkddLiRaZmQjg5JlDWA3Lx4reHdAVrdA88R9DchrLAReNMxhAa/xbGC1IdoGyDRw3rThUUhiWWOO
HJ4jdmYNoebrWg6XhKbMr3LUyJdxz2H0yGraUlemdq6EigZ4EODS6RnTATZ7k8fWsmZI06T6btGW
9uasj+p+tPwltEsfKwHPRRQqjG90KCiBVDtp5bOYIObjvCRtvo5jLvimF/Czv50rB3Bqx5OkVWqG
90qYB1JfZx+MR0aARp0OqJXS3h/JRHpwrWGZWf9Suw7qcIIU+Tuq4MvTwtvTeQZqGVN8wWWgVeMF
1TRVCeTYN22F2hbvuiAv8UBxJP5Xl/A4FXpdYXyQ08Nw65qW6164pI5mwOsM+m7R4vOE+wSl/a3i
NRMd+jMbQoCmfQSNNjdEKuAxIaJ9HFdY64BJEdBFsEFYRsmIYWzaHXCJCEz/yvalKhkacd9Ud79B
S8tdB9tOkxPhFXFfplLw+/ZLyTBO1MENaAkdg17wzdjWWJl/AB4WBJVI0j05/2z8O/KQ3QKzsTt5
1ikFtARAYuIBZi7ypE5p8yDfR1vOtJZb6hTeTWBAnaDyB7cUB66KYK7bcqef0JblD4AgvpYd51zL
Ty8de71voo/ARS0zuQc2bXo11iWvBJXkB6udMZp9HQfc+PIRYacVLbYz9+f0k50qaLTwpIptJWUx
czGAhnZi+BLp8kLASJUFrY0XNV5P1FWj9hiao0mW8oIzmqXjFGU0vHbnGqzEVwg/15haEbCdub4X
6jF03/eEBbfO+6xo39xjvoePdctbxhI8B6w+abdFtXxK18RSPUZ8K/nLs4GEjf8HquNebmbPePFl
ecRuyVzOgjeXlwEkfp5nbkPIt5LSMarovDQFhLSI1OBIjqVkQSsFx/kuhXxnG822h1SJLYHBnIoK
9O7hhujOBwhORyfLF5Okz+U6WYY9Ez1kYqL0XYnVqryuDcH6HN+y0mdtXJfEDXMw7wediLPFBTjZ
GbfeLnZE+c/XByS73eFUsWawrbvmzXoMOfpa/Ht4er342y3Az4tOpyrP5Azd7Ck3iymIUxRvV+7s
Fg8nwylkfEeOGSPuEka5EAQTCVYxJHug9THXbPrnUoa9wS1ds/VDrglpW4vqKfIPWHHKbFLJLv5G
yHmD1IBJ6znndB2pKJkA+HHflLpxtJTtgOr6X9rnV5lKLMJ9kHLpjj330AWVR5TLM3LP07JwPE68
Zd/RGb+MPvt5cIb81m759ooM2IKn+/eb293RrmsAy31tmyfDlmqIo0fMoOTJ3NaRn0/OH0ZBNXAf
dHNuV7sNOVPn0Rnz1/qsMFr3vx0blK2JW1WdKCPvLPkbDMRjQPNXinYn8ck//KQTd2aIfNyRky7d
xyz4EAM6sKAFJyDOTui05qfjXyvl8D9uPBDhxX093ThDblRsHXG8Apfv+EigmeFazAgVLqN85egY
A+fbkeIXscHl3z0otrJ1uEZCtdiTDR5ssqqB0Z3tbxYn/WYixgqcHj0m8YS0OA4PU2LzzubBvJsQ
XFdi3/C6p4HwauH+vdVnnywIsvgUPN84I1m9Ei1b9t/ZGRlUwonfcqWaFxPysX+RspHmxeijrRNS
Xyt7xy/my8ejDXbOwqvCp2CsTaa5L425sNmczrVhqAyEErQ5rEd5VtGcUii7DmGH3b5g3iDTUXKz
erzIKutgU1o5oV+h6DSZUOvEbRobZxnekeWOJZFXVXXpc+Mh6SkeU331TxN8b7bRx3SiC3PPZlQE
b6KinUliMB8UOzo1e7fMpTPh9GNY7yHpcMp2kt7IUlGLkQXlPkfN/UEz5ZNf5b8aBKYxg2logSZ9
eAEvlRPqfLuxZrpqI0mV7DDaApZquli92JSz4lDmmdvx8ez44v+CIIBIVirR8PHldSspTN0bUg1n
6xzZkM0ugpAGyu0yh6ol5/HqBJ+umYKn8XXOSN3P9K9N9Yl5YafaFzQkfj+1UjZND7naoIyrpaaG
Ld2nvUPEXfgL6Y8C5TLhvVigiyTC4VqUyTP+EHGJkgPBYt0vTh51R9xoI7Db6qyVusr2UOXoScwe
WTPC5Rc4z0z/AtaYqCkf+UIWN702tAR9ceMylA5tbWwN1WbcpU4WUa1flacz1voI/bEEArRAVhrr
j0oFmhSXZQf0jzUU5P/CURKYkOmtE9PHlynHsTpNuE1mXXj4SMR57NzZ+/GhdEvfA3GfWfnc7PpK
uPmCW/xupzjqaum2CSUQC4e88iCBaOPZZosXooFtQSDa33iNpSSVthc+D+azHvOxFhs+K8K1ikZo
vIdeQqzWPr9KPfb0P2O0MwGBNqMWgc+1isKjFGpHBnJBqo2k90WfcBr2G5gOv+6+6ZTBmaDbx3P+
dOPAJBA1WK4RD8cedd2BzmE8cZFk5xhcVWcQAk5f3jps5t23UUFFULCIR01/lS1VnzP4V2Reo+I0
xTURAy7+nLXocgxA6k5WAHwR8UWlEXUBeMqifHAl7PYYvQR2s+eCorGnYmoItNgZrjadGYv6PsmY
0Wb87M6yimcKti/1qbPX3eW7vaeoIyTy2B3FdXpDW2sNh9Njggh+F/Jai9uotzeCSgN/I9Bbmk1A
cpSioM5UBUL1537SGdcgjarQnJHmVlSrKLwmTmoYcgAGk4YyBmD9u5JIE4n0/dhXAe3PioUoS95B
JdgJeHTidSOx9E1Vt4db4CLbsd7pUq0+IpIU5QtRPF2syCYUwyJSrWcNrJDl6wBTUPnLPhloygOy
cLftfeOVLFYeNF0Z9KXjsbkEOuTa39GKIYtPWJCVJQHRmGAn0cGzkqVT4W0uaaPAAYA92QeD2/07
dzI8AO2h6XZgDznlStgHinOSrgvHVrXD8S31e6y8UT7HRFM5w2hZKAMzzVu8tjsXt84uWOfJApFm
XTZRb6jiv982JE/zoalpXC0kxzrtDTA08LQDMqUjRMzhJ/7qGrPFeoPZuR90Vd2p6rUiwFxlvxjW
b505RfGyIwRD0izTkxy3H6ddfZw8tWl6TW+ReFDSOGeq550vm01r3dQHuXOKiqBfUGV8b/WT3437
KvrkHek1+ay3750Y/mlGI9JDzQDXNVKa/+VMQqwhdEgMFDuHhnkvm3hE/G3OB5Ja6iBx4mLiM+ND
SsXrOBcN3qy2/GI1c+0/uwNTaA5WoygUjYzgONoiGruFSA6SR3fmn/JtWuyTFPI5Hs2LWkstOx37
W+NvP9ZIxh4ojn/t8h/cfuHrSK3ToDkKjPLkqDqgWL3wm6z+7Oc34UpNHOVetDbDDCpX1f+lrDWy
VQQR1GigFfnEc6qvbowQoxLMGOVdwlwkREJ1iHCCgpSGAgAviu+SxkAb5MUYXVfdfY8Vk2ky0K7v
8REEPdh1T8Iocwdlh+glruXRs45bl+dOqKmrwITTFvImj+MDkW80h7Z7f+6bKkAWJf++o2VOHLaW
mqi4+91QV/8Tm2ESlx2g6EXRgiNAHwSonxUgOaGLu2HvP9WE5sZYzfXnE2s2MvVwr9+z23yeEjFJ
kYTK9vrgMJW5v7T6J2KB6nnSdNKiaSKQ+zfRBUIZRSijSymh96n4ZPu/ISnx7OsQNjB1Vr2ItscI
ARjGbjQnhA6uIE6F+WyGAwOYSSEbZxR4vhCb3xRcB//o8lsxM8scWmz0LC7yWtm8kzJqa8tZF9mr
lLL5oNGrCPGFiibpZxWkpxSYm1ykBI1MhGVJA3AWLb4MPmbnfrbt0HKQmlzcPoPUdZEsQXp9a0a9
lqwSQWnMIvw8BuDm9xU/mhe6QoLXwcKYqgrLa40+0u+i+oZU6thAyLZ3AvHSZyarEgGInUp47lgZ
n7ictWT7qhBHsmWdSSbzyNstO23BvQDDCGONIzxzJS1gFS5fyXyztrf3VDJG4OxK21HxOf4V5fQz
PNKpS28s8iX0CyTy0m/MHuJJ7lPmCraiSr6uSR0QcNai/xVxFiB8iAxLOHnbUyQZs3uj+XPwyfyY
BYT9XD1uDAC8aluKmxFaKTornch0clZ4KIVzhRLKBnbMTcI547fHdQ56PwY8oaB+x3PhQaswB67f
9gmyat4AuV+qR6IRQicl72Onh1NPkhG9ngBvKmc+6PYpBRhi3d9eT5p0tJ/ZM+mrSylFph6zxRan
sixVJxBEBp68fC3zAEnL4IVYqgBFWGbkKxPHDUAUuuDsL1XXIqcE9MGRwb15QaavEel9S6zNlXot
5DOoYtrS8U5qXwPWkJPt8d2hj1RcronY137CTnHNuMw+8RnUbma3qqGiRQWYG0/t01GYLymMyS2r
lQe47vUtd4NxmdnPZg3MVZ+GHnjxg1kY9Gb19Cl9Tg0dwcruc7xIqzkW8T+BlGwjSL84s9jSBVEZ
IZFb17qu5Dm8h9iTzqnktWddWKJucQTjCNKkazElrS6mIzZnqjaEnesr8GZh5hHDNu91PwGe/i21
ATQjOm2xpdLDcldY+++4bG449qMeYamnA11cJI7BcdWS8NKsRSHtRdvhFaI621QgSKPA65PguwlL
rQ49kIDOqekTHG4NbI2roE3UHb8q4UhP2XoU5IAr/4MKpDQxayciVkpq7c2ubG7LPqYMbT4vxkNY
McA5im6beF14OIr24OdeeCgasQ+mUGpbRKzW3dbf/vDqReI7DI7PNnqVZPbzkTKe6O2VDcJc4Kl/
4a1UEWIbD9uWaHpcZKiVCsI4v4m6YZEoaDTJPWw4PEXJOaOvQ4TCUJcqydT1AvBnqtywxFeJ7KTU
WBd5c70CdRVrDqoYpxb+D4ZDSRgyWFPspI/PcMWwhTtaZyhoq4K+ZgpIAg/7WTskEhW8Sbzx16yd
D8hBWTHqFyzDUV8HJhQXWtaXE4xdYY9FviKWj6eSojDJQYs7kh+MRwQSiNS/iDMlR0mcLvglr5fD
9XPQ36xkr9Ke+PSXMBvRCZ2HdQTNPT7sP9PfPWb2ULmDCjhp/94nFbuMcdIvctyYDSuZwJ6gf3NO
pGe5VFOSv0CN6IHH4VhN3BQ4GlFG8yPxLeb4QZC0hI8ytArXbtIqVy4luJCu7LU6ADUyoPHCiAkB
MbRpGgFQ/muqTJWucYpUz3AkcsMSjRK4QzSeZhb0cwIZlfR6obX8IWrTvhxd4+x+MfkYgBLM/WnP
zxsCNXihfbOj3ch+SY7pR4tMf4ub/TuLcLNMnbY+Ei536E3C/+j9w8FDaontSeAEzTq2xrlUI0cN
B3Lcfd4AlS4fwYNNgZAN/1AQc/nwb56Yht0Tj+R1QI1oqUxKnoPjlrq13qnh2iWS+pzOIDFDI8jK
FO+6F9xpkp2HljRrZhLqrZpYwnhSJBE9yUlXK41a4opb+JxdaZRsZS8WlSkNy/owBEwndONdRBp5
UacFsxEc0UaSM/G9vHi0GyleSplE2dNqM4+sXA+d/AM9kOe36lRTn9iM6QnNzUOF7X7AXB5d6/5z
1l9MFSeu+owX0af2udXC2eFYYQJPuVgCrx5qN5qZhubTIejTm1PCJutmLaWKb7xgaecMVStnwLYI
RkrQA9mtdoOT4zMhToCvkG0uw/UNriQQrhr3AhTWisJyuYhmsnGhp7UW2bzudGvSABbVZnVATDRM
8WjTM5NVnJyJMF6S9/o+Z6wYadUkhj81VIQASKzWBGRvgu2t9RYe6vBR3tw89el6OxJREqnU4BCh
/P/GI4GDZZ7nTrdqLstKX1ylg3ACNJamPta8z0xZRz4fnD1zgR1lz13KKygp/htgu/6zw+UhAK2X
a7BCY34Pm+Dh+9MP6skNgjGSi1W1h1HnyaQ8blEDEmSBoZXi2BZeYiBo2CxueLsf+GXclXxrdV5p
JLjBVcuxkksCwfAczeEXdU86S5rGiD7PxkVSh8hvtul50ttR7YtL6FZ+KK+svPDbXuN4GcckMcmi
Mjf1Xk32bo95GgyhHRzn89SJb8V5fOxMuUtYxO+DH/6b5qfi38TWLHLOmySV0Kc/cFIXzWiffJ/A
O9PtNBUqCzp0S84IBoE3qQ2EK/X7jdRJQtxA92393Irn2dogbKiQCEWDsutYRfgKIpisBWoqaa2R
vnyLB3EzmwBi9Y+LpgWJ1X/AixAv0Nc8q0lqKT+5xGhaOsdJB7bkO/wY0HHiCmJNbbyNqk+vnTSA
GB5GN4fOKhldPgeA+ICGy4yam3VhlzaVqubvY1ehwjZ84b2k7qgxh4ml8J52wrZIwC3MH68QgEXT
9M8yZcPj4MHLh3BfP1uWaqI0Gv5YMXKGCQXS7v57o4Slki/auZcSubov7dEzYaCs4ZznrQhUl1eM
Rsyn/tlULFvqWvMWoGKGOWSReQFLkSzbzRuYlAlFLfBFVEy9k7e2Waz7Jef7YiLxBnmx8fA334/U
35c5ngXfif7oo02O7VaIy1kw2wueILagdqSDvkue+MWREQbj1BEnmyTGewE4DMx2SjOEHsBSbs4N
4wlQW3HvL4AxD61AwRxDRGVGjg6LKo3/zsp7H5qeDhvvT1gwe9OuvSLrLU2Kvlgy3/nvN4uG6ykI
s0868qTAPWK7LV2UaFsl608rHFhvhYJJMdZml3cMXnAPzyekqPSJvnTfUy6iAj190DLxkM8LD0cH
ohtFfQDUn44hmAtjbuVZdY9nHPLUMQuyAf8dYYryNTNqBhdnwIR5gqRHbzdDb47/7rapVq1xH7xz
94DrZ+1+njv/7dRoYTkUEg2DxgE039rma0X7UJauD67SKVP+rfLIfe3jC4bgNR2ccZRiginaaJOv
krikn6g4BBivJ6YsTTVFbh9Ui028ecej4T7i8xH/iHFIO8TfsP2vPtZZ1Gsjyh4R69SKT7gVXj4Y
z2hDrdq5Yph1tgQvgexhI0HhxyUUR65Y2L0bdF+KofIe8tkkvVzM6Ldi88j/lDm7alvMosJafeVO
8Ua5rDbQoWrYsusqRNKCg33QzETamJYcx0xOzEC1nfJSkGNkWV75cHvnFCNXW2TWmx8Bwi3DohFl
Wrcx0qpgO+bxeiuv41el32kMxTXX6lNBN2XFKZvumgAh0Llhw2NqEBhK3exJAxEobgot/GLVYid1
oYByuQ3LszWu+vNqZjDhCu1fzktVXIV5U1y7ct0puqA/+bfwf2M6gDONSGpF1moTvOSgu/XKmKew
BiiiQJiwS8lf00HWoYk6XWxj/WrQX6klpGhwCbgul1NEYTyEdht7o3d7GZvL+J0sG6/TWsTvCr85
/i2HL1P3wROl1zEWqJjVaNouwQd8tGgtUVZqssueuhFQkTjyjsJd7MxWrB3hkhPkMizyFCwLUvod
5bHDDxIMRc59sPkzIXqZtQk4YufORcvVYCTw+bDV8YNPnlbNzmf8gExLigC+zmH8MFyO2aQuNIp5
E52cU5mFbpwWf/B4UpJ30CdanNM0SIUSgVnE+fk/6jApoC0VoAVv2651iVZn6iqjrt+W3xDp77CK
cDKN3KPOe5xAqLcakk7JWF3zNSTlcLYrAPsZDJeFxcnZt9tVpOHBf+2cgq8NWOG/koe72pfs+qQn
oqBK2JazMpW/hgBQrBf5hnPXhAf5qrZUgf3c+3bReiAoLTAZ0NrJ4t0CqRBHr08w1Sv3GzeNNcJL
MTaldhgKUcA3VO86hLrn4tg/1V4HO+Hz561XCxIaC+2w5Q5q35btsqJQ8YCEtri6uJS1F1SVMqYk
c8H8OBAYtU4Pdj2dmdu2kqUEfjli3iwZYRAQBetZl6w36VG2ceSMGdRYMbhUM6cMuH8Q682poiWD
0itz6FECf9hAb310ikIM7DOIw9+3uO/XRylZ3BokRYmhew7seBy4Zpt8xrhcZLJ/SV2VN1BeV1pm
lU4sJElQivGKxgh6NhgewMTBV0+5oUvfyNzvBjEKIPt7U3NxT85GG/+OvKtANITHkweR/nWfbsgw
lg6L+TuLsG6yON8dOueZHgjdpoXfCYFejM9W0k+lpfknQTg+/8CWZ7ZPKYPl9bd85+KnOpCqSpuO
EUxZL/L4DtfHEOTMSi2ddC0lVmHqI24nueSw3syriykzdrxUxX6ispD2CT1TDNKGGlPWfIhoAXQX
FpCeLJgVV9zE5a5Y9AXzHjRn5EMUUjjiHPWXOEkT7EdpADmNe749D16n04yl+YkxWC8C9Efowanl
cvy0J9VK1pgaS7OgfpE+5mVh0PYzqqzlLHG8BY9m1Pxdkbqy/Ex1FeVOKY1lRd3hLZwg92zwF9s5
Tyqy3sEb/564FlsD2k56+D84RpQvS1kKIVwHOPZArm1q0PoEnVB8UyMemp6o6xsXtGgn7uDIEDpJ
tKHsWCeev41V6iMjF018rFvMlqMsB4DFUCBtL6xWVDAbK2W5WhGAn9ObAHastkvldLY4J2FLEXQq
4b3fThhBzmCUwpfPUtlbP/O5Pco+xDG8orGMFzbp9f88lKXziwRPyZaPrkSXJpXN60MtlNkfzKOK
kKQ28BsgSGaR+24Rkn8/1dedtSIv3sLm4MNnq5l1R35yzFIslYe6W54ewUuqi2+NTBqvCZc3buEQ
yXsRURtOZpBPhLZhWUgDK59X8pfoJz+zYk2bPyzrcQe6MQf4BGNvN1sHzdSCQ/jdhSi6srpXxfUk
P/B0wd1H6GfSRb8m3JKgSOqdm5GMPlbt5YZRqUUyuKtYWoEUsB2+fdPJ1eFTWLG0+zb90xg0i/z2
bFOO+wanYieiQmEWvdrfmpmNNxa7ABL/Pi2LE9/bCwj64XYi4Aks2Tm11cxoEoatG/ZUlBO+f35o
XgguDja/UdQgyvUkrn7RbWHVyn02HRLK8zZognzKrfeNGniZFrxmC8+ffNQOLlgmYVjhTN9ES15p
oZXU//OFKOEGkizoOtBPJ4mJH4iWkydXFSf5CIKQJ4PLFG5taqZImb+pdulTvrL2JfOePY5ddt97
59+5HkSheQ3iZz8OMVMAxdeZtyxguykwEwiPu7BLPaYvtFWmLTmzOiSRP24C5RurxQ6/1geY5ipJ
ftxK0t30l73K6GbFon7ZIls5cmtV0X4K84hwrDWXALGpPg0NS2OAyYpsRNcf8SumzHoMl4rlsz/j
/8GSxlBWJtxVNzruPyKHYy10IPKYmIxS5GxSiPOAZRaao8KEL2DwqtgySmZqJENU0zCYpMceEFSr
mVDBHbt0jhl3cw5QfFY7cHD/wLPu2iKcqPYRVFYpbM8W4+zJm4pyRJVvwyf8S8MkYyPkeQvkZ4+M
Rx58wdt5XKzO8GMUhD0zSh3+pEt3YkrF7d9/VvW+b2uLTOA2kP5Tuh2/AQdNDVxOk9YCHWiLTLDh
nehsFfpCC3z322OUM5lV3GShZDA/QvrFrHFwAD3+fRSa0wfKpbe8uu3a3+aUlnR5GTqYQgGvTXUk
IWhe1TeD2t6LWjB2wLApKlF8y9Ij2dawAhi4UHfXH2cML0cwa8wy9sJepakuxQENCCaSwmhDu6kx
679Bv/EoCbWt91ZTXZcs18StGKBiBS6cSZxE0ZKrjHnSYO38a2q7VUKTvTEYIRnLSdEKc41K2fJ3
SZmLy7Rhjyb8PWPqPvYpTXHhd4ciq/rroooCl2c+HkY4nOftI91/gZale7bziu3AcbDGgGohTgRV
q99jMV/kXDq7sjnPparyuMAeqyQT5vFmkfrPfkWZ2OYXjQ3P6ItwjA/tJFJndTa7Rpu+asL29AvE
MarRL1jOJtEFrgePakeAEmiv2I0rTP699jpOnM7/8mstoEAFxhIzEIVouku3nhVqFNThIE/xYulI
5Samx6E+J5uk1OMQpRN853kdntgPv7yBx9mW+0BOGRITkgnKIi92OiHO6kRXsL1QhlVL59KW2CeC
z74364I2KTlYVpGQuRCuHH+cT9829vuTHiAI/AcpKGlvDfA7GVna72kfgvjRE9ZzzBK6z5422VXd
MLrxUcKpOu+SqZVlYhv+uvbUEBoJwA2ZAgAKj4OfvxYNJaXG1z8Vzivo1x7IagvxL4Q79IVqs5K/
5Gojempxbo0Uey/Srw3+bmqWomdDRUll0EU/VQdmkC8INEL7P4IUvXgZkEGBEBZ+mLFsXjIslaBl
Q9kyeqEPgrCt/hc6NYwVZpqDzsZg4HWPtbAB+hSvJ2ljz6CTLV29CQvVnNvw/QVLOwk9reclyWor
iB++fa+jcE/X0Hx/6PluO/CK16CPs8lVZ8K8ncMDz7u7bdZ0PVpH8R6cy+1YERwOXNSTMXUKjtWn
cxuLViO6gVO7BQ9kIgLuaqmz9uOpV66g8GqNZsn77Jo/5tF9K29r3vryI/bOL50VrRdPffA2okm8
QBFxrYLmIHt2UE6jS8GmlRv9juNPI2iM6oiBYUiu3/lO801P2EcIMRWJ90b4xlJ3EhK1yfSmET1e
doSE5RBUb/glSx8HQqq4ahe8s60j7VrrJSD4jJmy8SeYdJ1bH7g9dTEwdbUxSu0zmarr33iwHx6l
rvLFckI3t3Ph6MY6xfbb70GW2/m0/yxH2dn9MDey4eQz7SPo2fibE76N0TuG8oySm1yjntJl0i4n
kPif4KiuCtPBJbWnnfk2I8tuZ6WHI0jdiq6+TVWYpGit+juzaFVeUwM+u3pPEG10A8gzWDUkP1bT
SlfBHLGr7Mu+jEGZ1ylarX8C+Rw8Qpz3KowIgQfeAI2ioC6T8UYiR1JrkKBzIDj7zDz+fWkuHB/5
kg5WPNLnuO1FuGGxR2kF8maYzcaHaA5d8SeEDneWXHRUAePH5VPTHXmxmWavKTN3H+VZxKVO05Iz
EzA/yo3jLVsYYpLrVFRo7CRPDmtD5J7YKdRSZZ3km/xRQ6zaLslnbGbN6jB7Qd4AWLw6nK+kQsqI
6YEhBeS0aCZO2VsVr8qsCP5zu19zMiZD5AhCTt12rIcIf/YZOEUjMjyTAVArYFzOPCkVBtj3eq/Z
Ecxve1NV7R+bDdAUWL1JAdMuBgGVfClmJbUXUDOs5vsHUqQyoOCxzMyKEiak6Ql5x6MjwDqWlpry
LAfF5tAyTR7QhVGugCkvGUe2Xp5RHy4cv7W6rgvctfYXjijalGNF1ku1ygylw8Xgkv/cD4bWobrM
37Z53tTLhmJK02hES5/GTJw9D26/SuoPhtxOVjAoty2rm/bRmZwoYqDaI0vWrcLEA7L8AiaJu8Du
yifYYR6bKfGGf2wvZgwbUoPZaLi/47q/4mjr7oj0zN82Cl1I1o3mob+C2JrwL6GruxkXTI3pOccy
U1Sz/Y9DfZAn3w2X+uab2wefTtqXUFtohgCXVfImL0DjTw2iuU3ZmR16RVKbtM+3R1j5MiWkv8en
qhXKf8LofBx7T/iWzFRfyIG/5xgTIlf9/3+cPXYQMciLnneOfVm39mjWR9ZBaBbVXl6Bc3kxMPlH
09rIcUGrOBvecInIZowzyM+Im+CUL3+IMdB1d65LOFgsBaH4yVBEHr5YMYwB6tCmV7FhbOEmemFz
XRcCP4jfob+sAg8eJdKFUu52R/L9oOSo/ETT3q6bjU1eOIy+m++l4Ccu7tL3JLSebhFfmbQE0Axq
T3zVpf4Uhav+RSY5VcEk5CBSNSTwMEaX2dGDhC26Gn/fpxm2sloQ4YfBhMzYo9VzNpHNFLLOgosB
xjHmDhR060ziQ5coBUpaE+OgSI49izX1ut7mt9w2pse0CVnL56bsCMtOh/vgEj8QKP4Iz4OCBa8z
ddwVoVPLdgPAwTatE8Lz5SpCCTUwRNVjLufPq+J5kr8u2E4gMaUXPdkH1VO89OcRgZG++3JeGNxQ
b1Oi9Fje4WbU/EZO6dQ2cnYy3I/On2oiZH9X/lSYOn5OEV214G0u7EZXmGDPdAPBuqcZkn8+6SA5
xQ/vidPow1lfSY7Fv+bVPCJVkc13aehA9x0DKJaNgqkhWlIyiV5upW8oFYezgReScX9qguVlJGio
OY7a1imxNti5jhFJj2s4mdJG37N5GRjixYPd7Ap5/ACEsrwh6/Zc1nNUvQdMeDCtSHtfvLas69o5
JutSXXbHrKxxA3NiCNuy1GGGLr1lvm+rBKHaK07uTGg47SIKlI5Yativ/h48TtOmjGUCeYjPKy1i
L6+vHZdUwb4Aq9dsAz2KxzSosXgnBzQgWX4H8o7BFtH9lrZY/C8kEtZ61Nx4rIm1qSskPWmI6avA
9ihjDXjWYvB1mq8diX2m7Upxv+emI4D0j7Je8QnLgdp9rG/ItF2G4wS3J2lhm38VVPZhh4ok5kVm
+7uKM4Xa0/B46eFMqQtm/Z7cQBsRFLnAUFSrLEJV+m9ti6Fuwptcjhxe81+fLsHoGVKl9yjaQsf1
C2SoiOY91C9vejc0U1SWUnlRFepGzFxUNgdgkVzoqn9JYX+A6FZYDkrilxz5DlfPYVT3qQur7JJw
5Y9EaBDQ6RGefFLA/sJnarfT+w1M5Af6T0JiWh4eBHthadJDevBGKUm75DLGVFl0gRTG4SDEDz6m
vdfEk2Wm6/5um2rQOjsFInLximRmWg0PCQcQBzZXsy1bBlLajIdpx6LdQgEe38tB4/tIjWloQq3l
LIr2BPZVnp5XGmisT6co7uSdjumsuOUbjws1ZwUfFOAts8BqWzOXCEeQzS34Ac74e9hGg9tiyWRp
2xqrWTy1TJJOvasSKvmOJZI/FacRKOv0Lhz57yzf25dSxXAnvUAWvUZcOQ0YkLibqJJx2P7Pmbnv
j4JM3Hl1uJrBOuZI5TYLYs3TQ7L+VzAVd3G/iooQ+6TTF0kXlI5v2yr12Ss5vRY5XyQJTetX9Ahs
IekqHfw2FUp82vU7JimBY/0ZQoA5hJgsf3wI2zBNKdVhJxy1mX0Ks77ylb6Qwlyd8UA5Oslt7w8k
fTaTPB88p/rUwTqwEkaN8TOe9Kd8IjpoBQnVxJzw8Ec1737J9g4f/utEjYD94zZ6/v6+/FUidqmr
FWKxl/viPWTvXwrxF+sT9RJZa9GJEunQs0T/tAlw/Nxd81qd7BRetyWW6eX9c11JOF0+vWyWKYLW
S9yr0GUdg0vJWUhBBdDaDvyNFxpGS9oFhbCqVfQlCjdk+A+XctvDuSiGYP1jManZCMXtwk3H/AYn
kFyfDI/rPafSS+1VELqEba7pGD37r+T5NuFoeR4XkzLf/BzvHZ4M4KSNabTz9DJUz2l32pbKIwP9
zavFAt78Bb9bDxw7lRIotbHhs9AHG5XuH7/M7lSkGXgVGZ7TzXwKGujtdsSeR5MiNtPA0dL8898I
w1PEuEG799AkntY0fRMixBH2kNpS1ittLf3gwXYUWpxz4Ieh58QH7c3uay3ih5uI6JkFABn4vOIT
TvckvQ0KMwXTaTG7QePjmRfQcDEngK4c6azCbZTwmrpnwUPovjR0tYR2tODXW3dBcoj3w1Xea22a
ElElVzTBWbFpIBOa/sacmxD1Y1QCQgZvLP2rYXUTbBQdnIcOCydyYyPxdP8zL7tPV378f5WkLDiP
MEJcrjCVKDEqtHOioikSFlsYpCRaZRhE8UkWdOUruwVIomCrl0IA2YyIPdAdYztBP0XoTq3xVXcE
YZSs2sCdVFYSXXaMw8BedK4OkqIZYzFWyITuUk9jmzQc82Dbrk/9A+C935oJj+69qOYHmBatoxvj
ltTTMR1YVtMyG8uk7i+P7KBE8Yi0eVEqLs45OetRQK71r0w1z2haUye3VIhAyOtoZtcJAfI+qFYr
nrbs8cIr6l7pwcMElRpjiJGIUg07eWjZtSTtwx3e3VAMj7uThu3Y7ctbiAKBtNjzwz+CqDfiRZgp
7l5fTp5Lo5yhopi7uynTI9Ql4XIgFwE6fXdKxgZAOTWIP4IXIN2OSqIibv32akpZQu7I/4ocAtCg
e/I7wOuIAlLdC8rP3dQXm+gbJ85pOsa0Dm/SHjMqXAo81TBllvve1WJgaEkpuHx/UuyYl/nHeBi6
rTlQOZcQN2VYv9g7P/FLTFfLs41qeiBzdt45WreMvlhsywy+9v1sBxcq0MQMsc6RbQyfah5cn/MN
6l73waglP3pPP5PNlI3W82/SdGnVKah8HYprnCD4A+pufWwouHEDtzF5h/NWq249EZoPP6DShyUI
qbmkuYM+eiMLfVG9BW5ktCvYaSz1D/QBMG+BrUA9DQ/u0j7nTpUXcQkyB0TxdRuO/R8ghPBMcpob
s/RnxNpMwiIUlD3dlmIVQIB/iqEMXseo4mgrmX5OB6FE18yeLLRRTPKgRInVfsdx8o03g3KqJSuT
hTE4t+C6uavey3R9XB20ZpDeuLG/uHaRpLA1FFV9kBcvOaDh5TjFXan0JRE2ZsSpBT8VRPI6c18C
UEXUj0phtbPWFog/J/HeD6Dv59xiJ/mzH97JMKmvFMDB3N6vQ8QEX9lwdiLlSTuX0e4QJFbIOVum
YFv5IhMEoQmG8UpHlhQcPRl8jUuomcXGo3CDb0BtUT00wUbBuXiQfK8s4sNgoNNNGyvnuQxZzO2E
UQJbcWt4GQ6pchSCd9Wq4pFUKqPtYyV1+gX9Fc9cbGW0sAbfftlAtp7Zt6EUDDxfaIqTE1o4lpxs
udJaIntpu2exBmCcv0e0eg6ed/d9fuatZlksKo2r+g2jAd/3yOsEYRuv4dpOatbuYwI2OiQC3o4h
5QseBH1HokYAdfT+2wxNX/P18+nKoWifVSrLVV9f9aRaObnkFQJkvQzfEEj7QQfyxDAPcYU7lXXW
9vFFZ0Ax9BqtaZ/T5CBl9HvR4ILvUzPzWbsn08Uo50++zJlwUhU1EECmsakPqZ2/pYlm1V2PtCG6
X31XmqiE+9+PQ8oEe+YzCNf6bP81zgeC4uEfSTh/RRrmnrkWk97CM0YqFbTWzZl9ndFxLofhtlYS
YMeLQUmja7Z28YMoF/Ls5YNHQUdsa0d1Byc/ZZgGQJaDiuIhQuHOhDZCybBULGVAP4e92QRy3mE4
o4tOw02O/gJJ9J2Hzgg/qkgtQZW6LnqVrrygyVFkYS6kS/oRevAdxBuQj3glwaZQfRYr+Y5LwP/o
9aPkEdNLIfFtcIZmIshGNI+XFhbwpatfajLlZBM7hp09woqyUDrLYI3XngDp3dmh/M8mNStzT+U8
aV8u/xxAU/NFwi56zPNy4jqSwghSJ8aIJOYzt6yVwifWx+0ocaxQRm3b99Pe5TtoWOi9ZdHbSmxN
fOHiPa2UW66tyZm5JdKz0oXu6rbJyiSF3rVZq1vIdsqxcZLtRr/TmTdI0HfR8nd6+RmeQ3Q6uSlC
RDVSrv58iVMAhmhAsPBXW59bbKwxlmYYeLWY+3hYEYrdsqkH0YN8Lwk+0zL2pLNb109Vwd1pFCfr
CyvpKy4CUV6b+MUhxzAlOmRxTRjg1a1eNQwaa6eZHWnoNGZ4ik2svrahl5fy9A8W7fgzunPLfxh3
rv8qREBfQxyHSxKsNoTkXviKY1BB1ccIQbK8UnSyFazcBgjG2V0XY8TQvq3vH+5OXHns0WoPPRKT
xXkr1e2PaoCEuVSTLDR0LiQWwDUpqa+DGnFh5zVCvZUNDjGgb3uYlSIfGvmXDGOya+eKsLz5N8j+
eVuoDJFjYRyk2MNYXOe6QVZNk/yGrwIEuhUP348/SFwNcGi8X/xEjNNRXp2oPPnrXCKgxYiZyR2P
ssBJnXV5Dl5zqGRqlscVniyW3RIV8myCwOa0FE7VjYGiRqe6aLNgvGH81fpdOIBelCLNqtUFmx8S
MUY6BrGZCRwp7EWLtuE74dNZG82/wQptkagNkJn2rntEmnOK7ejByE2MplZUoQm+gzTCQ3vi45Yt
uHUjttLDoy6H5mQO7mvuMBN66bPvo/TE5a43K8w0Atj7I0rop/KLCUeLjn68jfXX+aa5sDhLp+b3
ZpxX9Ew+TLjta+vVTa4uM5HLaelgLS9zXw2i6PuWqQrlcqaSi2M9kpZpUHdOJ8BcEqE6Fh1DosPC
FGKi86ZpyojHB9aXug8jD+O3gf0P43xE7ukCG27WYcdQYLUbzVa60+MpjZm/4F578ggEzCpJRRIC
i43QEbYC/JyNVCeDoRUhkY89A/+X1bcGQ41Jo1jVLu+yNM1mUW3psGvsff1E8KsVD6bnQZ35xIL8
dTkJmI/zcKatk9h6qQx+k/ViQ9gtTUq4wKA5sRXaz6QiIe7Mt7z0bLVJFPipzsuRweVYYEQqBbyf
5xSWbSqI84RuJO45l6Rf6x5/uJ4ToHvj1B//5wlKQ1X6G4GB8X1BLdEFEnRifxvg2kEOnv9WmK/h
HAlGrsr5ditA5As1eQE2e66pqNvQCv3qsKqaRcSc4D214zVyH5LHlvlrO0lu2dX5Q+s8tpMu16wK
A5UoS5mlkm6bVvzXCbeI4/TcjkDjjIQceiWFf+mRU8hXxyvTiAkGR3G1tvJKFft7HeakclFA/yyT
Fs2ZVn89cPrdnww8P5ejGkq21L3Z8HWjSr0GDbpOgX0XN9qzHFKsCvfww9SGmNGnWgd+vfNdUICn
GfowVARV6WyS0QMQlJ5dkLcSCgvQ9Bc13WXHvYkjmveB9qb/lPOuZ5hiy5DEDRFZCLJ1XaNZtm4P
bhTlzrUJpd+veta6p8WoKuh/iwc9FYX0Aumnm+FAJrPrDjgBsRiveIYFXZ01+oA5pY/GcitZOLz/
d08laMNhaRuPmuOiCz6rpFxu3D0sNCP3I0GxHgVzUpmKKnmcV4PR5BxIrtIUr5bpnBe6qGQyOC89
FGQZWpM5GFKyryHqm1jiK33XNkWJNMKNG7vFtvD7MgvKWHq6+O4tA41D+vVFf3FnxJ3nCItoB6xQ
Cj3gVfV+V1GkjxUQw0kaAopDaxrTTbtk9HKcI/5TFPHsk22ftGti5l2l47F0FAVcQSIg26owzRqw
D4EAZLDp4lSmSX1A4/z1fW687fxP2ZxGDkG0ZAyPwaRVe71l1kI/Zd4begNdlP1m+RFdrBDgG5D7
84jJztWdks4q7+V0LxAeItL9NlA/aU+aOAerlxQNZo4Zkk5LGJbpltQqCjo1zz78BW116EdiPM6S
JAN9/Z1WN/OyyqI1HEgXtM2/y6YYTLLcaUaoISlNQwPmlDgU7bYpRS31Ge0wu+IYz9X+NSDu7cqY
02FAWsqYQA6TJInbD8psmxG39N1bzg6VpsjA7y+O+3Iw4D003JVS77pJeWNmNSogN7+HGVztaJJ6
VyIdEd9BbLPCOM922lmvWv0iHRtsDU7p5vZO7lgYD0GwmOZUT/2vJLKt1I8jI0QWzKmLPgK//93V
wpumaukjjgx7T2PDuyaO2aNlBOKfVdlw8GYqw45izRRoQ2J5h/hn60Yi5m/FTrDxeqQyzl5fDrbd
YKdxoveZU86g6ElH3qs9fRA+/VZis0MfSJj/dgy6T5BU32dyx6zsr6t9F5TSdRmdBW+ZTeVPoFnM
M07SZvOxBmRPNs8EqHsFFFmxRc7JqA5whgbfB1Sbxx2Y2wF73+c5RJssmNgBQzDbode2HIva1YS7
4Q1mM/bvwPXojenyRrsjbM5VNkMGW/F6mOAcc0AJaAs7R2oINI8U9PfNXp4hgftyBZHOuMgrLXpZ
M4TtfdDc3mH2PqjrCP8r1jBB2bL7rjSB6J2fk3huAUka9sqFaH0L0eKDn0OGd5iLbzX1dx8e9/1z
qhJbQIYevTrsDuq6Urw1jtllBSLw94US5qk93htaaDUarQed8j/2RFGJk07wM3YXrkZQkMW0I43C
FxNNi7TbOVw+Bskv+Oqoc7xlwep9ydPeh7bTXqY7Ks8sjW4ppTSLdGO3TdTWbsyND2UxQSBxxO+O
k1rQNKcfuQOcwpcXDsAQWwPaa6Gw+IX0vgUnBVyE4WUcaEQ/3crfDorNw1eUZBMPbhrVU4H/NJFq
b9FKZDbUtA7SEsjq1KmJMT3oq1LpYvjaNKrHcYPNML9lC6rFeRofW3hdzGyI7z+vtcfWHZPoW+CT
z7ddw6r2i2vMEPiUuTvbdMR8ML/0cZns2kCPScGNRkF8o+RhuOHVk2zKg3Xq9q6jzCE4XeCK/eqi
lftXKqmCRTmQa+q0PuDhEcrgFc9/5fumbXxAduxfp9N8mp7UPcyy8pD57nwcp+e3FTAuBVGCpoKM
NCNgnoV1wwajL9WoqvcTkwVmwySJR82yAkl4IYUYWgb2mR/Mv3rH5ivmtROM5jkByDUZ7EX5laBP
98//9FpjO5+B0V7jld/qKpTCoyn68MoOIXlKc5PO0D/JqMFbGTV/7hAjSTFs2NUjrK9fbhB0hKcg
VsUUCUiJ4qbJINtbM53t2SCwZNEL71DmD0FmirtBrF5HOWhBLzRlJ0y9GTrVjZqEfUiEcIbiqD/L
85VtL7Yw3UZB8db910ScSVb1RkX9bF6pV+utZ9mXu7FTlPBL4xifrtwx1oxNg6FsgjaJ5U5A46aW
+2bhFwkzUtKqJyXqbLSLA0GeGqBN4OT1H1qR3Sl/bS8cj+x9bsv70kRL7R3tt44J974pssfM0Lu7
+RL+/rzs2TF7KPpU7dRfBWzI+0Dhcx42DK5QMCyRU/dKhHTJenpour/fDbp9rs8b+cmcDqzuGFe+
rM2wmgqgiMPtXPVANh64JxjIPyYVwbnj3qgLPcLdFPS3roU0IxUF4753jlDtgUHePMGcHqpNi6Gr
dJ+W0kuo09DtfO7zBS68+jKBpFlPkW6GFh4FHAQooRDqAfJiJHaZBDV7vSmrYIqDXWA/ID6LZAJr
KABptH6DLcfKrCUY84C4wCrOLGfU08Xrx+I7g0jPaQ+9xnwP7ov2TRmz7OBHU7KshQiRKy05vsFT
S6GM7R3D71z7+8g6nPcKTlVSpV29HlX/Aofzb8UGD/IRozEe2r+1qQJ0ITRGUhR5LGH5BbKWRQu/
Yf6/b+cSPt4w06QYPqhNjebqhpFF2lgsIH/Kt9dhd8DfKNEfsuz4rhlb6b7KdYLsDlRGhXdPN7fd
/6+jCYHhHJ1P9tiZ4WK1dS9nJkH2Ze9EVAPXKNDkXU1weshzz5USidHU0fxleDNLIjnEnEbIYQt4
xxeqOa7rhrYE2hb/oegmGo0p4miM+jaTe1c08EKu/UtddFfGUPi1j+Fw99vHz9e4j3mVxwGIqIl+
9fEzCOsl+gkKIy2TMH+TGmUtPAOc7/Iyf6Y5t4r8qWxzJeozTwYs6Gt8O/mWetD7YiofDjMyTbWh
7isNMAAocoPA16gzYk0/Z6AVUquyP83cb8nCbfG4bE0gwsXJe96EM/6UgprfTxH7RT023NyLTl+v
t36xo5VPmcmsSc7HfN0Gh3vkofJzSNjt2+DCDs7SEaIdnw5zn/zeSCve7kDh/SR4vaWU0qkjLFfp
VFj6NxkLBJ8SrQnnmlW2zB97NlkDRb+u15/mpMm2FU9QB2SFx1VSAOy1ItJnqE4kBg23uQAoOVaj
AGCguHiTjO6JSbnrD7aul4vBmen5Gqsk5irwCnXfcEIW9aNG735sSoJcjvb+ZG5OkgyIJVL92p70
5RAH0kq2ChUOvnusxKTLWOcMmaOJSz13YBX3pgf85DQFMKscx7Fn3yCTDgG2gp7+kxQ0J1PW3RJD
sCj3Qqt395D37sb++DZhd026SSMpcUwRl8cIG8D4bTnCb+Mr17i0SIbyX5xrw4ZhXMV9yG2s/FEw
t9nU14e64YVHRujmSlLPkEfatAIKeSxT3xTRKjkkFHwZAiV9FgnoL/Bp4+2lC+r0PYoPEsl8P1G5
YV5BGMx15F27Yiq/hnEqpMYGTB+k2HCG0/KMlaZPM/l1yYOfgQn16RU80NdMd/eYWMHWr4GVGf5L
9oFJo3gsmn1m2t0I2kHDNsS9g63loHwxwDDqVUV0x1ZQpiI1SikZgck+0P4qNJ3RBcExV8bdtyV6
yrAdP5PkqDiSLRNu0/EKQD3Z5OpNdoDba/mKug6CS7CoSX/NkrDFQ6V4Dpgar+CRB464e8GFKXll
8RCS02MQC4JptLl0NUvnW2ghNLextzJ6RjhzN4/vznK8EH956PWJhvr6l1ijqfygtgXNaPKbyHLB
Iz+z82klqGRV5PmpTSyfUw8FPRRrOz14ox46XQfv54vtDRuNrKiooXHXK1nRaD36EIKJpwIp5thu
hS6HTKA677J8JmkxKLu7QyW0Fd8XIuVQuE/Fotl1lBeUCdL4CkAaPjHFChqJERlBbWdF+SQcv8Fq
UdNloX1sKEYX0CsE6diPTri5mz72wTuO7ngVnEKJYjcwBgpl1YfJGAP1cnK5d3gOVDkXYlRjIM0F
DdXfWd52bnSHhBzVB/ZyCLlqskqZL/1GFSJVSPgkwo2N63yLyqwPutPGAzTjU36J6DLn+43Ikv7u
nwImFDbJvDnoRvLWyRCv7YsEYzEBLXuvSuQSFdqsBvFwwbz4Ks/WJ49stHBZrPk9gzD9p0A9xlwR
vNfntn3XUWyAlbR68rLygUqPcV6iORoWx8UCGx4qMF1kKfcHiA5QOAEXku9vh9Dz3Es/s5xeLMPm
r/hGg6oiDb8HHWSDPNoe5NK6a5miNaRYI9c353jWbEP81SF2ANcf49zTOfclGcCECOMYwHYigJSe
64MJ7/A95LQgFUDABs4vmQE1sgffvwVnrlbhgjuvCjq7idEyvvaGjw1T4WZ8a+OzicH7YSyzuyeZ
FIRtV4WkAAsoiBUbs8Bfu8Cc7vPaIhBRV5C68INNID5BgT4UOLPvcQeOLNf+chy3DwueTjW+c5Pt
2U1FdDexl+P682dzfl2ueTd00C2awmvn11Fm6RiLUhtgHvRmUNOZf90AbRVdJwBHNKNiZV0+Pupb
kbatD6J+zedizuQJfJHBUPpkfYYU6SXL2CIOjYMCRaOG87jnxOMT3925VEMRySqEJtVZCC2Eaaze
skT4ymjNpQ6HYI4V+/b8z4u+h4l8ubc2+SvpPmJnJPpU/xEDV1g3gQV+w2geEcmpvqiqxJBYv+TM
y+4nwx4Trlp8NLAhOWntIf61dVJeX9whVTYjhSfYx5vdCzVAtEE6v2c3K/0w8F6X+Vt1nCBpVB+H
5ZpweZr3SKepsnGe+Juqjnb+0VfRT+y1UnKxbRQhpbOcu9bGv4fedoC7kyc0r2Vg+nCQkVY2tZE1
ypu5C9gEs4G+ocNauTf5E4VWQgRZSudhruiXrK9cc1MUZZHiKC2swUY0mD2PbnVvGu7mvrfF3kAP
mF5VuVj7pc6MbuHVUq9KHp0OhJyEduDD5eBBfZq6DZL+e9M5VOo4Rd4Y3cGz+CT0nG1q/ES8SmLg
jbSZUPoQLrc8mLzPapIwOsGDDEg5J1NJGRskXubRVZDLlDamwQF8HTrGNzVL7c6u8xY9FUfM8r95
Tz75uFcVvAVV8aaU4APuesGMAH+bMBLXpm36+Bghgy9yQhoHgI4mn56bdO5OBSxLa2v+NLw0MvYJ
OidDnWc/URbdJuNDU1/aQ0lXil3LRoIhrXvQ6SMoitqC4OZ8f10ImN7W9m79NqtawmndShTQaTZe
Kpf6v1aucYT5y+LHP8DR3iuMdTTtB84NGRQYr/EuYZS/FeWEj4I/tZLISfG7cTCtOxCMsKmBWiE6
a+71gBx8CjCVPnI3BUM2/D+hho/drj0m2aM/IJgJNdO3i7dqYx9Ax+sfO9sqyWy6RBbGogEFfkoy
VZrxO4P3WkLv18SbUZI7vp5YbaanWoCl8A0LSEXYGiigH2mnUFzdD23RSBe7Z3b9mdDFPDyaayg8
QT+YZaQ0CBFMMQ0wb9NTA6mA++UIyadlFMzmIRkEAq+8dnq+Ss97uexVPpDklxFQyF9h68SgVXNR
4+JT5EPXkHz0sgNEyCMFm0L35frnCydWOaxn3LuVMGRCriiACX88+6mIay7OwAUDU8mTvIe/n+q5
y4JeMmDNMW7SQMnDyMqLGelWjrDXs8Sm2WhqJVUbrEMpxRqPnrJKwwHgaRPHoSgUo/fg6V0gSyVh
30/A70wFrpF66vieTxxNCArfT+PvmakYaAZE4EXJdsQ4ZU2vjLF6URiSHpZ5/abAX2Fet0bMiksA
PgRL2SllLAXS/9w1qmWGLcDFwW5N7XnaMSB0TKEtZ0DPWTA8oIbvZALmtkalRqG6PCxAGz9SrcTh
6KdkK9JPcRTcTRrfElHvVN210piEIQGRn9EruDBmPU1XrRcwc0YeGN+s+LeR/xHZeV36UShEWa9x
HKmlOYmWbrnHJMovmUY+B0Sl/7QgV/9qFdo+23ap7GXbHxTdqutcoiJfnkA1CehXutIEDmtJHvDH
PVghJo0BdzeZmdQWixPG4/7WrXho/fW1Yguybw0j+8Mbl51sRQeveZj4NBvtR4eK0Do8yYLuBohF
PmU/VQJ2xm8VnvOm+7tjyfV8x+jfHlTqFvwVZuHazgkLFY/9fLzsSIeBdCagrR38g82CoecUKyhY
VBuwtOPH2p9qdlbbaS780gsK80dm0Ucq2OGSSjGjl6ha2V5aboGni6ACPSe8qabJKRn4rDo3OrdI
3cQC3PhfRNl/Sr6xZQWBtXd2LRPtWdHuw5wzSTYgaGiNywoVCcZsYns3JqjHz63B/eEpmK8yDG5Z
IxLjMCQ/G/JmZQpb+5fPRf2um0TC7Kwp44jjtbgmHsGNnHKNYQQf2xxJ+/KbZR6f4V4qJROxjn/A
MDLKFuPSzr1tqniroaQ7OOvMZy9p0yv7k0w+XGoi8ZpZGcMu7tEXqRNGZgAaFBzS4E/4w6V0FAae
204rJOlae/zNul/XVpPg3x6OidV/qLb0sGBwj+73if+n8BL43yRF3ugNyUae1wSmb4iTCAFBKRgy
pWq5h3BA1J1QjbB0ZZsESdyaFSmFcK7KKO7bNYRbD/PtLpemwv+rt0SQq/IFNpTo6yDJW1IUgUzU
zQJatBhhQi/xtX29X7Xe/Yi8jbUpGTObQ0OoDkX1ILyreujReThYYbYgl4zCVsofE7S1pRwR4STI
oc8iksuKz2gDpL/ZpO7psaQmmVmSx1eaUjiqfciQ8sekycho8sv9ki1JaEH24qAUr5b543Hu/ayo
/vQEPMcsbSJap5Pww/Z52pUkDSrKBml0uClRfTzV+VP2ZGXEzaWMhW1Xtev1Tydma8LsluY2GQjI
9MG73bgV8DD5vfv0ppxe7gLcwS4TkIBKTGSAHkHumUCh6Telf0/QNGwDIRgWggkNn9N+mos0IuIy
1Zcs4KE1WWOWQOCBNvTiPs+38ISawjx+K2ZUXfQ4LCHFNEdyQhvisoat9ip2zZ6+/t6e/y42zYNr
dqq6+EXFI9PxXFJFdMwoIh6RH1a2aG/zJDdGbMGOgf+0f0/FWDA9wZh8gGCiLHtfleqwtBqIKH1K
HyMu3ddCmAyF/llJG1zfYG/5ZbwmslisreDhojzekQnj5XTvsyfoY+kof0guHwplVez9F773/5yB
Pb3EjPMvM9979GALsbt3DsIDuS4xPcuNTwqBULr0Eo+sXohohfeTdyVejZ81xacTVn9RmjfQ0HyW
niJSi9u5EbjFzdzeaLaWXqrovquonpqcte7Fnz/OaFxg+ISrpV80thHZ3oP3b2KUeuyDNU77daRu
iEaGO8jK7oToR3GLGMq5Wpj+P+S5ja9Vpgai+88JBUIgn5Fe5vj/N9G17EXI47GnU9GCu/NbWycA
IIDe27mYSI14Zs4CFdrPb3vntdYnZajxOF2gSmdWZ+QNEcRc3FWSvEppDzGhUUfcSz4VLwaJV82h
Nv0rNTQirdb0KTOmKs+vyC0IX+QKlaBHZKeqwp8dCXYXFK16yLMPzWGwxmgi50PlNF6yP5MAlwvW
QkeT0PnfdNcF6cTFmnXN96f0GvSTot9vD4Qq4Dpr5ebeuam25WlI8z4Q1VSdB9aYherSUF9Jwz0x
EPqY9BvV03spM1beRbdO5qYdv+ByOCinNTjp5iZ36wVqwU8Vp1dv8YvWp/pxVAJZE1pl7Sh1JvW7
BjpwLTEgzKqIbrWNSiw/mCz745fEb2WJsrW+3Bx/JNjb8kLMceSXKijDI80E14Ee3KnI0mYk7MXr
QAHXmCnq+jp22/ab/htFnp3RQOWsb1Fj9udl0+TuBoDxSfhQlt48xphlPX1s8msKZgZ/+qHV7FJ5
ap/TJywtHCBM2urUJBSQCnHlNjo5afJvH8rCIVBdNNEwEm5jQf8+TiLYmGNJEDOGxGkPogso70c5
QgYGpQoPAecw8vHmLu+dK50/SqVL8+J9LpztMTC90XbkmVOuX3T5qOraYCGVwph3ZikI41ok4Uwm
sF6kUoRAVgCJgZ6KktLBvPnRbS9mZ9nkLm/OyooStGWuDHD7/iqt1ZS2+QVOkngPGPfuS3kGi3b3
m1/m5GW6mryfdn37eFiYdOMzF+QYoMTl2c7n8JxTyOoZkylYaewMacikamioMyAbKDX7W0KGExY7
p6bjjHAUzvHYhsgnEqAJsin7JEexaEPtccoBzgqUD33SFCQXZSLWs2JZWTBQor5BCKfu0opcFKZc
S49jCjUDdSoPEuQM9WMqCcKpu7ssTpQR6LNDv4OVwsLGSvsR2YkjwXHai7QiFIVjgZiHxpTl5Wyt
gaDMgzRSn4uI5jnggOANCFrcx76urKrn5mUGXyVX6ya/LiDBn0UIGp2R+SlEUxIAVeseefFOkter
Z4c5EF7/eziFnsimer1j7JaE4Y3m4FsiYnmHWu5jz8ePyhdzP0a9qLfdFsThs87Axipq7eGYK0R+
DumP2qwRMUv/k/W26wEzzHTpbpZfCA067iDHBgzuuk6T8SqM4JVIqo3oXTIBmjCv7EjmXZ9RDP0T
6zWTQHLQcMVJH2wFyv+2TJD8ndkeuLh1rr4bP0Xfbi4KAW66qwGkOeoVrIeLaQPrlY1VlFyYV+nE
a0yLpKxT5Fn4kD7n1bJ0h46aiIYhp4c7OpN34ZcQDNzQzG94XO+ofsxn3Zl0cMzYSje/+gFrTXtc
4Ke0mqhDTYNreWgMYud/Bx5NTFY5qhL0WdEwAgiw4oAjIpzkDmdjdPkStGclvxHj8Zg0hgyXFqDU
5xhXE60RjHhR2U54w6tjX1NpOPGz5AOoYQ6w4Wqm61p2c7dTZzfn38Vf1xFnZilBH0q2BlzDffPj
kpfc4FGsTgAtkqP+XzH2m4XmTsk3ObvwcUwORNoqmX6CgCcNtLKFUA+z9AJvYi+dLO3DFlY0jvth
79KeqS1i+fO6gfohPFDzL+MeZCxgTVPw2C4FrpHtBijUzPVl+wQLSgbjVh6FVY+u/vp5w48+l7Ux
eAlO+Yk9pfySGTXXg3H+KDQcAHu7HCcWtl7nUOwxU7p9ABhosgRlQrpjryB2EpvYW2uFpXQhnOhg
wuzWTE62KspE1vwd0RUqvi9e001ylNIVdhL+hCnA1YYSbGaPspG6j7bsffsPMRhfU41/77O/FirT
42Vw++tJz6HV8TOYo2wgc4QauMqPTTrOKuiJFS/RtUeM1iuDU6hjvIbZY1uG1u0S/IahwnlQrnvB
pVj5wJLWpVsnM4XBbSEu7AT4ayOt0PHC44/b1o1nLewQGNwDFCe45dI1klpHE6fzI3wM7AFZPmm1
DYTYs0CqTuI8hdSYZGr94aF325+jk7BC0/uFDj05y75Y9Oxl9P1ozQrJTF2iK2umc8DcVW6gvNdI
yFYbspx9RJxrwSD/rDP7V9fgDD0+ZAoYYtCbsk6T2AU2GtSkE+H3WgafIHkdUuYyUwpVxVSPtVN1
5BsyYQ/VxXQWON4IY7vXKjdJ4goSf23WNIz05fGWmZPTrTisK/CyG3zsyWacO5b3OO8GWTlfK4Gi
n7Ss4w8n+VvMYS5ypyKdM1kbIhhfDZdeiVzrlM/JiCY9y3y/P0MPjbtR4WcrIhhKAa7dAwwL2kLm
+MWLhdEHXCcy2tzzd/tCmJbmajF3u33lrJDkgzzjomeHnMUXWzzgRzT5T2ykqcN11vqz31+gAeCU
3n1zacv9qeDFdI9vQ5hS1+sQRE0MUng/39vYycxdLYAk4Iofl7ajbumDSs9z3vg7UYjLGVt+bPax
YkVDkzUf0181s8H0JM2TdEHH8VtAYZqzbiB7JQ8OCSRTFLh0dfkW1Djn25Q7PTD5E45eyTHz7pwI
ZTDDnZ4jlxdLUN5ANhcW/4UItCRpLyg2Px3OfM/riwA63S+wuWrCPSRSnp6PMRx9/dv3vU/aFfdk
78Go6SRRDlFX4aISzPxGq3Ylw2FpUSXoGk3LRGeA11gyEYhIdwc5/FLCQq8OyX4ZNFV6jW9l/2IV
z9zRWjch4EQirUwQKlDr2ETtB3b4Z43QVn7LGDakyiBrrZ/eg0g1YEJjj8E3avyYgR0CidRn2JNP
+eyqbap9Q5R1ie7k/HDXPFheoRhxjOIrBs8vQFkzqfzUZ1EoDFA5Nlee4LgodgRY/14APiV1vaZq
ftoJeUWUuC/7hm33SZWXT/wXXgJWx7Zwj828JzK+DD0ESMuHQjRqJ6GE2dwt3MeZIZ4Z3DlwAvhx
5b/RS7u2+Y1+Yj/n3r4qB3Ogq2YJxanQNhhvekEDO4e3vDdl/GVQ0OxfwP1tOtZTWPqlzbUvZsxR
ghYZsifvSANIecCootRxrLOs5TvXAZq5BpD++C8b/JbS8suPbkVht4aq9oFBNYWldomBgRFHe93A
EoODpnCC8PUZFFLUPHGl6REbGFthsRxjonYiR58Me0sO9HzgrpRpNQ8PzjyQozRgBHFwVBlnqAjS
lkK6acwM0IgKewLkH655a2MV78s3U1FniGllGfJlzPqx/kChzmV8uI5Qw+CBz4cefW095QFFMTkG
5jZ3U96W7msFdDIVUcTSmJ2HVjH5lVUOkgXo5Gvd46vMugKU52e7+NrW/sjFfm2gLsb8P79kZqE7
wMZi9UrJ66nPhNwfD2LlMndE+cQBa4CNKnmtK0XvhVT8F/ttHSQZnAxeUyYw/wea07CRTfg89uHK
xhXkL1UdrkGMdg25nuM4VFFYfdrUd9OFnRM53MFJDsLCRxrwfx8f5KdzOiip41HQfyIGiOo1NzMJ
mZIfQaZ5hsGAe7bSyhK+RJQz+4B40OI1QSowalbW37Wj2iMLTUInv+GbYaFQca9Htqjljyp8nv58
rv7gVmd7pXRnuxETYNGeyWpuVVbZDm2agarzOrQL3KV20yOoPH6Fw+bpKRtGww6VTANzjQrhuBAE
yiYgAuouwgy0s+N6p6KdEKt+xPktpfQw2e9jNV3oV8UL4WYpu+S+Gbsv0zRClpPK/O7RXkMcjaj/
6FI79pOHxuJTZh3kzNGzP5N/GJshN8ekPzAO6wA4cfBNNftNrBmkTb4zrMFmK8Mj16OUK8SB7qhE
VarnY7Y5hR3b1zVH8b1RQCQcOh9ZumIa3qeaZ6xx8WTwmWt6FODWa0O0FJ21+rDtL6zL6WcIakFt
kh97cktsx3fo803SMcmAu7slj4JLCcVMHYYWdrpDESFcrhrISz4oPGjNjjip/Y/DLtE/x1kIGogm
gHMMBMNqDCmxwnAk/MAGbLlGvmUZL+s1wkKdeKck/5ofAfsJThbg9NMWIx/yQvRc81AWIkmmGypd
+307s09hDn7O08msdRCR51ZJrXCh6Th+K/q//JbW3Ui0kEEpE7EYT2aqhgt/HP/Ib1WTtfXQEXlt
MLSIAJROiGblY/baV4zjEEYwVtJYolRFuslZXxPoGX5grVUKIvT2axPLqXZzbIo9J4qNAoSJLfKs
6ykOrXxE348dQnWOCfiCzOnJSs/XRmTjFYnM7DhrbkofKUmoQFG7XuY8EdzdMnJ1vdrMGzb01fav
I9USYqiOqlbv0TgduURcDwaR1ATc93hDn29VQBOjdWddqi+FS2hSc1ZLTYGIPSyy1+iAjpHPK4Yh
VS3ZciZD4T46rw47IFwJP6/lUpKr260RXK1u247iHmNB20YV36Hf3CnzeFqkBLdvE/Lhmi9O9d9+
TQlDQfZOEJQCmxCzDsl1whgC0Mty220NQI6AlAQsnpJg3lNDZNA8Rmt0NAeXKQSdD8nrNFkmSz3a
dbJC8HbEBu8IpI27k6AsX8ViafB70O+Ui8YP8jxOVKHtg2fnc52N6bmTyWL00QJBFxQvdisVpdVl
+rY3tLNa1Am3YwN3MpoTUtzAN2viI7H+Nip6cGM6fgtFaoKbIzUrO/XXhN5O8O2sRsh5np4m7IQo
ZsZmFY0bhdBbx9oQovdxNEyLO6JVMURuAmeq6dxhNJriSlY0hL0HJn71cY/mpR7X1WOmseub2t/D
QqQ4LzwARNa80lNTVWoA0+Vbnjq0+yJnp+HI3KIBgnJ+++tv3PrZKTwgbrllUM+DTqoJD8S0ncWU
larZE7O1B2cqzKIOt/bz27VfVDkUYPZwJ2KdOmO6WeCvsU1exRszRHYA1KRY+FzPCS0e36fwe++K
jeNPCY/j+zeWQaxMd4d8CsYCc0Kdp7a2X0fN1nvAas+7IsSVjxJz9PM21wzh96OYzy03RdeGgIDf
qVVa0KtSN+tC63cVaN3JKNvoPwP1CxVLcIaoO3uvrSzUXJreFocGn15m+GbHg20lBkcLntLO2aLl
g7CGQd3Zy76z8jwfunghekM+L3A3Ge9UmpA5H1/ux6XRKcqFssN5SWJ9R8/VBZUhZhr1/YvCTTrg
Ly4UW3XnBBRHMahdzlnp+g7tI8rr6h47b3XPVy2M5WDM+f8g1L2+Le5BIXe5AgSRL5h83pMVfa3W
pMHq59WVw1F5uOwy+xbxdsrhrrrEppJ21Q6GnEC6FBLls4RQQUJ7IRM1DnUpHf38Bi02IWTkEOSO
bgfle1QUBg6DNL0z2IeUgrxr3dP0V8wCR0c/By/mYz8LqdZixaB4Nqd8xp2JnNsJWmTO1vjvZTId
Bft4Hjzddo5zfQFIHCzizewQuDayFl2OhNas69G5NLIPG5tDyabEHcsA9fW5Ctxtgm16iJFrUTAI
dxWb39U+GtBpjOryDXmln/dVTGrGkJcVF3aTe2nzkJR4utdFIyuU53gzpU8rHyCT59OvOTOch/+o
7XXRFkY1f2Tqq5w+djxnEN1v/Tkax0CLGYy8mH9gVnKEQO/f4udrIu9EZo/4bKAcGBFjyhYocBoE
hxnP8Bl6mEeAuCl+dFISEJQ8B40BN300p0YQnZZ0BdZN9LtCxkm6YbAqXiFTs68A6JP8v7cZ8dqm
5r1LBIZE/Z2J9PoeyJGIRL5RGK1Qcp+zyrYgtnVf3gkVHD2Dad1Bg+Gn3kzfmUCY49bz87/LGGAw
nXpsOiqacShBtLLUaPO0fLGU4lAkWm84gboYP7zoetpYACD+EuU9wnfve+Zzj8FGKAIXY5bgLs04
AEQeaZLhnQeLafntWeLjhYPnSmPkZl+ePzXMh0pP9iHMGpzvmp9Byy/xeGL+xqPS1SwwetnUOB8C
8xnKkWLPYgXYExZ3FStoRM2MU/BJibBtuAtA5y0f4acr+ABt/WzV06Ex0toE+yQOWtu8MbgCRskk
KrcTknC3rTAoQWXLb0eYWhyApEHg8dgI00wevpf/YRxGd9yL06swVZsg/ybqlWdhif+fNMV1R2f1
92c+R45pZnoACHcdEm6yZIVtuKUoLMWT8Pn4YZrEwVOSuYBLChuj1FZ8dR1eir6mEm0OVDFRwsm+
0RPZwqpYQRu8delwp+MfwtaFE6yTnqQdGGyVeNyXYx6y7NK9fLB+N+yOI3fP+5icNwJvVOVjQumq
OyUvmmHUktb9EOEbw/VimPy51fcjR76oBM1j6cPSfqb18AFA30LFO7zpd5acZdenUHzysYHWu6lb
xHEoKJIOBOvxw3zO9T6r/EnUsUAVWYvCwon1cxdvUIaieH5DGfb4zl/v8QbZRiZjy730HtKqrBcU
6MrAku8NnA6LgrvRrzQS59uCrLiZ7Lf1Z1Zpww1aUHFPOkPBG1GJKP5OshzB+GQwUOR5PjvaC3zW
uaLxanAGSXLUQJOL0TQO1kVNN+9GzxLmSadLeG7njxATf8AF3KRmAnsAGaYl6PmNtNK5ccLnL8sl
IAEKPCJKrZ/TI2vj1UZj0/VCu5SgWs5JHWIk3yjooEcTsWIW3bXjYf4NjQ+Qa1ZBqU1CGf3K/rKV
PAstz3QkFZiu7rh5RLkA6F9QfRx3t3JhjD9J9UTseiOCjYKalb2M9EVm5a2aTpGczdjc2py9Wlyt
EtiXKaRNSAtoYR91Qa5YBCPHhxzUHBRtqfP6KOmFiE3mNcyln8zfUCCK2/AWqW9cMRZrsyF9SW4p
CiL0NZbO3E/Sy1KYCHXjFzJ53ufrU4F1tZDZy+VoB3+XRx6bDDDQOeAv91O9ZU/u7NN1VGMt7t7H
u9OFULPymQm1xjan5lxVXsy/DqBzuCHCMinysGRchYekFKJPTNLbn7X6GUUurvyjIyC6aC+PVfeE
ZkRVEegE2Ie8R1dbx+slnn2F1mbC+g3GTxUTFLUxDbLcPfNT2hwKgH+V4n93JTaLhlD66cEMOtuM
SJCmBSycgMlWl5d3e68x09JecXrae/0cad+6Pg2AOKZ0opzc5CU1Z1IM09YPAXs9UeIYq4rVTfVJ
OzqRyLRWlHhj3ba4HQ671Lv/kuVYgKtzC3lYsPzZH78uUHq21Zi3TSspAZVbl6FTrwPkqCVE04Ld
KP30MX67wmHmnUyzBdhP5mpKQkLMUWSGe9JE7Qf1OAbDYzmh/xpijPFbI+Rh3X0jT3T4XjT3QuT5
aEtf3OkVK2+hMCbgqM//ommagJ1pWSMiC9n067jYUcUbA961GxMVP1QSuMIYMvy1gIyh48r6LVOx
lF4Btidg4R5n2kjYBEMONdYSPUV0Co4esaBqcsoyZ6UbnhJD01rzQqfgrLkmpFnNGHA/tepm0Msr
xqmckZ8Dv2rNRHHn4FoJ0v+yGaEY8VGSs4UzNz9EVsAFrlvtN82+9FUNDM9NJHp/M3NI538z6BIs
28lc9uHpzFx/zEeZzd0BsZo/YUqp5Q3HJkq3xziimO+MEa8xhF38yDTAunt1OKKXHVQz/Wiqkv8P
y9vUL87kg9u12ETfoI/a3FrT+hth+Z4ieB4+eBFQZNXcpGDyWquhJIboegvq+d8QNyKE05ekHF2i
2vVd5Dn5fb1IHZwia1djiZetASHJeoeUzI+o9h9ecPWZLylk76gmP/KT2uXkDEyZzzUlDjsho+d1
fn8rVuK0GzQ4HCJPcA6DsYpjJ4d5WDROKy0MRsPY2kCDVtTNFqaZawy9iz8GiCagMXymV2qb4H1l
AF+GKzr7n4L0zMz6KoHKW46nJhR2B69Zte8z8/Xvg2N+01kDXVUizA7kNl3pWYZW3yTSB2MYA4Ri
1jf4kk4Ideu6jjkICVxKnR/PdIDxDUL1ZzLnDqRjCfVPktuJwewtKohZC7aWuCQP0N18v+Lcrfoa
JVVjyELwe6FtbwlVaBDyqtir0DFWDsCvokhwrfDwU76R+gnMnlOEBS1DNzN6m4UFN8N1W1SbKYqJ
4GAxzIXwzir21XZEN3VK+HArZO/iHPoYLvtEP5A4rk/KYHNBN+ngC0gYPEqL6/DOgX4ycO4+ZHHL
1RUqsdndtlOtTbHvHXrWWVibngeAqv6iZe4YmqTYAD8dBjYFfi5VLyXNk4FWe6EsQOfKHWTagVY8
iwzmXAJ61PDaj9VPgD+N8/N/kGJuKjPtV51oiKg0XYsU6TUgGXPswMiKZXU2yIwxn1phDjNDZFMh
L4CS6zXOPD9xK05DFO6GDLCAolLZeIqoEbh/IhEVZbqf3+zkiXoRM7vHhcpH5law7F1eafnnawo0
dJAXtfglcjKlEt7NVQtWBD9o5dQlt8+RGg/0VpRB/7wpQviX4PRw63ZsqoeViJU9PDsh3zUvhBJe
8cj8qDeis4Ymgt/+j57w4kmO+4fm9qru80HAP4+k0cGIwyNyOBJ/w7dJgSR/2ORJ/my77w1doJF5
Is/H9R92naijgav325g8LCTXj5th+zO2SvNC61p+BRMQJgwaVzB3b2mIpZqW6z3T0GTkalwfCLeq
lWnwMlH98tynSa+oczeWA7vwM3CyX018elync2Yidt10jujy+bphwsl8kg05HWQDELvUVWWW7lox
0M9wVaFpt7JO4+1ncgIfUSEwkVMTchJ1uaKylND4v1gJ0I4eB5nEn8C1pUphtNoPcV5EoFlhoch2
8Ygglw8TX5jXwWwocYWK0Uf7MQeZVGkAWMn43JgOSeWSe95kfQRHhtJ2ScrAMxa86b0RhJOCIYTZ
TpeETgeK/ntgDZ8DzLcQgVNbR27MxLFFp3IWSAd9bWaa/S/Dp/3Q8C/kfOPNYIaJKb68ln1n8sO6
yRy/qpzBnyfGemAQRY4xxfuBY3cXEG8J7lYwFXa6eRRNMelD75uICa1kTLAmHeKGGiIR8cizxT4n
iR1JzpV5ZAtb5gXqwRSri4Y6iq7NmMwPr5jFY8qBDj6aeAadDGrfY/DxWKbLniv6THKehtjvxu41
0JRwaLMD0RZwuTmVRJ4PUsERP7HyXpz9bEsIhvQ0fTYlK68IH0J7uRJRtQ7GdxME/utVTI6GFLBD
c1P9JdObUuIqZr9yYawY6oFDKXoIkv5b6IwYMZXOy9n6Ab9OmvLrmFE9fSj7yTGOvBvN/0CUEfod
n2RdWSRlH19p8xiuUGd/nh6HczFEB6dXgzlCE81WPRXzpiti3m0DSYSAOg32zyM/mdiMRkpodQD9
D3bwfcjL1tvfn2g19mxJsOKg16ADWKUSyYrRV58x6WZpC33n18aivBY+Ltp85rRKp7TtUjQfQDaI
fUDvdLU6R70iGJojoE96UyC02QZ3PfwhwathQFHo4Kbxagmp19la0nXftwfRtgI7TU4pU0/APPoK
5ooMP/V7AUMr+JZJLv4K0T3g+rjCE/DNcl+8UfSk3r5maNGzrO3l5uHi4wM6icp1gxGXVgErIGH7
nMi/M9ozvDT/eTU82QRHz67qoWZoCBSswICpP/0cKP2Rzfvz27EJWvFGeC/SAcJUql6wYFKsOJxD
XVWa7/Vd8FrMyj7/jut7KiNkzY2+lRu5BpbVdko+l+Ls2MjshLco6rILSTwhDfbowZA9MxgsFt+7
sopapn0QgQM0iYtY6NXka/SVRgvSUpA97TjE6gR2V2aVXRsEWLnBHNNpLf0DPPQweTvLL/caPGAX
gPWsbWraDFFMvYxqkMqJGnvb/u/nJbdIzprvBcBTv0/XaEUkUyooe3eT33v76EsEhtAuEXPlmYTY
iInXaiZtDoQtz1ws+eigKlFUJAqKlPqVF4Sk876SnD58t1k6FY+AGkSGCzurPfyY6qy0zay/bWRX
K6+LG5fg1JnNz9jTynTp+6wjlzXLQI6EOsI3tUMzxegQf9akaOtWKHIn2Cm2JbS3wNlyD3hQv6b8
pnm26o2RhuUS0k8HH+ybfvV84htnFMcKe/QvD/jGlOBv8x0Iin97e1YmDos7WLkQHMHBo9GSo/Ov
OIUZ4/I2bgBuaQCxxt41qSf/u1JvouULUzof3H40+PelXnl5pDHeZuwMuvqlQD98vta80wslON+j
yW+NQo9fB9xi/b16HnSsvq2yZrx3ffeKLCy+0e2+bmD2AlI/WUWEFo0kJ3o74bgCk1ssEwhDGvCc
aaZY3oV/PyCE1R7469ab5TGG/EumJrjKUgddapFhpS3HFWhrkYcayCeLR6k+Zp+JGPoxRpFPJzQ4
XEr68llPV9B6oOktTAWIQyt6Nrb3D7S9J/EHEWBYJSWrCGzrwQQ6akWPbZq/TVxFsvEVnz23jqVq
2aFJ+kS3EkPmnfHPJ5mhFzVZPt5W/9UCsqO3ZtdGZCXW66aEy9Vxxl66ftO4XcX9LQ39r16HwVfH
rrozk4je96OCkLOjq1A15mwth6DdpgNSG/9SuJHQhWltlyvW6bGqKUMT0WXoPyvLY6mAp/+VJQV2
O5ZOlnqYb1aZFls2f3RGIDdpX4SGaVNc3DG90OuePMJscx1ucBl7Qf0Y+toWNXpvZZaJhlUyPFyS
w9ki1ZMmkYSYGgy1I7KnMWP9PCgy9MJU93qfI+1mUTohIRD2ZcFxabvLJmbxt//9+R6p1oyUZRUF
N94O1fbrtB9+Ub4Q/mVG4H21RAOv85tZ5hwdQHYWCW5AIeVS5zE+C9LlecQVxME1rTqtk2FrT/Cw
2HCC0s0PPcvOUFE4mAbe/jlP53KBUyFXd+cXL1pVSdE3EzK9MK1uYvY96Sy+sDJtjX38OpHiOkPJ
cvRxVR/GrVuwECw9MnGrYnOuXPl99gfd0fYUx7prURX+NnvWQ9FLcQJRcxHEmkFlJUFTIO4LjXFJ
CEWcEzd7jrYx+5m7TkaysZsnMiCJhKmonti8PUo0XVUs5vNOR6cVoMDp2jIVH4qPkKq1a2hbsbOT
Hfgh595nfKnQXjrFDalQUjHNnWNNWONDi5/ds5ys5JFHpV2pk8rn8FqoQjnk+zjpf070QFDVO0UK
ynWC2tKuYDkDsku+vW15q5BeqxC5VpVE+lRld5ktDB4C4AA9RnIBFwoxKRRBBb3GxWw5f62EZctZ
6HDQFdNzZbeUvBlm0J1m7R3ZnJIS/rShrwxeHliQcyIhFlTz/WmZr3hz4IWjbIYJrrBy+COafXoD
u1sCcGjXTgj8QfhxeCAalRiY0hF/ggE2yzbeF4jRQ/xBUA7gp5XB8NBY8y/24QgbEjx3z5Y9cxaJ
irYPNDcTEFdTXwZaOTybnSq0x2UtnmBx0uxA7XaoKEileSvNHZXPxjnCRBcvrvvZmzdKi6HuxVc5
P2APHnCUd00Eqbbgy7kLZMGsWdP0MYeMAqPVpYrNllrPaMU/uYZ9sL1WHY7rswMYnkK91BnqYagd
BvwfuLVF+gtmRcF3DqDYsS2zJDh6pSq+g82tsk1erF2FO1Wgx8FDJtRfZTT1AabQMySOpdRnAEg5
0pcSsCn/BMIrLUyqLYA8xha41MEmTyUloZjPS3nLBFpIzxZUga8nX8dH4VIFGoyIhvg4lG0FUvBB
bXwOlFBsg53PKfs7XhtulYCj3vwdkuyXGjPs1l5IKctIz31FCPS9KBQOFKov40cc4yDr9blfKG7v
K9bzAYrLl+pcwK+6+EALYjKcFJl72PuhcfnxKTFF+o2CMry/+mwnl56RyAE/iZqG2UxCQXXs75w1
e5ihrNFWSeMoQjxXgXgdV9nZUndY6rQLNSAtr6gae8/KjlfHkdKfc6YkkkmTxrD0l1iD22E5tTik
S7FFHbJ3KNZBJiZ2yXMsgPOGLn00twZWYMcvkneygpOOMI2nM62luxCEmpsW7wPv99O0+BE0+Pz3
wOYm3JI3e6YByi7BcXwSDf+POCZ469YBs0r6c46Enjo+MX98f7h7bavW2vnJfURM41oO7D4GuU3j
6N3fOCDhkA4x7KTDbCAlUDuDLu+zCmKxpwdlpyozLiGLLoONgx2uvvmU71d63sxAI0XGmOYlqm+i
ygY7YAaqfors5hkUIITtKVzZh+dOJFBcgzwwn14Thfq4ZxpLIPLTr5jbXWy4Vz9eIaBvDbm1HVqc
BvGGhbAQkN2WXkXNC0EcPmz9ZQTjx2cz042oQ5NMt/TWsFGpDMzYW8v9rJuA1879zHCDAkoaBCBd
VwdrAKwpzibURxb8nUklAB8MXqIu1IZ8zaRB8tSN80Lk+kWoSc50mXX9pflhV2y/E7nJtFkFcZeW
93P0Pl55oXz5hf1Sbmt2aXdrOdb/KRmipV+ggocoQAPEGWwYCFrCtpNXUiDW+cyG91UTH6ddAZgi
b3IJwCWzFLHVzZKBF/Vrsq69J+VcGT4ZtAv8ODX0US/P1nkZaHsvwRtZq/xFb0A6mmR+exQYBUe0
ik9L0JH2hSduZdB109twhAAcdJ9sVfYubyT3FwhN4rMrfjKLM47ExkootWCiAoK6VN8VGdi3kSzT
vibRiSMIplfczW/OqIrl2AkM+1V3ncZmjISIj8MwBqFRR53CUVzL9Y4BWIfd+WgfZWwSeIeafzRm
11X1DCXvUfBkxWoq/1mol681Tbd90jt+9LjAZZUDG4GH2997ijmMX5EdLvseYQgKxjF82VuiAhXA
J7oT5SLkzCged22530lHZTFku2sKYCC9uwLBSJZ9yupLejfJhzhex1WwYVRzZSSgIgoPNtR2N+jH
p7YMnyoM3DS8ouode4zmidPMI/kV2a5ZDqR7/3qbfxbN28dZUV39fOJp/rK7Io2KXaCrgknCsvvB
0vEq2oIw+e3KMb55VeSElzW9CW6Ox8hhDeCEajsxMLwzu/+LXrlhezs3W0IZk2bPYRBEQPreBO+x
MNYxmZv6r2S78osUVodlMxxj6RTHEXBcEdeIc00yUgB6l7hJb5nJTCKp6usfqSObh12tPulqcM7N
J6U+kMLYOxMj0kiJGayaoeigMmUw1xllF/dII83iUDDzDIbiZKr9wtuWIaXFkPkJpZANQZAFVoUB
td4IcnuiBwNwDyl2tFRBhuAQqzfuDiVeUkGc5j0pyB4XOiskI37eXRUcphqRr2F3bLPl7C5Raj4G
k8BPdcBS7lGxxCama8PlhaFVP2pcvuJ12EguV5Jh+J8iNmyXxr8ZkVqjVjTB/BFnK+0McPalTH17
2DKDA/3MkpZ1FPOL1ABeNyBFKRm8YDM7crdwbpcJFYXnZih09jGc8+oOpTCupNfLEQmeYhuGbUWn
8yZKvr/BMNns6zqM3lmMoCRjHplYfAppibLFDLFrXhSMjnj4iSmVX0FLfbXgsDSLx01GfC6lmZdv
31hlGRpqe02E1Fia8XoBuykeE0JYSrp6ZBXp4XlyjPLFHVjYHz3bUhRQIQdwNZM7qO7xWJLvQtTi
ZwYMWis0XTV/L0MYWsVPSF6j9XjtV+wHQ2vRec/O0cRH0+Lidpt7pvmXjR1zEJK+e0QcALCdKYMg
hkLxLLsEfqClKXjGbtXOGS28UIzzJxLAS+l9B5WEOfXyhPSU2WwBOZXqrrto/EpYyUzLoMpVQ7ik
+yoBifEmtnJjS5T52aUc7TJEy6rdyhUbwKU856MlyZ/xWqsebhqhaFOoQ0xmrcVVsXiw37twCb8x
6xDcFGfk+86WpeTmGvMaIusWROrbEBcF4/SneUDLc3778jH/jVMn+XiIh7ERNEM8WHfEMFim/mCH
ZOsmXahhADiszFqg/Uj2um++KMHYPiuhntZlTXughu5kzs1UraqMf/uuv0ab+XLY+P0A1t7Bo35F
ppXJM5S14rgSX4U4QJ8UEyEcy36fKluP9YyFuV5tdfAKlQuKVijDXdz2VeSrerux4GHp4zzSPwl7
EmTVkgXnUe68XKH06okFFisY9YcjuYYqhRrUJr0nr12AnrEIAsW+V+L4iBORjVcvyOLKknAFvJNf
Gr8jHXh0mg02lITAzAE2afVsts9XgRgCavMpMNHzOUTvwnXZUW9IPNwN33n0FlLoH0xWferWZ3ZW
Xcw9iUq65JIIvLXldsZDJCpq/1iSRz7eWA/LM2J6fobWY6ma++zth9rQq61H4728uMPwr3sSVVqN
gw/D8AgXRdfz08nVqPPj7xC9Zuy4GsSYz4WZ5Pii1S9me3l1kbrtOaUay2OzAtDZhriI0gLk1pgY
KpENYdM3RIJk6W1Ve40yZev3aZjD2TM4aJaMDgHNxTfy6Qzattc0dmY7ANSc46nMeW6DvfAu9Ohp
sqD/PXSr7yaNPQTYlueWsFunD5lK/LYbikgzFWvp361wVCCijK6qCwbH6In2hAahyrPpFE3fqovS
zL7gG0BXSCUgPHlBXavZFjL/RJfErZF57eKu3YTAKva0RK33yMPClFL88JHOuQhfp2GNlWnjurq2
eVKYT84XhGBTiIUEHrPLVZcCFHItbD3DqQu435IpG/ICYbcDtkw0LHnjjiS0NKHlsLG8W3AHUMiO
cdswAA9Ak2G29iY5WHgasXtS+OdnLIRBcmvUY7T8ydKs11W7/qDtgIvQLP6FDmoaXidVV2xfGZGY
OSh/jKIyjyhe59zHhB9T9MqkrjArHG7GX5DLxrZDioJHlP3c/zIb1prkmFvwwzqmLFgLoEVH4rok
h6V00xnkDoiOWxW1QIGg0woJrLlotlM9J9PTxL34Pj3l5tQCT2+CbCTxGrjScAITqGa7daEPomCV
6evyB7JpgxXfhwxIo9Cm57+DcRUyNY/MIQ5/Ph2U27XANrRznhEZEepOxFL2XMjM+Qh0mDmSe/FB
aKKbvHMdvyY9Y8NqP7IVJi6dPKlR7c6Ae3GJ6u4z/4Pl6FxNOlCteuwRO9ynrffk8Baqw1nMruFZ
2vMdFKOOgzenIx6PMwMBUdpWYutGG3/S1VhoHTiOIeb6MJ4qEWIOYZXK4ntcVLNOKpniT0vLfEtN
XioJmOFQ/fDQFJqHun2iCiMl7nBdQQs4q3fs4g8evB4TTtqGLF32P6SLWl2CA7d//h5/NXTcmGKR
K5+NZNUB7qLs0UDjQJWkWcBCzCWZ+8ATjCajTWTGA6BcWKmkLKAm9QotpR0qEvh5Hln9QN/h6GS5
4VhA9cz9YAWFYqVAvm1S7N03kUAF6sxVOVsT+/ZwXGYGTbpixGshnRzIdUhJz8d23OfmsuA8wTwj
lGiiOXP99YZC1FS5hRoC232QSiQcqKy5DpmoWKVc/eDazdaZfh1ZXr7u0lds8dQO9qwht4E1+7RC
qpnoofJvGcpFgL56Jo2soYWosgANGuXL8FVnGqjohXOeCkoTh2p9furhXSq0N9qxIHeln9WTpUnv
N48NXIY7ODTL+fyeH/dAWQM/4HxKdvr5eZazLfybvvQkqnUnZc9hjOpRMN/b4U+ZOz6nLdcekuzi
Mw7xi3KIQqsanbTJJFAS7zAV6fvaHt2ghv7WrwxbYXq7XV7UDm8W8EznZVKCh6aFn0hUvUR6kUrf
8k+Jzw9jLYDV3a9POpi8RjuXdr7A088qiGu7ZRMAwgATaZp60jExyXglUErMEUowTlsurBObhXwl
VfOGRG2oDYfVp/5fMNDbq9P1xtS32BGLCFNDsIWqzZeA7yMOKMjZKMLTs6ZuLD/dGZxLgolaZCAW
zdePEuShU1dNw1cSDQ7CkEv8TR6e+NannieTzaLlPgX2ET/D6gYuLXg90LXl3Rcog2iVM6K/dl4u
+bRTLDOl78iOM4/Uh/h7CwFRCSuvSG2Dz/6o7MLG+rxH+K8qZmthaCf2KInndbUjMB/u9hbS+MMk
ctARq5hHszzgjx6UqnfFtcQ04IaHqTlVhMVhZor/GMmVpb3fPNGmxkKzz8WkWn00kTR+0IYloBEU
MVuHsJ5KID9BhkOcEHTCyk4LHMPvJ/b1YaPhLkqoGmqmuJg4fPvAygjflQF5YrfA641dI2O+GaG1
v6rAys/teBqhznyZQwhD4q5LsF+LEGTFPdBpdktCFM8Li4inWNcvgH/OUalI0z+aPqa7d9A0cvzm
siXZvuH+eTv1xuub34tVNe4S+3UfzN/EJpRd+AS7XsqYoSKF3u2sZm32jGSC/PiATD0f30sSRbJF
iR4BOw+CjSrLCkCK9zeTjXBbzgwN8FAGGjVTmhTT7nRJNVeIKD8PnrH4UGBLmmNA6Y2MTQsZ7BV9
x29dvhQyHIBrjsUqYnd3K1BkahcP3B+ctB7wcqrro1/wYGA0dMD5LBXg77mND7iGhQ6WrH8JBwoi
hFiNuRK41L0+PxU9VABYo5t/NY6UmF97Eq4S4f8I7ocNcgCRjgWIIb8pExqnQVw/BzIQI/STDF1j
1cVyGFaKvDB4aoQ8LzlzWWWhBOIW6YPJs5m5GYxjBwnZNHGpNfvKVajR+z2mFBFgkTASn1TGKj96
7MMMHNc/dUQQNUUgPfG360rUIhwnVXvp9daFgEoq/j7oH+LJsPjOXXpQmavrX8jo5cZ45/J01b0L
dXNzzBxlOOZ/oTrAC+wh3ovkdtvBDqB2rkMM059cPvwhUZzcsQmQlRFnK6q/zWzlXsyM+vh3glGg
iZZp85ZEJo3FQjm15RlGkBVSTWJhlTVy1NdIMmOKESpn7jGdjYGOBjazDAWsbxOsZWhCLBfAhXsM
PCnC9gmstGupyXl+EZJH5kMCQejfjeCSjWLLovygnCdTUAw/sqVRHnqsSGAsLWiD4/1J2EoAqHF5
Checs2ZbjjHrsgQvD0zAplTMeEhwqNhpKEDrxz5lH874L1I8RV+I9DpqQPCIZmoccN8gyG4asXDb
6GA/Gaq3wWCnHeIn7aHn0qT63UDq6Lvp7OPNnqrWaA+kyOSk2SLffxgMuev5kOsd9+YmyHKn+sXG
t3eTUowWphN2zGNS55jIKpRknmGcu8hysoRkClTorjdp40cLRdcjWB9UyNVYzT8nL7YQmwaY4o4T
zaOv9fpt0ValfLo4ptaiPdguMnYtMpxddimtSJv6Xnv8eAwgIjfMxQwRqUqQR6jQ6sQ5NT8Tbvgt
ir571cOy8G23UiM0QxohQZBY9FbRLU2b9E9JT6Foh8gDSSlmbNjFO/PrIj9+L+ftcl058E2xem1d
92k6D9PQA0nIpW1XGcpkmChlf6zI2DZTP2GZNkNasODGCSvzNHnKzHPv5S8VmqighJqplqefG7xi
n1uiZ9Sq6DguOTk5RETggwEOzOAYvFCirpAOvCv69cTK4eSthzdD2wyhlRVMPR4UE6STjvdvltc5
2rzFGeZtUxV7PIj1BSqbSocYk1mnVd4pPukw00ly0eFNO5mnQJHrpdesUD/71AlDI+IRuMZrH8eT
EdXqHTfA2EMtHx9qGnOJU5rTPsr0iitemlbszy54jo/zTBww71+hkIBmKXCWEiLfoiyiOkjw7e9f
dCDEUyUEHRpDVzYJf+dAa46AuahtJpgsiDUUcgIcpsqxF+yf87b9dNZalETDCwvOoZYG/v/vn4U+
Sw9dDd4yEMXCd7WT3CFIkMe1MCH6S4+8oA6gkhIN8n2IRfNHa/nda8/6e+AVK0vT6l8xPSBU+nKz
8xLxz0XxkXvvVJa9xJIV4SkjnN4kTbX4Sptax65UpzeAbP3KCvd3+S2zGXs4RZpL0NOrM3yq8+fx
quB5Pus16JyCWcuMiedghGV2qpzDT63LmDY/kQ5J4JAxaWyGcJc0gbI6wx3WH9BIqpPODsA7E7Yl
sMbYTq3N7SLdJp0M0W1jzIB8xXAtmbJj5MB/VbPkyPPCPs7dRwO8AkNJEoJT9w4FnXbX00vBTgai
51ykERH3C5HrTtF5AqbPzQLdpRBaIjE5RviGA9UuBrQC1CifPwSBtlte9qmp6GbMBFJslfU+ZV3Y
hFvcTsKbWoKycVlgC0vaFJ4/AAD6Lzkyzwn8AwdYZFi4I34HoKtpfnVmahVJKe0glW2sMILklDCw
GHexeSFfI81/Mu+fsbwMJhdOiKb2tMXa3uc/xb2d3o86cK3pU0QLKBNjHiC7iH8avpxwaZCwW+nI
o++nerzCbmp4857ofHTGJSHwdHeg/TRSd4HApe0r4PQNfiWzrimmSC6JWysFkXbOZDP3dMdx/aDl
xADa80UUXKbykwH8hykK+hQkKyU+IDgatUUDcTw8tUEj/KorspdA/NoXcVSYM0/t8RRTxYI4TTqW
E1lv64VcZggpnr3smuz5m5/sjawwoWpRWjZKFIAFODHV1nVuiyoP1Od0vvc2nxTluQBPwP9LIGSg
aIpJ0JTwopRb4N5snu1r7Lhn16qfItc8MpU3XpKAxiyvN4KxukV8qAgAD5Afx8yTF5Cr6mkco2PG
k4fL9fu7ofPcM0LM1XBq82BarMh7naZlx1rYq1QGtf267Lo9HMT4FZo3Khc2AI2YCLZ4BIwggf08
QqHeaLl65sdmB8ZHxLTaw+zoZivf6P8F2O3iGHjfLRbOnJSauEhynAmFH22Q6R81CRX1LvS9/sVe
9m+GKxane63eg+5tyY9DRWmVW5qmvkXLt/0rmpGToFk1DPk4dG3IG9pGkPxByJXEc2l1J9mOPZwa
CkXv42gMtv0s3Mt/5749I7i7Mhl//0FurJZnqJRQJss8XteRwnxZ2m8wmbLgooxu2LqMsIFES7au
xPunNRL7GH60+rbNH1ycQiAquGUZG/I75nP1SZIKyWhOnQpN/mzKazrGD2HI665OvvdjVT8Qei/9
G5TIg72GWPqsPnP/BrMaPQYq/Jq+/QMTTSHpU6ZlB9LJeI+w/VjG31EDryFj3mRaCLhJpurDYXS1
sJzQpSCwFlLHMZQB31XvLm6iH39YUn+IyN+YagIQaRvwql3yIKnmTkZWr0DEX+fVr46/3gMZ0yo3
8d4nN3spCSGU7hOiN+gO8jc17U9NUMsuKbSxOV4tC7SZvfNrH6ZE5SThC3AJi+CaTgi/gElu1IzA
gqHjQCAb4x2tfrgt6QplR12xRdok5NuckMpQOkLabtO/4hGitjc/uS9oVu6eO1ALX9dkCIcHiSzv
divrwYdtPWywV2aLvjeUt2O8ZGB/fyI1ziJMZZLuKoXy+xPGqHEwx+Uu2ouRJAGv2PGrMajCo85I
PJpgigs3n6hCFnSVjzHStuhhWKymxM8fXntR8Z7yn3wXqdYKjwbDRyH6b1YesQTPtzGUGN+zJ4MA
3IWV58O9+AN9Dv9j+LLWmbD/kv87IMRiw6BxrO9K6jhqdAt3xIWOKmCDsT2G3u0f3OPXVMKLTkyn
mrVPobLo1PPFZvsOVSYnVyz5JBe49+WWJKAUpbYJQiD44rJXN8SFKQy8JD3H4eFWBwSzUtF4WhRv
G04tSjSie/OxDKv8cKOyJ07UF7bxaib2bxkWVSYbE6KyUS7MdK4BYDjaT3/UIJ0klZ87NtEFHbqY
aEPj1ycNg/OUlCZlw8urQyzodZyR+36vdJh2JED7/iBjg6sjXj323R3IYQQtX6NiHtDlAkwRmAvX
E/Eh977vdpn9i/Dow/jJhCum5nqdU9ZwO+zn7RHSDoLwJwqwxjo0CJdzP1aR0oOtCkIG3B85MFvi
//fiMs3MRUeqS5PsopOK3w8LL9bFxt1jH2rOeImS7oeeA2q1IcRt7HLtZ2cXHB4mySvqPAoskcSK
DFYrXLkWcNQecXhmFtN7J0I7KYGKjtgmb5MLqC/bvGPyxauvn2+Ul1ioN9/rUqXD2cg6AHMpdUQF
B3GyxEoMTA7zjy3tXN9iZxiex4aHyGBtYAG32Coqh5I3IRVoPMON99ddpNQaGB8t3pMt2isD76tt
L8bKTafnSjNWXgxvHPJ/zXCTgZ6T3vkrvV4jCjbiJQ4kEI0bufZ7fVCkzS6Sv3wZFzbyCHMZZruN
mCwyC6mqUk+ir30BiUi8FFRwP1K+ootKS6Ppgdql80rAVBYhOqYNrux8K14mKFuN44gG+zYZ6fPz
GUbPVJmTBETn+MyyJeyECVNcurouoGCTo5B/i29xGPdyKjTH6fEZE89nTYn0WYe42aAKZIZS24RN
sXJ1n66/7O4/vw6/zOJQCJs9qzR3PUHvrvY3RGOB/9MTYPtKQA/7YrDEN5FBXm7SQUNgOR8ROGV3
aiLuhjRcyQN0/AvOx6I1EQhuEv4Ft0AcRagRbdqp21qnbLcDiFRlLnqGYsKPKaVNhUKYQ81SPJaq
14G0Y5r0yxyc7293drwQHv8fO9umyeiJunQcDlC608/Q5ebTlDQuoxTHj1egFNnms54rv3g3T2Tx
ADrVdOrwfqpU5bG307k8MTKYuQG8zObjuZcZQc2vTPagKYZ/0ZcsGBediVvWp3JbEv8wQjC7fZVH
9Ic7IcI+FIPTfPTNOc8fr6+kv7gf6/+SUkUFUtGqZnmZSeH/dhG57TEF5AqVFmkCzSzTYkIREfDg
0BosaBgn0kD9+GJonumBLK89634hIYH1SN0W33wW9PoRBUPssQlGpJo+Qxxm2bEUulUOjDHG+l8E
fEOC3wKqmqMW7sGKyrkAuxYRTw4J47/5GzHZPKHYNIegNYYnvLhjh/HFIA0Y5nJIwCBlGZLJZ6Eq
+UmTlQQWRJCB+QJ222cb4PuafsZ/4Jkm+5B4XtqEkwcNMB+vueI2UVtDo0IMDs+2H6FgRfY41JMO
oK+pJRc21flskLl93QeKufEhwD/eouvhlwFlYoiC3C+hERrT+LmbVqUl/KpNUayavSp7L+XFxFmz
51vJFLtwAIsn/npvDa0lSwTSGh3QRsEnCOm5wGPVCbSNaXo56d2oCe1qu+ky35HdGoY6cMu2izIp
8cP4xjnvgRqGcKJ9/hOHfda25QTYjnba6wLPv4IJVXodIDPgl7aJzNggZiIhEI+A12OSIElE0a9M
gZ/hRj5sPWdgj1B75vaeSSrsx7OkL71JWqWT8LW/jybXYOl0+DvuzAJdV6DRZVNRF+ak75p4s+71
IPx/pOfdjsJDJGLwjZA4zdV/UCbKKUJHdPGK7ENXwDRJXVvr9C61JzWla+KXOlNOtqZYzHOnBdmu
uFd4brkphYj34IXyt/ESLe1K9NQcu+ViE/dNgoc0WWYJmbXw+P75I5Kf6PDhgJBEsj+IkEeGjE34
D6Ik20vWZxHNWtnOc7JHwEzU3F05Q/0+q1WBfiDplCG85Fy/OoZCcqCVsA2029ZMJB2aPU6thjlZ
5gMrKA8OWrGLnUemWQxDZNjg8GR0sGjR7yO9OF/eoiDn7uRDQCECcuTkZwKrexdZT41nVrV04AsM
2Sp6ut/ueXvtK/N5kwc8rzquYU7iL28jKD/JOkC+IFBXiYObQV6ZmmWXjg9fAgoR7DyWy4d0/dNu
LsY68SJnvLIKZIlvuXZDT8QQAU7BPMz6gSsVcucHYU61FRRFt9rm48EVOjaw+GDw8sQNrs6eJHCA
3MojNjpdHhCaxqu/rBZkd+fNFwAdFZZsC/oAjNr5ljq7qFNkI161ZuPMmd5yJBg8rM9zlnFwB/dQ
ZwvyM4eL+14YW/oQxjOE9/cRG+UJYpQdlNkc/kWD/dIlHpD4uS125wUD2Z2qZiIFTIEmAnkXu5+r
cVyT2PhFeRLgAlzapUkLfJA41Hsof58Iz+JtVdZTOgNHxFJLGZx4JgWBPWVIrrMdyaZFXPLE2cTF
ulME3VBmDkGGvyu1KmkI9XSUCF1+3QS03/2GBAN75RlrUNSSh7kw3gWQ5KzENa5+Hx7FedywFCKL
3YB/O83v0BM0I2fiI4dzB3j/+tHwdQcAReE4qmRCWR3SocXnhMv1whJnL0+xAY1q+qigJmpoD54T
NLU0j5nU/7wXmiQ0hv/NlkBccdOYOHACClZ3ZUn+GI5hOQYZwu3l+7AppWVq7WBsopLYSFoNUKuq
UpytGi+KnLCnxaFSYDv3sQKdqIGXzP85Mh6uBTGYvpARMj/T0AzRbZamXtZEdYTKH7sBZXUsn4Py
8kN25w60CsCOu1nIG/FvGwp1dpMXVVvYRC0AIl7MGkgbKKGw57uTNa/x0wvA/60N0yWwtO2ZFLi5
CYGeapyHPeV1Irrg+rqY3JMNIJ6QtBoZsYWp8P0m9MqObKU3OIeRgYYdY0l3eCDHW3yQub0NVQ42
XAwx83va6yttMQLhxDSGF9QQnD+CfrOLtJyzQVDCXk77WldFyauoe3Bba+MBIVprxAe/By1FJd0r
pzS8laLaixyJErsU00Kt6pNRkQVuDNhryr4ypEDwvpAUCqouemPNEdN+43fGJVT5R/usHKClHL2V
kf4NQQBfelxCTqVDsaWlSytbroKNyZOf/7JukyIMW8GhrFz2lrxkduRiWOM7MJWYso3z8g5Ly1zj
bwTdFAEdIpRpTWcs2cKBYHKV6DhIubUoWRS4trIk1ool9LljrdIBwj8AKHTSWCJ0J2UokszV8u3u
hijQ0kDJf1cyWj/SadkwvoBrb1l57D0xYmMD6QkHoWhw/gVvq3WMA3F79IpK7kOjNJ9IVUQIQdAO
HBtOQdWO+MwhCg5TxMxxmfRgC9sphjItqfbztqGS8ZvWg1Yy7WeF7DhjADevpuAEY55BZBNix/s5
DJejOajpOUb2xqgjxQM4JjrZBz89C/9OpMWxwmGP0paJZk/x4d+kIgcA2mRT1eZ9AQdja1tQ6nGO
UfxYM5q8PSKnKpcaS+dHyIdGfD2ZYzMOEhJ+M+xxWfxgIxY4ajKdwoIgX3LvGIP5pUFuPNiEd3SY
2CR67xORt3PmompOMLWWcabdh7Lp6b6uLO1r3GSXEjfiBxmvige4Vk0JrM9Cx3dZAhHFFKv8RTw4
kIKxQtWBXxzujXrPUwwKQKwTDlkyRqlLRfklJ5y+Bl8smGYOf23kq6unOmqZvvIAU92Jyk452gL0
vTnetkWGrDSfuTXxNNn+XA6DayhBwClXTZVsLYUdC2YvbvInmlyCilguRQkIEUgogyfoRzp50KEQ
GVQWFO2+lQ+vknECAIUmJfRuQE6Gz72LI7a7VBWrNowXGiIjy2Wag7lM5hNhAn/arZVMLBYHqhov
AAhD7e/bIcY8k9WG/XUUzS0N0TDEoewUI5sj1lGqMbkqPto1u8qiMvSzXMIFnSDKPfO537aee+TE
2vj34iVCEDFEpkd3jqts96HY2hfGvbP3CcrtynqTjKaX5Hkli2yJctv2LL/5m9d9cCRrCQ5cAWWT
P53rSosXNMpjVvA8QlaCSC5ManotN8tQUKZ4Bfim0O/t0KLSnbgU15W1E1YLqvXnu0C6GzNRbAIJ
lEerDC2Cx+Hk7GDJdp8L8kKzEi/U69dBEgQN5b9dz9y+Mjvy/6aNytuoSPcFg5r7updq1L8VMHrV
nQnLMiTj1SgG2q71NQmhWIaINWp4ZezW/5fu3HCdO+FrNzVAmTlJx/6FvVoqDWyALHweG54PO48G
btRQtoRLpf3Y0Kg5fw93OwloEGwslWQUwrDWyZ9LzZQzlbz5W+eC/W/L9LCX6zjPsxkLaRUV9ug4
ZdB8DLAPJC1HzqDFgxFrUKaYvw6NLX/uLh/Pvi7q8Ov8zjcYCZzCF8bp+5naENrA8+DgLHMVP4Or
iGqMZA9r4ikh/kGx42hwYa+TlwRPlCQiYXjGAN5wUHgguAz3Ay8KSuf8Jjq7skl1D0cWEOMdu5hF
jeBNEo9OS20JMu9a4rEhE6IiH5HnR2SGBLUnssBhoCOuHiwZ+QJqOPLdwu1PQlk4J9tilOA3bToC
xV9IiZNSnj7ScMLNHsGIcdIyrCRCC6QvwETMq/Y7x2ww2D767L/rN/JvWmxXDlqJx1//GSrBVk/y
5f8ZwY2isvd046NFlvQM+awh55OwQDvx654fUbi7QNWoIfs1J3X+VjCvfSI3coXmNc66tJK3FX6O
h9VCSVTkLrDxvi3GrwDkVHUQxD74PTj20l1ePTJLWcIqLyqEvvb1birgO34A3TU5AQ0yGO0Mn6sm
frRD8BD6A5YoTw8Uuj5r9PMUFjNhstW1ga9A1kGL4nPQ3adOpbWgGznMbPuuocgoXNxoEO/S0orS
X2m3R6B24YecI871WcTzI9HSNjr6+F+BZYroE1WBDtW1LrTMfM1KDMk81PYiuKT80e4cIahkWioW
B3vC6NtxLggFaaIOl66z7TE8m91UvEbTAth2D385KwwvYGTELwYCSqZZRAMiNlUoKYg/vie8fIi/
+qiXI6vyU75uKtdIlLaZnuc0gcpzmup6MKEppXOpk1E23CLsfqR1f/4d/69dQUk8beJpD4BBuvYU
WxiGq5MEVDQMZ3pf4qvkFTpPRRJXS0Q9BCRYq0BpxCYeYm5JJWtSUnwVJPVGVOspvu72VY39K+No
rHv/JwFHoC0imgZA1SL1X10XQM7erMnQwkA+rFypTKpBYmK1vmo3ZAEChppkoQ7bj1qworvidkcD
x68aBma4T8cVpzdJEziGKuIRPhOg5svebLUDt/cfU7Hzbr4aRSY/rbKXxsi3DJIm1CK/dZ3SJcKd
/SHVXdn2Uml03fd9kvDRQPMUhC9ZRgkjO8SnAc337PrZXJukXi+DDnakOpNSC2hYF+ak/yzq9ayL
KK6C7iUr5/EOVEUNHUkBrhELH7aMCdYRHSRa44KemZv6JXMqOYc3xjMCqeH4F01KPFNhTJ67+0ui
JXcPOGBWYjXF3xP4W5k9lSJnGXYrEly8kWuKG4Puse0kEYc4Bmku5mYzEgvw9jgjzj9MgQmkT6fi
UgWd5kh/7uNe+19bG+tbLLpxf59CMkvKghbYHiECuRNugDF6w2jJA2FxmFgHSyXCbKdFkXdezekf
+AD9ZZnhNVlJAMcyltZusEeZbZCfTA9F5m8XqYfNNMeo3WL7tupJhu7cVE4WuaUKaVKnYcDLNmPb
wzBU7/VKkSli88SEtH48UJHCGQSg2fOCxM1W4jviG1czXjOqLursrxkRlDwAbZNkA9S+vFM2GMRg
p4szo3gX28bQc/VMduodPh/zd2Q7eHKdFovs/qjIHuBwKAALjoycFRXRPPPJteaTq0+bgW0XQk3M
vHo3owTCmExmfFAJOaornVJoF1x0rwIZyVP7nD4M4ShLD6GrmfqcjGGEW/hrOFYUUW1BGwI7T/9i
laxkR466SBbJH6uUG+DU4noi/t7O/gdDtqXun1qLOvD9KIa8knVYI0RCGJ3zFuwB73WOr9QeazY5
c84rMe7m/SFa5EIBDDC6MZmEXQAWkyVVaUymiNttRDAFKthLwpxJq0owtUM+k1S6KqjaTfz/YnK7
myKDCzeh97JB8o98i4KF7+qkGrDcnoEk6+unYpybmYLME9Tx445A1sPAKE9xElpmxg30oTzoOYHD
/4Ssm0PaQ3ArHIn+Q+l25H+D8UsSvfwx6yk6Hrc0wO3QHlMmLJxFRjXYW+Xx07ORGA88b9tjBA/i
Yetpen3KYU0JMWEHTE0b1eaWY7RhMfX7b6jDxSA2ZKkjldEZmtA62Jz4n02MeNkXvagPwrvyRthD
BYEilaFp9rX2OrvmdnVBI6Dvfpd7QAGrl6XOZ2q7IwZ+nOwfxKWJZdtDfaENqYywdIDgL5PT6CIn
vDuvf0zc+CGHiR9Xyjz0i2rO4YhmtWHUCuvmzEluCESAJgybH8inXTlUhDMtI4L3ya/MrzZFPf36
781Ppaj78piwjz2bANIMR7g0UWX674gQbeDmKJBp7qrZR7oz2Zjve79wwKe7h7+GwRsTQfniRbpG
BrNpK1tOHWvPvGy5Xhi8zT2CdQqmDehZGLCT6u0GzSsoFn/6W4zugeJY6Qwp5WwYwSM8v1QgF9sW
69sIgChPbNln53dKldzDDErIbLi5zIHljPkl2WCEhGFG8QhfGu8fDDI0P4lbkRziWNIIm0dbCsFP
+CQaXFzWLSGkh5YKUZlncJNHA0N/WTGK3K4nBMcOd+K1cWGYBRozGr5KIZBQ/ncB15JOzJcEXenN
OY/pwiyVKdnk/iYewXcOGdDHDxYnuB0WmR1LmwMB/5Nh7BWe7j7d6qErGa8vvW8qTJwBVZhoF9GJ
KDf4G+abm6pDXfKnhkTukpbYz14TLTeaeNPmy7ckOD8F/U3R/53WG6yfTdvqRhALZz2DIJu0hs7f
YwyVY+ImG1ugDTsc9lxAoYDKDX9Lg0LGRiAej6YDV9B1EuxQUVN06GAZWG9UbacwffdnLdcHY4Zs
xVps6NBMeJzTUiGxXCLEvuQoMs6r0wDX3Fnv5BkYTtO1t/MhuSaOtLAEB3Yx7eha2LQVTrO8SlWP
QlBy29zk0grOGHnaQj5BLcZATop0865wxx/cc5jasRcvdLCtQGRhpog/2Ff/gy1TalEMZIIqMNwN
AQOG/Jkr0g9X1fRQhDn9EVKQXh77EjHX3oTsyRbTYPzjCDBK62hAAkIyb6OyrJPtqZRIvEvx0wX+
WioQlC1WSTdVhv8J+udOaV+mg1CiEuUUoAT3GCc9Y0nPyJOZLWjzIb7YbhFL39il9lUwwYhH453O
ygjIGAHYCEu63oDPsw8VeJwVGwtZCsTKJ448n4dQS9GFZcAaMYbhgRAE96V7SI9n2+OoUBxA+N11
fLKMoGX2kE+Z8FH9UWuRC4AGq2fXWoRChLdx0uCSCMeEjKYyLglWeGyanq/wkJS/FQ5MMSj0HIpM
i/jWRU2GN0wqBRT6uAPU+dgJ+nIYnyNZknwminY/MJRi2EtaAtBkD7QZWsCvNrsqbqvJ8Oiq04A2
nocjBNMKED3peHrYMYhFyRBEoO6Ulo8Yb8L/YlRLfhfcogbZpvfPxQ3UH16JhQjMB0hvxtwapJF1
o6LdLtC/HiLjaURBviZXxC6ZEbSUNc3+rnpMgytXZ6xfujjLPZieaWXyMBLdf6+52ObmsW/zqKbK
ElFKG3lZoeTn4mqFlxM36YvRkurJhJ+3ixzdUFDRTKA48+Bn2uBNkcElj4D0LwzNv2VpgP6X3lUx
rPfAq3ofYqG28JTUHQp3rrB3I3GirYgCm7Nv2nFkrCnbMstJinPW7bSNIEwGZ17iu5IKXOu/NH0X
7WR1fr0otTIiga54QsmG/6ns8j3mELNTIV5UZgtc1k46kHpJFEmWDtqonb/4cjuVN0d0Pm5xAeG3
5bfzF6u90ZGfs2cUxXJ/iaN1YLiYsWYwm9DImhZAxY7Zd18y9URds86l87UznwDHTuf3rlCqd9on
4g4DogF5eY+Vkx8mjfZHghxMgZAiwBJboPQ6f1xhknMWbUl6RLoqpk7PqF/cBAkS3eHbKW/tnoOA
QoCLVu/X9Y7WokX2hw1xJCZGtsfWh1mu2R5D8LULthwhSPbZJhkVdFz/8Vl3z6Gw3XKCHpPg438Q
BsR3rmGoYKqidNI4SNzR6du144fnqjGu2P7UFnyhAx17OXijkrhROE5KoufJvHgucjGvF9pdGmz2
A4fRB5OBTXUhf8tJo3wbyOgQZ+lB02a0QVlB7JxA+swTQJ1+4ZI/d3hf3jG4Y4hFGRySDkwvUIPN
F4xjvaKNrJ1imv5qxbW9Pb42sm5V94zzrhjF/q5dZiO12/8y0dbDNpf40KK9gMryMlF+gP0m50N+
6u9AH9UCqUwSUdxdj6Hn5htUWST4OllXL3CoGH5OK2Jju1EkDRDuxr0q/uPTJCbapzAThGyh8W2i
odDLssa1u1CTDsYeJu65LCDhcLuri24XCFCTbw598rs3EE5q8M5IOLcMs9tg5nf8bM6PnRVCRamP
FXqvPITUBQgs7BfARKgKzrDuNoS/ztqg6ZzHRKQEZRHlsMqf0R4YzMslcRUsWo5p0IgsYfKMe98X
Bt+pwjn/OvFygUSfWCgSx+mdYJwltIFrkN1Yff8DRk6GwLYWUzPXOdOmojgtF8WiL1342eQSnlVG
Jfyy/Bl6aoygm7Diupz23UhZnOvhcTCErbPewdXziIeGEeNloPIsNdQsvO58w0n9HbiLVQlz45eh
a63IkC5LdLU9OigeODUtM+dCCDuWgTLBvqI3i8iDoFabGc9uMUhIik1c1zeB6PP+gRqsAnzuQw1o
9NVT3GFTq1ROnLVZ1pw+kx8lll7QaMJTH67uBuIYx0mKgHUYseW8w9ouQngiKueea/hFZg/QS9Hl
ywPtttjxuTCzDhha6vhNUXMFr9JBb12Sj8SjSQqRZOvQ3NKs3PnH8uI7sbfn3O4qpZsZrqbnfFWh
aNjo/pGycXaOWLRKX4mGVrYzhDn6SGNDoZEmAP9uR0095epOGkQXZZgMb2f9WVi2I9ivjINjrJAr
m1hyTdhZhUHOYHnsw4e6oq/JP6lLsIoPyFQmYQOTwXqkzjBwgEhNpnGoL71/xe8iy3BAGhoSmJEX
em1iuxb14UJhV1ADAKs5mH58CTIJhvRCOgW2ESUJfNIKmzVz8EMvKra5+MQZ5mfeoVP6zkwpiZH5
Yg5x0G+TUeBLGjGkv1w1Wyxk079/OUCyrwEa6KY9P51qzyzTxgvbIVnCnSXINgRrJDXwDFUCOlKo
o9jTvCA5nyjM3/EShCFdFwGjgSCSUCK0ui+vAoUq8U6TMA7inbk1iKNBGnzPxuHsz1OBkig+2fKO
Uej84ELXbqHUJR5fvcQePICqPYwECcD+qkNiA97WzcPiO3pWLQBWZeUQKLgl+t/3K+Kgrh4TyZqp
URZplWuX3k2Wq7VxPdEbD7nIO5lOiaqbLf8DgGi+4dWk0r/aOvVwz8N5mQRqoXPMO+pHJPn9LdHQ
K0pf3vQhgvh/qvD/0neUIjjH4U10rHcFHKVs77iu1wcNNrszTFvSjUcOqv33xVqqg8qCT+eVMsEt
ymxHIbAV2fQvTJcISXg0HaipG1IKHEFfYsSGPQ3uOyqlC7aAR3SNXAd37tLt6d90ncesHkQ3rl1d
XpIfyt5pUz4svYJH1WLXl95/Vi1WmneabbUINYpluO2hREGLTjGC4VoLqQeUO0M2G+rcaO9od1G/
BGiwW86xuanPDs9tU310I13Cd+Hgi6yaRSSsp83z8p/xnBY5qfIsKbyKYMBnfTXd/N1jn50P6O0a
43EOh+ZOoQLyXllZPqHtwGXGchk1hQD5rYNAtO8WJmCp7+PRpoO4VEJAZ6oCRnfycFzSJaRhGa3X
NKET5QjTUQeyEE0Y6EwF6d5fCvLs6c2b8/kaspixwOsrePB1W47vgF5q6pri2jyOcyu0U9ctKElX
C36QGbumo0llrWmG9Aqs0pG5ZcKkTqHTMXOAmuoREuARn5iuUqzXVgBINx0UeDN9ycetG74IHX/y
ELiAbYEF14jB8obQzaPfXpot5c+Rs9cK9P95gOAWJVABh4SjrZIfPudZOJx3RKjqm1DY6MpwKz3M
+UyT2YkS35qRO4IjPuddOpOaDdLfTaTNeEikUckzYozRie0322fZuRBctyNKfQ+ljh/+XneWjorj
Ckuif6X/GDnalkhOIP7YkbYKAagcqVsLt8ByjsIs2+O9L27YHouGF74tgQf/Ha5EzAbNpsEnI9QW
HTh28Adpqaf+PlOP77IWHO6EZkN87WerCBbxdV/XNVlR7EsKjZxR8E+aYWb+LzWWJzQr3AmYWsdA
XXyDoRDHtmTemoLFtW648SFNc958va3Fk9XmetGuLOlpahhfs+GyxBfXonAXoHGBTu0pTDfKCmv3
dqYwb4ztrP7DZpdhUZZjQ0jCMaIeF0btiRBSYf4Jo3UgYwWbmK1stsuHfEfgad3ErLi9vpQb6YFm
rCY7nPaviTT8X3Nc1RH+FkO7D/W+PuUmFlwLrQ50xVmxCn3hBWP3q3kXLbWeeNnbvnYeAyP/CSEj
sZ5uB0JteHSh+NEjpPqP+tQYcf8H9xCCKdLAxuUSBJZsdhTJftxMTZKenhz1iEL0xx61PvSm3xGe
YmoZkMn+Og0Fk6haOVgF2PZQDChygTLS8HFhul3L4p8hxCZJ1O+9O0RRm7blVdmyVn2h9vmSRkma
xSzkhLdNyqOJhV+fgnUi6RutBDysZUkWa7nYYUsju0uaZK/XqnCYCUmtiBy/HNQIJGXMV8oiN68v
LKWLWdbNuINFH2EFMUulcdz0fbz3Lc8bEQb/ZnO9XUAYrlAB3nUytvjtqLwPu+2r+7YPcy4kKAf8
RTOIrO6xBh91V4f0zHjH5UvP8DFmPRhJFMKn+atcQHLzEMYfH3DjIbXPU/dRMPsilSdFCfX3S2Ov
q/V/nen5mZ3amPU/3uQFKll3e4fHSlM8ompCuP7EHEzw64xcuNrwpiYoM95yNJ/+O693ve9D0Ue1
IM/xTiYLDluOOMRse6lh/+KWbgYF+VcZvq6YEboPd2uyTRfk6MWsCoGUZ+ao3NPgszyUshUjF74R
D7dJYlsIskLKknhYLRMk15pppr54mS/5j1RwlCA5xmQL6Q/pqy+cPgtKm/9sTUXV/MZsNm2GkzGE
bLukidoWJ12FisIo73okEh1mpknxalIpDJo35236aDLPc4Z6fI+fxFmxhm177JNlU2F8QUx7rbjo
w/CxkKQJobdKSaSHqXuAcOhV0ZTiGgykGywW9Ot9mcLdR/JZ6hlptHON0jPrBiuXC2GWLE8w6ezh
n92ryZRba8agbN1kgP3v/IOxHjBBkzV/0iQNtTmd+fHrH/DcsmrXpB4tkU9YnI3dHmKF3Af9KcfY
6RWL5RX1V16CJcAgIFovI4QvntsVHQJFABPT3UL0QAWA/xCym1LGRz/P7LyPpviuoGpBv65VjIAj
SurhjvXpQE8bzzMDBjoUK3mgv3mgQ6RXthu1xJ1ikacVv8vtw0Je2UZMIzPCByErFbgH0AyEY0q1
L8cElb6GlUQ/U3a7ojAKVIFHTBXpLyoJwdRV60qWM8aABGSw8nQHnh+q7eKiE5zkjMXMARc9N/ta
t6MqYRnz2PCsg9q/G44jMpxdrNcBErVYkrPiBUw/hoxzAYkx/Dgo7E+tvRvNMc8+j58y0GmUSQkd
1B8WS+schYOT5ZDx+1rfq7IMTERr5CEUK8d1Gvo/e9FeTsJ0HQ61/zd9D/ay9jC7enmtZlzeA/AG
RfYCgBTUU178SvC100yBtpl6lgcjoKja0cn19JkcmUa+Fz8dMKrIy5jlb2MhMDIQAnd3yUc6Br5K
lU5R/WGzz99VrAJlbe1kWp12Bocfxc6QmlsXVghtJp9cWEi+LCi/wpk9ODD+H24UHR/IiHN0kvzr
1eBIysdYvFFdkBvOLXBd4AfWLYJ0Ptmqhfa9tS7KNXHlKXeZWx12xBs/tScipzLC3jNy0oLrlDqS
QOQgRsmr57It+hT+sSfKeP2CMZURgyOLiC7lBzYw0KExNQ/ZW1VMWgoBh5pPXgULHpj1Au7IqAue
gIbevGlY2mdEUIsi3jPQGF5JFChUxgHSzxpbTLu3A3XAiXwb9Vu/tUgB2NoATYCvKp9/YtayHt9j
S7ONE9S1UEXqiTc8n/4W0+549BJESKQvxYWFI7E70O2KDM4iIXRD22KKodqbLwubbUTdXosuohnZ
snbANklHPw2aciw+2cwWw+qALwJgR4wY8Kr6Y7vtcDOXQG6lRStA6Ve9uc4hos3MZma28xfBCSSv
HcoNJCJ2JdArsM+pa65bkE9f4PgqhHxx7gWnklZkraJx+rNwBdcwYSU8kE0CZzKQCaXMHFtpCsoF
/HAxy2zY+vGs0+OqGfpP8AmrHyM2evnLE4pp0NY3Wgkam/fWOPmyCb2DKAuy0CaTDssS0PzdmVeb
2ZfWb2SKSJJxt99+Q358uoLJF8yaTebsmo0U4s1EzAkzeCgH7NjFgoUzWjvUmlEuufA+ll9ih4Lc
CSvC/nXk4yPKDiHhR5Rn9itRhj1zLyxmGrwsGzkRLAf51ghRH2TjuoEGG/U6dVaa4n8NCPAPk6IC
rvGIGyw3cYG5grFDyxCEXdgtTp+waO1j5b3e68llgWgWkRIKpcXwHgvvV6nCGtRYYDK/V668bD9k
gCk6kiu1ikNqGOr0mqNDLatc43uTjDbdLQxcDv/HHgCK0Fw/kMwHoda8BqJ+WEPK7gCODhqSnczv
Q0h+P6Q43qVgPR5MYwL9gGB7Hbqe5h44j+OTbIGbE+dl9zli0TfjryEH0UmYQQ1x8l/KuWca+gDP
6diusBp1Jh44nHgIVQjkaPpUUXW9cE8rza4v+QxD+aI6mqM91pavyIBilsgL/0biTTCnkjSnu8X7
DL8ct1vLdsSRW0Muob8f4psgjsECJG1nGyWIac+JcLnf/986BY3Ymkc8CJMqiWqqALHqrIB0/F2d
V/4C1icgAFJRO7upp1qPtEshYk8MfK59OdhUaeBle6B6+mnQ03dSF3GqogRKqrP5Q0rRO5VnlG7/
Jb7RUSvr4adAgL3XQ8GpL1ttr454BTyH4ATTRM+S7KR+PtRWhmSuSOUFGAZBLYyRpenH8ucxomfn
6kNCyBBpyBtZOl55/ZLWC9gIJ2+73sMHsgfRrg7/sds6uHntrl6HQoaXDNDuJytBvET9d6471qyE
/VPgUpj+KmHPm01hfjy+BHnTqwMzRALaJ6wEMPXV1ulYKsXxu21t0XO80G2nSJv/EPAjTeKSUo14
Ji1156fu8ak1ls62BpedO34UHpAqLJYC3dgxZ5TNA6Tw8+9Gg+NCRuBwrplWtTokKSsWjU5iYbDW
LVcHIDcy64Tks7ZufjHgIm5sxOMEjbNOIPk457Z8irE5CEkZg0HbN8vWIMZAeExARGDXs3FGU8Wd
KPAxjDMrnob25CjZA0rGqKFtqcGXJdS3pX52tCcq+htuVGHUVOOEP7iXttntgZFpzAamUAIaxtak
jmCCPC2QRfyzQ9o1mLJFd4WMk8GXeSViR4TsD6PXBevhYKWuJBIl1menii9oWnw9GPrLeq8Dyddj
i7PzhMM3tOpDLpD0fLdplvnn5k3lvC9ZNlvRqTaU28fbVOmy3yRu5bCaYsPORHHgLeq8Facldn0E
WYtMJP+xP8la/TOnzyedbrLMGufN3UxG+DNrq2GUFQG5T+wmiR6BgzVlyC5AgMdHTMEXtJZ1vfcl
JJKob+D6iF2cKNUl9/ZieEFrHXoZOAzeDUL43Coq2odAP5T4aChN9EwDIvRVN/o70gdglhEoyAtD
4s11kAnwZcYVKCXWkvIAsMaH0/aekEM06QnOkMMMlO1LbEEbfi8l3WDEZr0s/cAdNVwKl8tRhIEP
0LK5kJc2AbqF5+4iFH5LrJ5hwRPDcY5DYuxMwFGhARvlcfACqvbzjz/Ikmfj/YysDD1YKu48GcOv
sJmMtO7PPmX3c4j9SOqRAj1BfKzjut9MNx0qwNzZNl9r3EOT2LuvIIP8Aahfp1JmcBOqvyyMqXVT
gqNLd++RQWRKf1OP/onvBdXGwfhowj6vt3f+uhgExvXcFYP2uJIaHJQ4JfDQPi+JndLcLDkJwVpD
Zpk+kZ84lExa8JblVuTOpxwbZGhISA85IFZgmSi2iMZQ1V810AdqdnCvF7FqAsSLPigvVpGd/hBp
S4F36dBZtrQ6y6GmVpKGQkyuPTHsQBtX31/K459SW08vmFtDZ0ZseRBvLlruYnLKhtxaPB1NQIc0
UgY1b8HIOa7lRNAklIbnuzdHRIEgkzxhh0jnmAZBAUTNyGIpNY0Mq9vN3Lh0k7BPl+7AgkoWT4Xx
6cUq4Xuo1LPug7DvNDqNQndJkObeeWeuEBKRDHiASNnAmbYU6ogIuYG9nLBq2Jpi6dg5qJS78rKW
8NjdEOQ1RpAUya1QDs7VbTqbqb1g1FrLS53tXlx3D6EralLws4jyUY3jdC9BzO2hTAXpawS25rQE
TblcJkSUAOufAm9ejHkAS8QOfpCkNyEnBS8A3WBzY6s5F2SrNNNN/5ygi8JzyRGiC/iv0rcd2Ubm
966dcr8GokPJ7/zM14wlGF3TgwlhAAQ6ZWm5/+xwbY93zmtEKLx1HSv3sLEZBxLiBgg/IdQFXMda
WJzotnZJAAh9jjCLeP4X4+vR5qrItCLuF+yoqv6Jn91dFHuEXcjx3OkUyfWz5ZAdxhksZiulmZuF
RvWZYOXJhKuSuGa9FyuxB7+opqoC7uwLaeW1al8WTPk+mKr6tZP/afPThPnkRW343VKpgVhpOiU2
WhU+k6G9x6im0jj0b6zw4SVVmowKfT1ZD0qIgNR8uJ1bVUqHtwdwO/31fSCOG7mABjcyH9N023+H
EvF9VURPBSzcBogpbm7f6nyuFuSTCb6xt2UFla//NJYytj/lyibBAVJKhnqjUbKYzd6ykkbzC9Yi
2syiz3IU1iIUNnc5nZ76FMM2yLk/O4cqYeGRTdmtsIaEE8beHdYHvPZW5KwkUSR3FnpUh8o47HDC
tZRYydvaG6Kpk5L2XUyQoIWjdSBZU0KjlUhmmaTi6yhEYc2VgbPDc0tfevn1ITKXzxZKVzsxIJsy
M4/DM/JomfUlGig78TzMH+w66NH6nTjjGYwgWoUCIJCSz0jRKCos7rZkW/BxdkCjG1R5Kv7N0Jh+
s7/OQOoy3A88siqacOyld1/pwkeGhziBUPkM7WmOs6sNyKdbAZ719qRk2h8AqGMTUa70pWF5Zfmj
vTQKJDlkBGOBng8WUGXf2Zq82fzzHEhRYYohoG2chY7SnBetd2UIiMR7solttfehrO80RK03omUZ
M8HBbVs5hEWAgbaSQHRitTDwsN9oTcKIeBtRqfBb3CAgkyVBPwhKgAPE2IWNFye/HX0E3F42KC05
qzlG3RxDK41b1EHJ/nGLBM6hPTGP31ax2WwFQOrSQZRKWIcdkWGJvIptz+Y4/rCPUMIc1iElv4CT
w/IHxs77xVKvUyjoC/jFXLE1FmzAJ/l7kEKqJEGuWvGF16+W4VDw6FsuEvfWRGkpi/PRCQANBzHW
R4XPY/xN8O09lifQnYzv7TSA6fy0xLPFLc2aogPgK47HSwY5qhNcjiaBxgUbVoe3dvYD4SYvPHmR
nm1ZOtkHBBJ0mLnuT9dJ+3onqHUbgEdPuW52b+SKzEyV6OddIXUWveXa7UU88Jty3S3XGG5UdQL4
Flz+Fqh215F9QK4+Ed1sFv/ZaHFhlwtMkqByM7tCsoUC3DvwT5BTCQ8Z4SURy/EXVYv81pzbRoRj
+lXfIGr8ZPX1upvn7lcgj9Sares/byoUhBwcGR9dELQcn8uWkawAut6iN2eoX5jrcCX0O5AfYbCu
sQ+wA1DBbBOfX37QiOAAizoUMK2D3x0rLxc7ZuxoWb+6/OsVviJsja+dacdZjyOCsaEJSin8m4QY
9SMUJhmSZaHnPH7rZihhAqRXC4BBmbTKfx9CuWGR7kloZneBToYj0A2qJkNtrcCEiFr5YWZL7m2d
KeK3+qrdHOG75BdVkuWPVcjX60JMHLVyqanYQQ0ynAbDuG7tGvs9+CgCcXyTEkF1saAg3BKXtFYO
ndT9tBcknt4qIVghx+VsVdwC7X0m3hdkRaAUqy8nqYK4P3IqbViAcZjnqUOloe9FBVh8lzrMVOii
ea5skXFl8Hsnf2tHGqNRWUJKF+tzX66zZWLaMLW7Plb8jr6Tiei12YH6nNlS+R/15cOkhlabHxnc
RI+EsZ6M3o8oZB2gyDjHz+tJFO7atgCu/d7YlLNBE5wN3VJ/3x+P1MlXV9zn3q5q5E69T2oOt57V
hAn+pjIepgeYwBQcdp2G1U7L5YneyAyANO5aiswSx0PbZlMFMwHtgsQYEyto8dtDSm2OhpvMstGS
mqo1lNdBr+JxMe9fbf4V2QamGaEnhRIV+jiLprQQkQ8ymZsqLfnXBINBevRwG6KTGPX8hfXBfdkO
9CyvdLRYikMzhmdwUDiU+OTMPujg947Wy7wVNnbCSbZWsjm+UQEkcLQ1GgdX1/71Q2aK6DLh/U91
fqVefIoltSYEu4n+Ao+1rBVqj2XU8fcH5wWJ5Q2YLxd7b9QOrJ+6Ndu/pPFR3vrAF96yzYYBZZAi
cQVAm3X4y8JHmuByTJ1PgpG34FOuzaaJw2sYlCQW8ObGNPFgh7zlh4fHSbXqi0TCdryh09JaPBTG
gqToW9OAkr6rneYy6+V6FDvXBtn95SVEiRNO6544jOzN9EXJfH3Xc2CkzQJOwswmMjKz5qljld5b
IH1G7sp44UJt/H37JnSpmVwuTYFfjqm7Mvhe31X6XKNreeTPD+LOmlMbxNtoOr8IIGaG2PJoiwqA
ZOEs4VcJNUQrTLThItdNQY1+foDASwE2oW3n0Z/ijUQ6q05Q+b8RnBvuZeFVUhL84tiFKyXI6iC9
5GmkvB+pcSk0toaM66Qj0YfIFyhdt9B8LHcWwqLiToYzkotGcUBrnjHxMLL5CsMNqx16Kp0Pq6kb
C48vT2Jj+1aULhMoVPaEGp4EMpRrJWcdzmCLg3d460GgtK51UMlDui1IOD2f9MdPMBMBLi8eEj8D
Z/Gq19OeYYpLOpTjayAGIrdKTlRnsHSPlu9FuctVbRp50uYZtK3YG+5Tk0pE3GS7Pg1Upd2Dl/Ts
jfXpwH/EvJub1wTQuvpIwxfUvu0JiXxWwbSEwZmFyDo4H3FARbGygo5oneVtcVo4Pcxo4Ts7kiwW
0tlkyiyjaYNPoPHrSNjHYXnwhPfODbIAUfTaP4+II99id7A11c4HCsqkxBJSjznZxY4pnAkQuzM+
5chyttxFmkkCmWyz6ECBAwR+XLCcvlIdr9DdQF8Z+kO+IDHcz/iFfgiRgwNcivssEHKUxfIp57gA
bRIMS8Ph6L5m1ylidEhDHcIjn/IgEbyr6px/E2nXvWRd2FHe4mKGqey7eqtVQaR1RTxNgX8ne4Q5
aCt5BML+pYZq8SLp9beYbGcl5EvpG63+Wc37izmPQ2wmHIRmKtG0I0IpOEXd6rWR+mj0MgGvNlA5
/EkaeRl4QRQt1BgdvvEGpKrQQdOaxpdjpagOJQDq/2jpI5LN/JSfvjXNPDU2AC0yutmfIrR4Oe7K
42JiKbyItkAsazqEPuxnAhP3nE26xIurVlkhNxFG1ntwc/55sXCIgVzlnNPS7lsNRqGHveZXWZ6D
6uuEL2E8UiDSybhWutbmCRiPssQX19BSoau7nXtgcMcvY+TxCesq6qFXganzFAKCOmGYQonKRC18
LYeZw9aGBEd0KuUTkmJQTGvI55zwK5dq2LUS6i3fIj77PibcuKLfZc8P7jFI7WsJ9S+PuU9aC7Mo
l/gceluySsA6Z5vmHaN/UJcgP5Q1Tj795WeFwN6LluYIOTRPM7gwF8v5iJZDeJkRnuqIpkf+fa9Y
va+JjP8Zh2HrwlWV4kbZk+gLrVuxnYedfcsLpQatfwvuKRR/n03Xslj1xxEUa32i+LZqHU9ahNsT
zSbycJjA6diqH1OdTOc+uE1V/3gOWDlBvPjpQmVU/yN+hwD1/wwp/+O4enHAeGeo5pAmIkSsuae+
Fp9AUAwl2mctgAT0v9e1wm1rwuX/hkXg1f0XNkoDgr+KKLSYKMV9zGWdYDdjHiUuiq0cn+jnkmIl
BiNuoX+Y1eRql0axdOs62A4OelLMSyt7ZmyJV2XYu5VPyRiDXCZ4KOKySlzPz6uvUSv90ttnF3d2
kzaKmqcU+xwA9vQpSGDgK/yh7hyDxm9NVQORnTT/zD2aWQuTQal6P1x5nttpxitqURul6qXTnfYy
QsaoqG0R/RTAc/pjteISeDv9HhS3Uqn6OQn9ULRvqauwIgCqlyhaTOSAfnP8oRo3MJr36vRz0IHm
JxOm0+aguLxVLygAAf0++R636HberVJ6b7XgQFaWR1JUEpnr+puzFhNanKMfzb82A7lhSUXOPd8U
OHWp3iO4XGSV05sS5WslQlXySAhWMwd7FSCLKP0CsH60IINnC+dnS4zO2Bx6bINs1oCkEWX3rlqY
OoRWdieJ17FiDZik3aPSTYILNtsrQiiHnzE7sN9dMrPueeILxqJHp5rpJymXNsWUVWlJwr5XHy0G
68JA2ru60j1j6uKse9WlqvSVnTdmJeKDDqnTKVbPobN5ybN1Mugg673XBXNyzmVtuO0xD1Irld+7
d92Qr98hkBKVahr6BCm6EyRusGY6H+snIb6zn+rHCCU/3rqDIavPs5Crc7IunSCJYQWEGPkw8o/0
YdKj7oYTC4npW1AeXCsH/meivqv/HhaD6YalDpYamGWfaszFTNUkdro3X5WAxxpJ+mSoEVmKZUiK
x7TR0JwBMUkg3wQzLQQhxG2LmzKuhvHm0ZmUphZr9rjTj/Hw6seAQTx0lNm4F6AY5VdPwjQEAKn3
LZQ1+zbEEw6NG5NJcUcqfItjuxOJ43YKxZ96cwg+l7/L4+HHTJuxMobsu7sSJCWhFQyIk5KSBOAb
Vskd1PFAJhCd8aA6LD7NdqjYZJnFH2q6EAYS/6DZgv2NHvfReu1uZ+t8UpbwVyB+rW+4xgKjmhHS
ucIWtmVIbyvD1hAgwjizmb7pJ1rdNAI2yS8COlviDrdyM/2mbN/4XXz9cY1TJ/4L4puXhst7sH+x
5kYTiFi1HDc4cS1c3Ddv5/Y5O3iLS7Huo+QSJsZc4StplFODBZCiU0oi1KLv+1c1gt911RKYdjrh
ByVClPu34Ygr4xLJ/TgwoGVHdP+3jcZaK8kXY0QDzc8AlS3onKMuT9lsfQw1A91rjM0QNOS6ugMR
OxMhLDRMplVwh/c06b/lQ8Rex5z20yXTYVfEA+5EDw1z1YuEaRGYqXHtTcsFKEBmyLFC/DjsG0cE
7535YXaj6LGOaXJqQbLMXW3puMm6gTJzcBD2SGGaI5fE7pQ0251cQf3weRPh6U/PnyS/4jjCbgto
NWSgQvp3G5j+6dSeWGQyLI+RyPMLj52eyNeUtIrGYMOBcMLvnjYsfe5DH7VBS8YUSr3NTwpov6/I
8nxKAsBFVYn3NwPe7+cUN5RpGiKE+2CXg8Obb/SoRpx/ORwERBX9ktYI0R/E9TclATnc8bZ/Yv+L
glMciKGEN4Co7SbPdY5ZlWG7glA+0lkQiRpIHooKVvCAuvU1Yo8ZcNUOnl2a0YaDsYQmssNgfZad
FnFEJjCyzpmCqHWKep1IPo+aCjrQXhLwcOAQBQkyE5mCwQ+txanEu3avnVwX19WSSB5VCLclJQmj
JqYTKdJSIPC7wWfbAHUwhjo4bvWEosdTBOMim7Mt5EbLx6l2rrQ49IN+z8fZgXYks/xg/X4jzRs3
8ZQZxQOP9t/l9Qs9DVkxjzA+Hx4Ltsjt+6caMgZkRpgTtKyR00sJyXsHURwJydFdUd3mwTeYIKiT
JRL+0RLxrVxzh3HgMTFULHCvu5p+Va3msfR+8MVASAThNHWW6Urp6JuX11TUi7Ke6Pecv4RbEPxd
YrP9nJW6FSMYGHch5wGx4PAnjuR+6LmghSmsh27K8NHvMSLq1l8Z7vBd5TCH5SW27mWJ6I3ApJcC
q81E2Iru9LekDnGih0n3M54cb/tYp80fZiJOpnLSDTIuDZFH7BzPhxjkvdLx48C+f8hLqyf3k7+j
hBXtS/cRnjNDAqi2Uqw1LSMsAgJBx86S6w9R9HANYXfxWpl7sM64W9pkTs698vKIggmdCu8j8XjB
xGu0QJfRlme+2t7lhhzZCYMzHOeR3rq2Empws24zlNiEl4YinpCUCu8J8hRNHb5mSJSyHR27lH+h
p5A3TlPGmDqxnAaDiRi3+ndP2BF7qvWBZY2cfyFjZqSaQ4YsXlZjdAqFMuO87vDry9cHFiB0M17Y
8x5Sc1IY/Hhh+aUmrxCnxQ8yDH7eIdBPLNKH0uOPEQWOJabdY2MObhFInAqieVlaoCsDMQekAVea
naNRLH9mGikleKboWNVbpMU+pIKB9wmdw4fbUr/NJ1IULcPkgeQ8fCvvkxWGATX4lpdwk4zPMpIa
yMMzaNyKjHFw5X/Da8nxUqwkqepmtcMUkPDOtztBdoaqcI64nkS+gphgVdG+05a5kY9xL7scywYR
Ke32T7pcYlVihfDNZDepspzjLzGb9enfucaYi/Etm31Q/wsG4kuXlX4jwvyqzM1JGquGaCxR3lIp
Nkubp8HvWfY/KS/7jCXWmO6t7YxWAsZb+iNUzHWxAbYV6c2vG9zK9m3x7vm5IQnxNsztXIQk2/Cq
qxNDvkoW7qOwGhwWSeiZN5XbChdhxNxV1pMmQfYZK5+xbjquJiXPiqZutloerjdJ/HuEEsSpieK1
IwDPguHd6Y5o22MmjGPry17hG7BRZuVtmq/6/I7Feq1qYLGIy+8cfQb1cuFEND7MXfgRg4okjj9m
oBgTks1UxgWJ3+Rf2k7GSFmAZk4n3lgnOYl9OPvQkE1FsRwIY0WKImsGwR3r3PduZk4f8oCs9QuX
/ZcCiQsqg6+5fDLx0tv5hCxp8dzjISbO0u57drHfMYddRlwmwKxZCu6Vy615UCVGq4hTxtd0zFvn
8/GM3TgKhl6J3QNFHqTALXiAUrlwjKAocYPSKy+HIHvkz6Galjw1bRykx4jQvyOv+ZZNkL5p4iu7
Lqo0L6U5v91zBy5NS754Txud5VhBa1cbGYD/AWMLtyzITak7FA7qs2xTZdif1TFopYRVa5ar4P/i
++L3OSqeHNVsVRfE8yQXaPvBlfOfQTQdGN8DrJf4QJa44RV1V5JPHAccl28UIMRL3zuujY93IMea
87wtVqjrG2UGGgrdIq8Wdp6PnZ7kAZD6ZWuwAWtDBzoIuOgbyYpTywM1Wwcl7afDup4oCERfLGnP
KALMgeltaVZaIJYwar3e+i0q1nwoTIm+lzRy7xwOEwaEsrbSonUR9y/O+Xq9t6AkKCG6U2+3Vzx5
6GugfyRflLwpW88m1jGFGDxol792EpOhRagPMRiAjYH5c+Zh2UiQYWlXeZ+5OQUkuyyKcQrmb6xz
/AMvmNjXGrr6vO1zrg3ge32CBbt89URHai1K5oncZyXBNwFUBBCBCx6SUh+EXb51ddWAvuKK+0SR
SRLV40WSRFt4pkZigDsfzeUAtMemFRePruHyrDshtGZYlztWRcrxQ/SSzZbe/iJyfb538x5r1sfs
zYOdXeWNM+rv68iWE99mPfnD1UGlJCA30GKTQbNQmnX+QYv4hmXkU/UohaQjGJx9Y+tTQZQYeXwu
xvqcNYqsyX1hejBX4o1Ed5MyTZ7SdZz9DyZ99YoLf4R40Tjhovu2f0bSkpER5EQFtek+KDMGzQkF
p19t2GTqceVlk/R/m6Tc2a0RicVWXGRUUrYasXhLtXlizUF4zT08s/ASbkhU/byNqEfktEAbSs1F
WeY8Hkje/Z8LNM369olyv8kn5cKd2HMZFdBgmwejTC61H0Fx9lDFs3aKO/od/tH3lOV0MQfFdgxZ
Gqo8wgX/jhleJOEpIIsDicmBHu59Q1swqi9/gtidYDTXHZGcWSMyoK2aEzSzElLu3f7R7uraoxhO
Vlc8F87lYTcwfQbvxtTXktvEOGf9qOCE/xiPwJcjiYowzhki7B0mN6HnPQCvvQcd73Ndqjer1qsw
4CASlms/Yo+zNEHGJgVUkHiHj2rkACIFMsk6hoKCBnpH1mQAcZt20OeObqBxsay78NDKWR9MV9Yp
GWudWW7s03NxiiaqVDtAgT/K/Krw3GlVbGefiZv1mwWd1PVD98rIG8qhlkEciIF1OS/izDzbg9b6
UTebCPOxncrl9HuEeZaA5rmt47c+JVUGNnXxu0CIgIVtzivnoch9iFV1hn+ZmUH6/1MtB+5bxaKf
LmQb2WWGzryfNiScvXdcxX2UcgRMObEXj+fUUXG3kdrdDwWr2NF+CovbNPwNbpYkK20t7tvphQYG
4JIpL1MWUi6K83fE0zaL+4sCoA0xB4zRSpsklcANhAQaKjP/605FY/S6/ag9Qa5UUb8vMTV8OqIM
TWF3BmeAf+dz5Ssj84BdEo9M7Ej37gsUQdaxD4ZI508KBgw5XpDGB96gnM2OBdO8cfdGRv6lvzHy
zoT3SbnrQCBlSehKP0qCTKRd+BCuHeOuv3VleCMZXvWXse/MEYo/zXzQ3H914p2Mz+0GMBnToLyc
LdX6rlprHKKpMVmaPYpY4IHjnhPxE+X2BrPzuuV3mCWSLxjCtiyJqCPqAXlOhUOE3wzS+gTtOlPt
Hf8Be0hcHGwGU/liFkFCjt0XqRRxFh0YN+gTqPUAB9vaYOMKIAH1OM+QKfxaRQr5xBvsLYzcYCV9
bBf4wd26Vgn2XBUvatahcc3GCYyW8SMXk+FbHFLiH8Cb6IaxaCk+6Uzk/U/dmESydMcYDUi+2eW+
WGnk/RaXMO87bTaCTBNeFvzgru88Zety4quouvZC7GC9u+1cxkbKEqlixFEraBfUaRVOC0VSOgfu
JSMYfRQRfK/1neGiU/aofUkB52Jo+7CrhubLB0SqPTaS7nFkgwWO6ti41HsWY27juEF/AKd+RQWZ
ADUmAe5QbCY8B4IL7eosFOXLeysF4QHsonsjbhB9n/9TYWlr5kGuG8vtYbbpzd9i8Cb6l/rn13Y9
zvrM7sZhLJ3lKgvuQBzL2bQM/+VAsYXzQ0Bq/P2ovhPpFa8JwmIC+lWCdn2Dfsw6Jw/azwcQ0e7R
iIUUDdPPxmRr27Wt4HS4kq7JCLht1ayUANQqsEc/NfFz+d380AEKcTj3zrgCXnLCvtPlG2myr0xo
F836ZJFcGdfOYSmBKaAZV1LuyCNCaHXn4jtutchsvr0hA3OFpmNbUCdIodVKbFHqMWWIqfCxWrK8
PjKdj+jezPpzw206ch2TML/v2k8CW4TlhotE2bQlulujhyC1JqgYDcM3K9GCXaUU9TebySMZ6pMc
ubqqACZe2edpoHe816xUNh2htl7kZJ+LqiecjUSjHeDBxPJoQ99SLXYnKEWTi+XX0Iz7DqJd1gaR
PA36FS8Miwa7zucNUhm2xrj+M8hrcbuchb5G2fe/DVIhMuDHojQoE7XfKHSrZDE8Ozvwr3O5xxTA
umXZQ5Ub6LAR4iNsNz7Zytpz+MSdbXFBLYEZtjhaS3tBx9i1fVWZMvstj3m/P/kMXPSPhukCrZ5d
ByIiE8P8qAx7rz4YgRwYBmjeoLRRUC2AGLYrf/YPuqAWo3JbZ23oDc2ur3fWF5/BbLsgzkou6I+g
YemOnvKoGcTBkista+N8l3/xUug4Ee0j+Ikfa05ed0xrfPicunAo2CL8Q1eQkwPCxuGn74bkkVXj
MFBwB+4RM2SKAdp2iDGbgjBzpHswo+iHiaDpXpKydTP+8sDJaDWFVBGgjzmIMnt4xDmbC1IyCnK+
aPx3VlrWRN2C9gwYNUfzYejUFYGuDa1G0aAKh+u2oXOOg9rpEiBD5/IVV9BRAG6SrtRdqeuYVfqT
h2v4jacApQkf0Rhv/qRdLquIYqJsApr/hzNDLYwGa7L4ihP6FQ7MHYIl9fOr0RSfmcttmOotJrT/
EG6nf0zw96pItbVRL3GaH7Gu895C9tiqIXvwBv8vVKPs53ZWAHOL/lbWaeKudubHpLgAecdegxcw
uu40VLRjO9o77v/Qafbkv+R/IpAx3sPzCk+8O2VZ84390lQw4Y7ZXVVxNEkA4+q0EggkYyWYgVLf
7pHj34zqzoXfAC8h6ZGz7ShtFes0l/B4fIk3TbdpKww+LYVSGR8OT54EVUII5PXO0zayRsGGLqE4
Joszgtw1N8T9Sd/MsCLA70EEhVjW0DDJQS6SRJMAngJajXSqhpmM5Xukv7kR/8IySsMeEyaZ8Oap
PkDecn8ySwZ1ZOP0jIcMRuH+XdS7y5ffEJesrpjD8ztC5g7rv2gK3wCRmVfvmi6XJRqn8bBDzAL9
iSwgRYDeOttHreeWGyYDIxEUEiZw7azKvENA4ZTH1Dbo7LGjGvR1mll1jsJNlcYwYVyp3oGwI03l
BFvecEVxhT3nP+yG+KFXefMhUO4+CWxtsdLa+NIqOLmYZ+BltXXbDc9VUTzJiF8bmSMTA07PG7uA
ibayhSTDhcEJW0bpSiB8+2QrkQAll+gjT1Di8DPhRvnb7riEIMFnNEW3NDTQabH73bbXAFAK/LEP
w/GWOGPUj5bmIsmhQB5+2Oy/SyHPBAL7/fRkUi/sxh56dehLad7N2cVsve4iBZ14Du5YkTlxX8ag
w+XV2abNROFdo9GeKt4gmHT6RCEVoL+bGlkY5UpwefI5z/OCTxXbnzmt3AUEd1ItzyXqN343SvQZ
guW9f/qUMYiMgR9ZZoCCfMIqjxIVy1IWADh79vW/aNKsf1LuHtuH1vxSLxUyIs/W4aI9t9xYKvMn
dSxKxvefAH0geuWp35QywRczGU7/SKiORxehh6yUdu5hTGxwk1jC3gSWaXFIpHo+KbQ7aynErU0+
2SP9slbsg8uwD7kW8wViaY5i+D5udxeaD21a47TOVc2zUF/HBTvsajWIgWmhJEXyNZBMygh2WZn4
wa/trOz3tNpn/2CcH9OvJdLt6pZeeSCf8ag5JR96bBaiXpSl8LEB4Ac/YSLUrFvm+0/hnAQ2HwvH
q/GoAH82I7YgFe1c5XOEO9W9n7ayTaIHnG0kPCt8x1KhGVhHR9bvR/EHo1jgUd0XGZtd/p4XEwwi
vHwZMGfisBbKwHQcRt4ICSkZrUIEuLpDVnXUL+NE6rczAjQl/SArULR535ihOxqWF3oODC2JwMrp
RnMbBfnNOBhnDPU4ycqfYHrYMKAx7bZNu8KzpDecCb2XX/L3DscssLpGosg7XFOUTvB9fCMyXw2X
pX83uCk1UqVmraPmXVrYbva5/pnaoIOH5yEaTvuOesaeiFZeXpXurPTFaaGRNvSjj42RTohn3ALO
5pxj54l9KMdL/ObbMyCAeUT/TMyigsjCtvlek/9koKwWtKaKxTj60SDGePXbayehIGKPp28wj/Y3
Z/Iqxr0VSI+H5WUSoFfkob/shSJtc5Vcpr1Z3VtwgvUJIT2bXzdP9wRmfXWaGoavHmiIzFAIuatX
yhItY3tEcnRRjMmba3Dcs0QRgKSSRMQZAYNZoQRoWVvspAZC6Xl6uuJyoplbnOOIaZXCIPki8i0Q
tKwi2k5MzZDAJG265g1mOIdTi/lLVrOnwOSN7Qcn/QI/Yh2sOBXv4la4fZeLlamH/TeaV5/CFNS1
POI4UzJDbJZd4cixxk9wzXZZt/OIa1mJj8XJpwi0deqFd3f2IJ8QKW5IwHM/s+Qfig4kNZUEOlpK
utm/kshp/fuT6AkKAR7XFQXCiWYa0zxGdmV4DmI2/ImhFgQNSzmE1ca0egnFLFn0B7cjzCcCFQ8m
II0NvUlEgnZ0gRu/ktElgLAuiemyhQkTM2hYaPDkMwOAMCm9fbzT+61f5ohItl6nCNwe/Vm9tsHD
rAVwrY0gW9e+XukAay7trtj/5wLMQBJuSCkDmP20yfSEkaO16e21tfMVszq8sqMvqYGhD1jeTulW
VAeRE3jtiU0ONMx8tzzSLqSQ06Fa0+GEPFABMMwGDXMePpg7lZK6cGeJm4WaMOMWA06aVoEZAqnF
Cw0BsAsUjjSKxLqxNodgG9vonGU9ZX3MGTD7M7piJZ+KU74zCBG8UUSJx0lUmuuNYl85zFsPDhPz
TjraQWN/RwsBWrPSmMFgu9h5nLuD5kqH0pYOlbIkk733zkL7cwrXe9z5tF+BrcX/QD80PGz01Kmh
BsWB7UFWFdH3QNc3Airt8rbTEAmjawwtVgJcFSdxf8JM4I7LMz+FY2u1+fsDMpj2MV5rsJA9ugTl
WExyjnrKCdZFe/G8X+qMMmM6nwYyn6xksAjrnJxR1E5usbs+R2DzedtxXqF8uPqO8DtmZ2nkfYPf
faA3bZKPhiw87+kdybicz4tB80tzKpmI7jDMOVHMMhRpinyKlJ7rqgzzmSZcuoOh0XdELDRbj/np
zmsZd9M5D5NG+6xFyy8D1L8laRZqiSWm+aAq2Y0cal78EnfzKPqbJiL3JJPb3yhLQUyph0QGOlUy
IbGsmq16uYRqAJ2CWYdFaM56WJLW9MpG/2YtH0XEvul82ITju8qu9A6aCrBYfZq6lcqc89G9GLRp
ZaJEc9/19jLOd71MQxVl8jTi3b0NlCfw51viCbdiQBHHfEdhpeHSzftwFDye9fW8slIuO80KKQWl
vt6ES0DXu3jN0JQgYliKPA6ys0mpmdceNqR65ghM0qmBLSJjHe7dD37gFds0fd8dWwAhYaZ/vhiA
cMowoFed4WCAc4DBAyEKJ3WiZRfGvfhPRbrNaMv/UG1t2RPULv/yfq2hYPfyx0e3U6hfWb8kI6qh
jxiZ0+ddJsfVFkJuZbBh4IuESaAmmga9OrY2esmayqUMS1q5h6iO1hfpzQex0kKsVfC2FEXXQC+L
7LqqEjSET6Two70w9roJYkmbFUV9yHlTbB3U7gd+iQ11uOXlIgyQmw55KoBum7N2QqJgWT6u1FHP
hhTD4M6dFW+9AVXA03nxGhRqNQBsdGmtI/7Sm19fvaxFioZTks6o6GrELVToev0WtsmXCPNPiO9a
JHmdBRKhwMN1RqX9zU3AUsp2Ri18hp8bFndL8vA9jEiqFzVHCLBEzIA0Djhf9VphjrGJ/NaXfs9k
n5SJATXXQBaQWUT2z1yzUSXri23Z7xvFmtASkCajCg4xc+FmdTRwY/OP1kejvYtB1AEIifIYSIEr
J7VAUwhUlNAx9LtQtjuMcgm1X+5qQ4RFDdfWbUjdIQ1WlpygQzOXX3LoacjCYLivHJkALjEXybno
tQgbgD3IXaxgILo3UP/fWypcG/AW2DcJauCUKt6104P5QZoD1giE6F5VgVAW4yoamwf4KR3ylhuz
t+Us7JW0VEFB1rUUBzJ8tt2d1IhIzPnmD/qYlw+1WXNx8Bcu9HOZ6hzwlHiO8C29XDyEyOOdOlCA
yGNFsZAUenYfVpuuY0kugBVEDlOwZoqWzOR+5Agi2VftBpOiNW4NZIPpoVtfWG10KzqUaylRb+GM
mVRi/q3PE6juQVYjhdlhooi+9gKcO7r5rcWJAlfGmSFjTWBTItxg63JquAR31Wgl60ajhhAZKZF4
Ph8Wf9iizkJKC5Z7g426x+dVdHUBTUoqGtykeOM4Y29K8zsVpNQzn8/THvwARSqXDcCal93blx4m
xP7Pzk/F8KQqXx/DZGTrKifWxezIH8D5QlgP2ne1OJ4dAz5PoRljg3t+1MRz33cMBbAUPD7UWMl1
YIQTf7i76whUhjASCxtFjUKx1dDQ9QvlAAXE8ZKEXkkvrk++1w7O2wC6Y2lrOev+3ykBlJr0bmvk
MeDB44aYJEjRtOhnxqcI0UiawoF/lGHmXRdIzqVXxgRFIV7F0nRhzzRmUgz2yxkKy7LUFrQx/u+i
WSCWckFu4TPTLa/mJQr9hhhsM+Ik2b8MULnkSiw9JnE1kKpXtCyggURldEmoYJaIsFAHW8tdkF4J
Ixh5f4+dbrYjXWWtSno3i8TpKxUOcvTXl1wHyRb/nBOwOTeH19fXWqEdOitdTlz+woSAEw8Mc4JP
b3cGGrnqVbX24nskb6t9IxU87LoJFqaiJ8L+wR9uQN3vgH0YrDWN/62I9GNXIbiOAewqmVonDwho
/z8jzWNuYODRW3veZDzmAmK3PHeOHJRglK4h2MPL9y/OzTU0nIZT5MZ5pq8NEep7DhfiNnAxYdFz
fTpnkxlvGo/2S5U0lLDmZPjQdhNek7TijcGgJD5o7FDTxwD0EO+70TXpVoBt8/ezPVlhEoVkTTpZ
idwi/GkeNz3mMskRg5MCv4W/1HTx6MNcQmCBrgtJL/TZllTSx8bFVa3nwvniIRrCetSw2DG9VDE7
CWDMvw/V10nxnuSvmmVJG6s27zbPPVSCbKWDEb6cEJm2JYGC3vUrcxinjBjO4K+fiOUqSJXqnkwT
W7x1EDImA+w2jqZuub/3y4lZ3y0nqZP5azaV8lqXg16JHWvuvmKIcYJKEOVq0rPTSpm/m/8dtt29
pSd2TCP+bnOhwWT/gdjfR76068gzUeuqeh8UafZesPc0cphluPPzfE8T90vejn5nGxnC0wV+h5dJ
Lo8XZa30cutOfp7ImpYfGTBjxzKjiA6VhH5b87ylKhWeZ7FaJBqM2C7seTtPNYZtNb33ChMrSHBR
k/nL6BeEqXVXbtuOz+R/+o6c1DQpkbPyEA/QagORAxMebkJAaJwM61zC89PC46Af9eWt1Wpv0WRU
XtSswGOtssOx7fm3ADkZ4ptS5BOqm6NdtfIpmuZwyB0oBds2CnotNo+bzd4PMfy6lt5HxODqrxQe
WK2MwaZAnoKqlFNWdhD55GwVVzBAOF3wG/dntOshFpkWCg/8eZpWDzFM50Z3t8PxdzUKKAOHcnIM
vn0vKBcpRX3gNRkEJ7O28WT5oxhitCJ/Ug2v3EAjVuNCFxxtMe2Z3ghh6Z2cB/3vxpJM9Ml1zVPE
YWTRS2uNET5ArUBoonyL3GanFrFM9axVcSJpRQ/kOtKRjlGJm80Pvkull3K6c2pdVWRVVCqoJUP8
aYFZwWRwAuS5CcLQ1+ENQ7TdMaSPv1/CJrmGr+Iwgniqh6zZVYEBtrI99RWoWfarEp2Qrd/rFHH7
avy4k1jA49dFF8RIKn9Ettn8kWgoKHI6oAaYTWefEx8MmvHStEiCS0AZUNNqVIDlBJS9494i/N3R
K0veKTU4Ytl31afbKbyx7rhdTLkQcklTCMxitHxEEUU/8AK1WqmsB/U209OD9KLHO0yicp+gcQ4B
ukx0euVFku7kmJ5Q25+3eLrNtFT9pG8AfF00szisUazO8E95l0Sf36EdIn1ZMbki+7+BPNs2FbEd
CPcrOG5YrC7wbfaW8kXxqqEUgaqrZ+5coFBaETmgYDu51ud6jT3NE0QLay/LnFX1bJEfGT8TWen+
t9mVIQ/8990pBO8SHT2M3xp+lsdmmKNJx1nFGS3s0qWyRkJW9Ir7KaGR/Bw7zQlxbGsCgcet1iir
oapCVkWv+jEZOTYXSYf/nogdCp+z63Rd8o++heJdufjeRfgNo+Bn07Jow4nsZYDRvEsOy8nXH7+j
vxfckx9GPEfHQ5hj9khrjwUaDVxN4b2n23aDMcYfhZfB9JbKWzJhKEYMcwjMJhc5iU31/5KX+/0E
rJK+9w++fF7L1L1fy/hSw9I1GLnALCY2DSVs617n1y85Mwvg8C/pdYqX0rSsLelrBrzJNGJLjpdL
YULB7zWFEOTk9fvi8EjCVEM9MMaS/F3YU3lLaTPF8dldXZ9d4P0qhZrdpxe+ngduYjjW0eQ7KxM5
qwgQ3CCmkUtOo3E1DtxNlokc55AQhdtbza/Y1Q5lM+VgjQBrYe3l83vpxH+XeOZKESDxA9xUd85Q
o1q/mwUtUtBQ57BcFoQNZt4v0riBeN8ufPokXIOarsvNjQGJUwACbSb3OXZ4Nca2AqKMPnBXGFvk
KFBPCOFHyNmu3OHXEukpdG4mC+D7fkTWbzAItVm3MtmDtgSg04fUe9fSSBI/1XNSFZ/bmmbiO4y0
Wh1126HBo3uhBUGsIWii/LNCNQ4xtt5fECiHpL04ti2f6bkjyOiBnDJlnyuti4gFwnkCoAY/T/ex
1vIud4DbMgdifORZxR/jWoTWj/5kPuyfxls3CXXI7qPaNL5yQC6WACeEz1T8sVaKJxZjZ42yGL6h
w2C3/s2QoCp0n8i1VNsqhLrw9WxcXyB/b8La9skhpV6o2qhS61MRr3Sc26PQjH/CW3gluT+yTssP
yZsaLr030TsFn4nHTz8iShRky9dVhz6NMllV9/wKg4rrLZ2QEXdDOHWRzHUIvUml4r3rP0EAbLSS
vWFxc8YkPdNeFlwRQ7flA1dN6AMMRL3EIGH3dSEyN2GxLWJEJ89qIwa8xzxXHVpuRMl0Aq+HuA42
eXOMC3h+r3r/sZxDU2IciuZM9bfAQBznQO53cP5AE2uw1M7KQwe7q/XW3O+19j1o+CNGRzv/ynxT
Pq+Jua+beZQ28tHpomDC47WPqjn540qahndNdrd9VWfcfH24D+d8NbUmOzeGvvNA8SFNEVjHJ+mU
QM4gL8DJhvkFSqXs1OPyi2L/kqgEdhA6588IIBWoQgAC5zurmBQXU7Stq84rl6J5klyI2PFzJ2U4
WyBAWB7zASXA7ZZqfa9wN0tKCi3jzl0GaznUk5nNgJRptpGig4XvNMHoIYNeIMhqcs3CgvDgLQAb
AfcpYJtRPKVAZcqiq0DOB0BDZqB5j5dD1qsWlKSaUacOTB4GbdMYLD1DBaeOdbB32KNd5xlA2bCP
73aol5ctg2/9EkCbHHTpI79Gim6ALTLkVyF6rP7SIz3WlhtHcYnn7q1QM+K5YxSc7pnQGkktIitw
5so39ULUUQp7/2N4Xycsfh6Pti4PD+Gmb0yehidnDuxUkUAmRvMvCzyTubsVDtlP3SDLUaU12SN3
ouOixq9a4nJ03Lrep6Rfxz51AiANbdnLow7+8stg+568JwWmFcrfKMRRLV1RkGzwEIEuFtWike8e
MATPnZf6+59TCaq8w5JGhcNOUhFgfacFjm+lw7pTI1/GyaFy1bBzt9GCWUJ0KE4eGJ/GuvRDQQZW
/4J97k4E3nMtFllmcAsGzUFAdV581tRKTu6dpYoPQfPHmm0S0MysrDyW7KZ1E/ckb3C52uCxeqQ6
4UFD5FlxvM0j9xSsVAOF1K6muXhx1qy9ZeFmpNBAZayfPRlKfULhPaeceUoT6IREISxvCfdPURHP
xMZ5zcXo7Hqyz6ZsHuqhbKKOj9X6pq9Q4u8E6Lf91bJ3B6ueEvhKgMLPEhjjXXjSiEpPoHT+jL0F
5NL/be0rRfhK5Ia6tXW57tnVAWIOgQfSKuXbnFPwafcc9lNJSZmx5n7NaoAcpLHyWZ2BpQTRtgL8
krl/APyxjd8IsK4SyxFJ/pjTMtc3iKajrehfawJHDmE+6zslGQYGUYl9HFfbVNjo3aNiNzBxgfSj
lQ/hgG1sQQhB6GT/hVtl0RhL3B7KnqzE0bLG2o/eQ5iUnURyjGoVAv1KszOF5VOhRLcbVGqDZLQU
x40HJMhfguNpvUX4F5+x8mw84doXwHTKn25LkjXS0x0Jf6/2oDFMDoV2y6r7Ah6I3dDsYa+4b+fY
y/i7IN2Nuks5/ASzNmsf5sVHEZs5+ONr3Ra5UxyeQV+7FnH0eR/t91SuOQJgsyesWeiKG5BLvGaN
8YC612LlxtoOuzqQD3tgF3oeLZHo9Q0PSELxCiz42iupxZ/ZyhlFqR/AIAKvfAvtFXSQhAn/pj+V
EORdk2CQHVrQLBUxvO253f5ao4zw+D60aywps4zE6U6Nm7jeug58xkqQPz7RBu0m6HNLm2LEwOsT
DtNgg+kPpkcgb9iwB2SthylOZkCd7HIDIIBFOQoEYj6Qb2r9Y83pTWhOQ6RLySrJdTpfBAigo8nT
FrWZ1CqcXBxO9stHQpySN8kLYcUv8jPTNaBxYyW6ws9dXCm5WCIHoO5LUWqYpOnIT3eNJ2wy9HqU
uR4o4+mbAGpufnIk3H84bChj+OPbeBRD8QiDasIZgr2Qx2NUvxWMUK7uEYkAwL+RE+z23XHSaW3L
T7eC9IM8VFxwVXYp+WTVEgySnZodBF4omAG5rQEq7LKu33xO3nNNaqrrqK22zlw+uXNoIVVxiF9Q
Y2zmzMju9mMrxrhC9zs8llxK1a7FijnkF1mqZUQikPmoWpJHSnyc0uFcMgqFJA7CvhxR/8EDzTsk
uMWRdm19HuMUzWnYa6MuOdobbqF1RsiWvZx4OPj0mNgVdZTnuxSo6XlezDLzTrgSNFyEemDw6+wZ
JcpxBWCCBqO9+19n08Pprfr8JGMlKfOX8JyDGLk29+PcCK1EH1JKwWkstsF3SE4qV8XXTjS00azE
CXxNe4Ar/yyCM35xEtZl5sKYVzWZlWwgZirlrjCzUHvjeFGeB/1XSV/MN4JI4K54ZuFpgFi0fxCH
70cMVPPU8X/trTu7bshN2010eYP4EtXDoKNVhAMPd19DHJIYEcMW4YKNYzJPBhXOXG38gZdKY9bV
GsV64w6VGytT9GPQS6huVOPINE8oGijk5PJRsipOEe0lFku+Wdp7udTNVPqMGZeNKZHqLS0ugfZb
HFYQBQBGJqtUl6ECk+B3EtIz6qsKIq3ErsGRuW+5gswFGssGLuJ/THGi39A5WcG7FrUuRV+kMszC
Phj8PoWCLtn60iCsZp1RHdhwpBaiiLL1iGw43It5KlyX+Vwiuit2AGrjmmJaFe1XtszTx0/fBBpq
1JAd4qZxthDflLP1EnDIXg77G4OVHl66YfaNHChtWlo+ea/Kt0/DMytIgBqPuTFPzZv0e/+pLshh
MXxxUGoL04qqqwxbplv24DEoO3iSMISzQZgFz0bCmnD33UDaXbINYl64mb2gWNMDuAS8oLYWtcb4
qc1sINyAK0bGEzgPP3LHUVWJniVTqivBeV923tcD+Ua1VYoYWWL/RqfQyWK5yGAF30pmpi2UWu/g
Z4zGFCbL0qEuyR+S64VGKfdZXB2EBaOfC8bjAP5T1aRuZ2WxMVfTSCEyc1lQB9fLCsJ3siIU2RID
HctuabNz5j3NAFc8TaMGL430SmF7c1qw3niaT2JuBpZCKVIk74Uk+zyDX2s4K+Qy+3tAwhjq5/uw
t5t/DALrCsmgF09G4wfAzNAv3meGEhSyT0ATdJ487B5PdRAvIT5fSV0E9A1VbpMMwN3Lx2kxwBF+
9qdt6mmYtnVwfg5n+QtMBMh6AgphzrM76zETBG2kpOYvzRqRC43fYKYTo/H6kCl7nAOFsBZU0/1Y
l/GzCDhW7O6ZXAgQoecjvwR3VOik5RTRWqTHw2GUoJwWzxpwWnEVldZw8ZUyhtbI3mubsCmaMDqd
p95CKBiI6uRTBWOPFa/Gj6TxVAT/EC2uU1ER0SG0ulvmuphHuWZvozC4+GRIF5LZZRDmVhaSVFUO
OzA7CQ5y+oexlfmLE/ivLlOLIr4ZzuMDWIPQ/Aew5OGB4ra+CKt7NFfVY5P0eM2/ynqoYrfpFneI
3i6UFQXgccWW4Cdzl7zV3an5h0AJm3Ukh8x5dSCzfDbWNvimu3UTCEJI7ZOC0eW8PLlCBB5L9uKg
sNltfXEUqAcFWMzbIQjm+GbXW1liCPAsPJqHdWUGEj+0alazPQiIwpzgRKHNZoOOk4dCkbcIJRTM
7jtYZUtxhabEqOyVEEXdCVn8V+7BVl8I5Ax5qDkd6tMwjS7OfwA8je9y93wp+oIJYvKTGiM6D5ci
uPM5hKNgLF4fvJs3fwATejD9/5xJY1LWbhbAcrkeJ7B9BIaKhNwCjO6j1TY909NJhngMMimmpiPE
SLS21o7ofd/xBWVdVZhgOT66fqcpsL8tG44N0l9OfjkA3Wz/yN7id+PXhR15xYyeC0stu0bRef7V
gVpHZXX8OhlIJgRhk0E2fmy5UKD+/hXalvAjUg2Vgr5T3ourLe2GONXTZ91/fMOlsW5zxc4PO10t
c1L+5hf1viWhbysFThugEBMUnFd09e/P1BX1xZEg24jMPH9V6qr3vDJ2blBQ57GOHGBuOs3TnCfr
9L7+ukpWvRZ8w/94qoz79JskAJUwHOliaAwon3W7WLfkdkVbg2Q7PlnDcN1IH7zPnQ8VNjkL24A9
eUvtmEsjX2pMNtPCZBq6j/7bTjHAX5NaZ/WnNxDPL3Zc5zoa/CGo5lEka3uYwtjX2+wSwGpW4z+o
E9QMpjUSnnfWA3kkCCId0HhfDYG4AAX6H6XKcoWgrgE690tlvNAo8C87cOGD6KKh7KBpmloHlntO
TvxQPV40hqGwiz4nw2BFP2YGezRKZouTNvH2IZhTY9VMtJK6S+WHOv4dh2rZBOS0EzPzWwDeilnk
3nKt8tYX1qYSn9erU20O6LEtfXXOV2234BEKyONys62l1tY/S2FxcqIzSgJqlg6nYD1v9EqlH0MH
TW/txvAFltkSY3uGcAv6++DIBYpFQFj+I21QAUVGhMo+aQihmG6El+TwuuHOzYDGrrvTi/4tni/j
V+1J7d084wS5Cfa2jujzv1bakftiyqnlSnOiK4sB95HBmVtZ4tJnkwyxgkFEWMaWCdLbUfc0kiB5
+sBNZOS1Uzx0TUXieU+Ejf+kcCkvSJ3YUyYjeuAYT6dyMHPIj9e6X5f6L4L0R1hr2av0D61hNnlC
C1/UAGjgx7xE1JR18U5XKlzBQ0BOFIugPidLLm2YB01ZE1+vu3UMJO6rFLrG1fpzpocDL3SQcqnq
lipZhkVFUj4h1yUvMH5dT5OsbrJB0AwhOwFM/CeAD1ZfgOf11OWjPorbSEsB78dGwrDIZ421VaCg
tqZmZ2uIZToyPcLAMn9YfPVSxB0YJEryE8wjxSOD2RIuwRlyifqamTDkLw/mUYBSeB0LoTMVemqv
rojybeUL4OeNEpjr1P8ifBzC2ryNo4dMpWNYekP5FdRTzCQAIlXJxvnQHuzh6fDZeCj/KcD5VDbW
rDIvRAZQKskrUKJgEATtzr5r0r6OXCcxZaikeKxAP7057t2bONyeVYbQcf2kO5D/3gonnJFVNZEW
cIonX2DK5++xvlF5ZK8s5nVlLZkRDx8GStwHmckvTpHF3y+KT3lkVP/+bi/joo4hmiu5qiWO6NSV
PUc3ZJBKU/IbMq69+BvP6J+ezoYWr2bOFRSKV8wPEwBqiZX9VKQRh+WghewhFjNGcN0lXVWt9x5q
lDguMVSqZqAE0c5c7vsg17ZajseS4vyzrcbfuE9Lg2fynfGoERFlwuxC8VGJyAq+SuGS0UhiSXvY
jALWQJ0bENf+ktYcaUgbfF168f4tYP6jXoHNO2vSWG9CYWeu/ZaYtMLfxKat/k4Y+/5wVgN6IiFw
VxOKP8M2mRdnWlEUz+mMg0bsIR/H6NpFk/Ohrh2XhirjZu12Z1dGVyQbu/dKSO4q6b/qUa40NKCr
7XA86AeKnHZjEwIDbGNIS6PslqICLUCnK6tXQKjttxb3XFB3tqGZbOW6CBoWY+7FrzzAKzdTzCzq
pm7mYb1+tZVwJbOFd4+m8J9w7VJMAuH44+7jUvpMCCnkk0LQblAbE8q4ojlRSvum8wgh0LTEYS3N
xiepIgaD4lDE9OZWE89atdSVs4aAyGj1myYt5l1IcuyujdOL89FA7RH0fRES4WWAy1VMPAX3YJGf
tnWuASnX3srG3qGzR2v2SFwYi2ZlsSXr3RaDaiQ4OS0yHaO0WhpZQJ8/Gn4hR7yjpy+aRIYnthA1
Vj9qnFmlurAGK2vj/CAd6wBOcxA2VUFPBT9imyizniflepXcUFef3/aKHKF1r/+M68RIWWdfa5AF
Q81FlZGsImZGHC2RZBZLXVc8XAWA4uGjra1UyAVw309RXz9HTcj9pUS0n7Ns7qkagaopdZfJwiMB
6IVvyUCOTHjhhn+sosKkDk/KPLDoOKEDUWfMnKLsMXJHOTViytmtAckw4k6+sge9xsXQJ8gZg09W
kPlZodcpXKDuZ9blY+Xsj6ewHvCLxgsPjuGEREoQtJ/kGtzLwj1jOGl9WPWzoEFTmuvex+nsgGod
vEv1hn0QrkoFoS8zeX4vQK/oW5ijyKjQj5U/ExLA2QNHwwv9nNQftTqlWRh7yeJU0F8AcT4+2fag
rZc2yAJ33qTklNrEGIxiZ/6CEKNgzY6mSCGQpz+hvqevBgPj2hFm/Uh3izm0Ofd2Ixdew23rLjeT
VxF84MHx1dFMmOpzNpSAbmNJwAkmyXGlx/YXUZ2xJT5D8ccpy/eA+eoVFRdDH6SU3sSl0NUmIz3B
JrvKRxBRomRlWIDuEzz2w/jiOjCE5buXimpucmIEZ4okiRMSnYKSMoSA5Qaw7mB5sSDwXu9pgt2z
3dQPbAEUShVAWEA9AHuT1K+avk0HOXM7DwTdmat38flvqxgPIbrIdkxIpV0DFn3T2fL95H6zANLU
j6ck7o016TBpM0ZR82nhQPnoVj9fg+XCvvmeJ2kOJjSn8UZochGW4Hn3+yZ8+BinW43n0HqRmETn
3PQ0M0nQAY3lb0Guj+QzL/FQQ/1xY3AO4DCs9oRPDR4dVXZS8d9T8pQ3nTv2hvM5pJ1erv+ZxBBA
phhs79ueyw5R1Pp1MLaomdIENop9W8iuVIxa+IMnFZw+WYZIL7w2LZ5K1wWqSaZfYKUs3wpF98m1
FMz6hY8YGmbgvSKWs+WpBVn51JQnXIzMYAu9OtYHYtuVfdxtkkihzMRjiXeiFRV/JvHPKwBZSBKj
SkVATY8SxjVOECemW3XGyUfbzPpMF+lrJ4UotqX4t7GCG62Wu6U+jgRryfkRh8qkz3lFKBQr5+Ly
AfDG1HbayZ4c30/2g2vCBfU+q17VCUcnjhoXqQMqoQqw0YA8HMDQ5nmx0jBy0QFQ4K+vs7qlBjbR
rFxJRONXid5t14/zBsn8OlL3gj3fX3dU9rtyFB/1tWy/NuNgIEGy7s9jc7y5sDwQK9+aVoFuYlF2
2iEfjbPQImUKRrdTHc8flyRe/1ry7AjQFqLlb9m6qofF9HjjhLAmThkW5C9lureL2hJNzZlERGVH
4FCcJxxbEbIYA0NZaeV+Gywj2HKvT9vfhhADd1hJkqFOXpueTpXBP+oA16Vq4v+Mrx6ZS73UZtpm
kzF2i+/2TArOKElp02Tno/Kx7Jrj9FFKO+CGt/oZjdJHRC1tL8/OWlG89OTWSC4UzNQUgpdiVWH2
KAp1H1C4bCT7Hn0rXtiLqZJu9If0Rob8Fg9UVPOra3xPaPpVzCQmZTJ/m9MvddUXBM943zA3Al6S
oJ/bh/V2pJ7KsZ2u3HPSqsoMjNyRzI6gKuRe8cCL+cqIGJhxtGHtpR4bQvoP5t7/6cQSb1T1Gfks
1YS9vtdV14tag8G7WPUDaDpMBIowdig/YqB60kbTTqIOgnM63tP5gt6DlAiOXLuJdiWbhnJmS0s4
yGwVy35DT0ETJGo7tnVitzg2ySkhBsFJBnW3RQ4FaJUsMpjDSV/tejUyCowN8RgdvmNVeT36igrW
5Golh9u3CY3jhiSlirLA2uRdthRqGu1cp8nRVA4nPIg/e//zuSS0aA00/bodIkMaRaKqKIHQ0gw0
6hFe+vh7spMYU6kEPl/3SlqZoLKWygaq86fVn2zcCQKon4JuAeJSESTnUWcyd9wmH9TJRCfavK7T
Wp6dsghmqHvnhE0AmaaLLKphFxkM89ubBiXkwXe/1XOjMOrJPfE117wTnEhX3cmQo8CMA/BF7j77
mbQqx3up99l6VoVdHHyXckOs1y0Q8FeFoD4fZhxzHrjijO+xxBcp3iLGxQeVJchcUoqa4hlekcek
WfA3nkxAaPfidZ48+jbTzw2huNnt1yxPiL2XuvdZZONJTOQiTwwLgDLYy/ttdbWY360Q77pfovHw
XJ0WDSQv17t1GSSmozcFYDZCHp9NfjI77gEmC2sor7FJfpRshnFqUKDkxKQLxdfUzHu4I5gKZmE+
C0HIN3kdNBEYu58dLCM7I4PpDV9G9eB/v6KKdzY5YOEszZioSyr1+jzcubiy+38w3KNJXDPKD1gw
nCpGp0tsoRhaKEXfMj/EHjVZP8oUD4iLVOCJqB+mpCaow3XWf6+dyvwyWNFpHz/LV/LaeaAdiCW7
MS7lgDvvhRts5jh1zsYX/+FVWnI/BoFSZ8gNjDyaejdKaE836CMEKddT19Jn186ZX1sxTWB05Chc
5jmSlW+pGb/9PzDTgqUMkV8opgA9/mVizTPlpm7pff62HhS1b/a8C9xDWw1AAH43YrpSecprXWjI
kS4AsOipy948hs+H6CBDQtWwIdA4JdnNr/9cdXEQCwuD7s6qlXMajpolmi7K3/OiwbrsUjvlOMGo
X+CBO7x3lpdXEurV2bLHFapW30dClF0QPdht8WXI1utDzYruUuDNHKYjmk709nlzUWzXoD9NaKtE
1aeHoLkma5huKlNRwS1XAfbRRnyLBPlPbGn+Kg6LRZY7hGdhcByxWQJsdCAss+xdH9i8tGbfzv0j
O9a8qTNDve9udjH0chdxiFjDI3jDYNrTe8MQqdhw676J1RvDI5smK2cOlDB5wAVyJCDs18c0bTzd
Wo3gfA+1UaV/17vHGQgu/x7FfV6cNCA+3bGG+QMSvH8o4zxjOx1MDNrLQ/QMsPu4WmJmcpC4rnjl
Efofc0p91Q2sDAMP7/QXcD4kyOq3Gu/2kTCrFaNnTyLifv4z0RxwtXC4zyV7/HsIpZ1cwmqfZNIx
7U4/RMeulQH+Dxx8uhsBy8ve+rHt4sWBzmFqEk+/w8/PiXZnxPgy61UrtMzQX+6DhWw3xbhMPlHi
RzAKmEj8AlSuLfDUsfjf1m8jV9C9DJadmTPWCvOaWkUuSh/w1NYdk/y1TSB0WC3V99tvEbsVic+m
iajaZZxg2ZPLxkrbOrqH7od+73TilYlp0asXt1Bm6EzP+c9UZXriDHMgVQgARfG2mBLmjpP6OORu
37Iyu3VGNjp57huhhhFivRCIipa7GXNU6+DX5jjMTCLMOh+D1p8B4p201W4YD6MNs17UxhIpGQIE
x1Ub6EquifA4zUacJO9BodfleooH4y2hc4hb674wxLi4moXNdd+qRJ9J2YEJ9QPiTQjRquLN+e/T
/9I55ftvoEwXWRej3NHbMZkjTgwALwIDbfcN67OkIiOqcuQaKG9XidWxyyRDS6oSOw9Zurj88Rs9
vThTvsEHc9zGpZfBu6zOe6SgVJgShb3Fz7l/D58/dJG7lVDEV8I6vTqmo+wsRwrdDikJcq7TVdlI
GGA+FCDG7wp0DMm13psKj0r+7Xp9BuK4JKArEJLLlVbw4SigFhwHq6hJ13VFxr+DuYJfODSioQ4p
2my2G1wpfpVg6Ax1PJFatQx+5WcykqKgU/ENGE6b1+JT33kxpZHbhzxIS72Jcdq3RXmgGEPfW4Ru
J3wCbjQGYwmhX3sHd2GHuPRO+JiapPxwaTe4JzlJjliX6tAArBvbxyzwk7unUX8X+mPizzYvO1Y/
LKzxY2P3uQ0St9XEGLEigrDwwc+9xv7Y0RtykWHikkHaWo1hJPHDh4TW2NEA29Zdd9LDm7MJFGFe
YcAxFvVjyQBr4Oilg68zgY7GrEtaNDARlLWdmMyI6PZsZmSAOyFjWq7u1gqNjPdc4TV99zI7/FTH
PUHi9QS70CZJS3noirD9/JhXymDEGAqViFTcb78gNrsI8nMrrQQUgG1WGeLA9p/fkWwRQtrVgW/d
8zgN6QsCc5IbhuuVGfpkzpVHqIR7Q26fcFpSx5/3Orup+eJeuUTaayyBh0ajVQYUFZmnNGsk1ZDP
zm0Im+JVwVju4095u+p3fgmveP2uVzdRTYszr7n21d0WtbYm1yQkC+RZWwQ0oaoryqEwUhz0TKHI
6WfciDvTe9fzbY5U0IRgs+JqlRZIhTrVMc1XTqnn7HZFLbNvxbua089FckCIViJd7jFSCtHQUZQG
xKtEs0aG880UDaKQ2czaVZzeQcNN+4B4nV2lp10z8UT+IE/ditruUPUdJbId7WLSY4iKiMGXjqXm
/MoV0q2W/z2VE1uZRRm5UXmRn7nPNn16TjSChqbFWr09jjY+FDxmYI9KfnJre3EHRHOojhG+N3ej
XIgFbMZNodxOSKe5/NSb0WCq/Y0HwbIoLhaXn7Goq1Xo2EEPPLohlLd53/VVnU+QnErzafCxRuGb
LNYwNRptQV/h/iXm4xC0fbXCbTN1uQvNZ0M0rkQzOwfqvJ/mIxSX9003uNwiHsv1GKO2ZT97OBlD
4UIbXIuz9Xz4Aq6w4v31vrsxWg9Ydzrkd1vBfixh38v/RPq5sbuL5G2jVtpbP6ZEKyctky9OLe86
I5lalROejZ2LlZ/xZIX3+UamEXSs1nq7+xglUSipFtyF2OvprCp+Gwfw9bLdPy1v8ZUYLpYlFf94
gfaB2zBot+is1Nm6cOhlyB4U69sy29xzeiZTigVmv4TEtLoPu3iSrfGM+gvpGHdb8+OD50Lq+Yu0
HU3qriWTYIQvq/Aiy/2CkUJF5M2ML5cFivh4l2io1x3IAZb4+Sx0resHGv6Nb4cnBQzZHyUT0Hvx
rMOx7D+aNg39o0Ef8QpNA1gZCQIevkWSYy/oeA0wG/jYrhts0/tOj+bq6UAbuOBkvIXfDRxrg+tp
9oCjOAVVwOwic69nP2lGPx3UBvJA1e7aejlhapPevFSM9vjvEntQ+hFXkidrSgbPxGsr6/LxOpCx
26WRLLMHELFPkxZqCVq+Mn1CpaABmuVtt9ylwKe6PhgYucR6UltvS1ilm85YMqUSBqQ7iVgrjzQ/
nSyyUl79a4dx3w/kiv8ggN/PnQ8OfAynNT0tqcvxVmQyIZV4kIx9pI9TWwHLgliu9lCBLJ7ibzh2
1a/5YICmfWW/r4SFFGJ6Gmhxis3EsqXi3NQ5o/zdgSVrKLIhKq2tuFFOUJwz/9K2gg3CM7SkrzbE
kO2wW6BPguLVy8U4Tt4Y9mDJbEacCoJxIiq5orcgTa/ho+XldxGKx33G6iZfEqmHesc2w3Ghko+T
4UmhvDXCKib1UjP39C/HASL0qPfuwpzu9Vv3SnQvtytz1P180Ighl2AWxUPrAL8q8gyqE4+xbe4y
x7a2BiqGoYn+S0oKxTyQp5otHMauI/+wqqjjtRbiHNUrDPhY9BPeaZ43cPR66nmISVO0WZiIuSmC
zY2ovaQvehHppiMR8FVyyJODJVc1/DDQRgSMSX3dkHMd53JpocCNB0RxQpSZWZiiKsl+wdZFkfIy
3XzqO6MsltTto8144eyVGE6HqM3kriNhRlFBZWzEDql8ns20P+JTVPXxYebZSqvyByh47/MTRnfn
8ayAc+hmV1TY9Pwsn5uGYFAdnZTKFfjFRHBP3KOOR+OfwdXzNe1rvvvtEWoA0o2qTxj9BHiUPCnF
ZkiBEomEBeqBYXs3oU1XUhK4L/5yXXVgJMoJ44ivXuQl12VyYxHI1Fgfe3eI9EOBuUGwPCUa6fIe
jNx+TIIw5Na+MnHDlXw5yMbyw3M+/RXqZ8CjnGgD2yqjH0zhbIcUr4hg9GaLcIujH4J8G88f3vYv
pneppTgwg6tXY9o2/7wZLMyD5GK0e/SMQIRXGCsQBxwYmu1Spy1cbtd3FbtOMZOsyRaEFb9LcdP5
GMpS5EVNo2sh8ZDNWMfDuH27qJ453VdPmWSleq4n5iHe+vOwGMDTO+lyg6PPkofKd5WcVxfYsuUH
c/ULUJIn9xSSiDNiUnGoJwONkvLxqaFWOylSnLSCyHN9ohOxroUy9NuWIwdvVxo7GJnbz38WXS84
Tt0c/9+JCSHfHQj9dmS2FCEv64kRkqGPEWlteCBRKMvrzikYYQ/+yksMJU0EbJ3PCk0lZ6Se0Y9X
MnpsyCzTdP8Qzobmbq7D+siPYSmNByumRkF8spVMR1Hbe2Fm1XTqVdsNGvuoIbfQKvi5xPhvmNGz
/x3A3DKe/gl1/QGkuZQhvGAPaj4jtolZ57gmi5F0FPaBd+Uzlm5F4D6Sbqvu0gnQdBi5IbELpG3s
Lu31f6P/QeWQ6Q61FvZJ6AoSm2HvNhmxT+9K9pCvcRY0VC4DHCGPPXyOufB8e6LIaHBh8HgyK6NJ
KLWqa5z1btz3ydyHvcwEN894mhhR5uC4b9zUAsvPl9FeYTpJvxH8mNwKBAd9z79M7VvhTcx4mVuI
EFoiSCmgdfZpgEhLR+WsVj3FZfIsh2TorDZav/g8ImxdXJWeTkLq5Tlun3KP9I39l0hDnj3VK7N/
fJeGePd39z5G/zS7okH5TvRde1Zs6cWIQ5K2hK3dsOC78At7sERx0tPGU98wo6TIaq7F1yWHBMVn
Tl7tApfxDgtsGGp4S/jlKGccqPE+Ta0R6d/9nS6Q2+tLM2q4OjaIwRZvKFDFHrTuG7F1Cev8tQTc
SsiyPr3tPn5eFdj9dpjZJAmktCLZTa+CHYk5MFDTAxfSaf4Ng4VQ3YK63zR5qBZzJxV7T8H1UHEw
PBSKRazMfY9RN66Z/2fxbQ+XgkTjNgd0trztn/QzhYW2ImwtPM/MZ78/EUirtCTUZwU+Vzs7KeNF
AYJ8Pa4338wVSFTow87lRu2hLw7oz9D54GMCVg4cokzbuVX9fJv3UAQZGmpiS6R5VlTz4JR86gzp
xiv0sQdI8OuNQkcwt9anRizz9awKTH/1WI+3ZeAqsu1XEBMgNyS+buUjpFuoy4pWyYnCNe1HAuPa
iR6PrR53WHs0/RvOJVr1hMedAMpgDSapgsX33PzWLy5P8hkTO/9QpM9cHzxLGZk7HNT3d3hICwS8
OnOo394a3ILBHuS0L6dav5GLAfnApZJkednrjhc4UDuPK13aJVeqre9+I9jJFziaCx69RcvgcLZS
p/8ZTKe9ouj1zhQY4z7lB8xKf3XBo+XzKjCAmlyIc5yvtceYxQ5XX89GNx1PmNUOxkD5EsKLKS2k
CF9RqxndhNbvooYVyS33R1XEHkw9OM7maGpjQ8tQfJNG/delqXcbYPDpplZTQ3AfTCGg8JQKGtzy
/ee++HaPsXUaZVoC491rASi/g4p8qxvfNT9UIiTEt6dqSd8mYbX71pBIP+5qguZ0IdGAhSKbPHKf
Sv7npPcnPiojXuor0vGfwnY4sr6TzRbIQ4xkP+L+0yw0mkTql8WhCnGIr9+hRJUucETbzJ0pr6hL
c3EsoUpzYPwSXPghg+1p4znR17j6UOYNpNpOMkus+bWnAR5Qa+rlzD3lsUeH8oQcH2lDo02NDNOg
FUEw3uwFVCs+E9uZ5+gGR59j5DNTKatc9/j06tDccOo9N2owNHmLtpTfqQ/5W7iVO9v9RI6JVSJn
uvyVRHZH7hnzu/iL7vbJ2/Q8PANDmw6aFauuEA8LBk+FiUgM7j+x/49DHeXHh1crfE3iCMrx76pV
1VDz4qU7dRsTWFbZYQmmNSqHvBNq/qXqvm9Hyf9+37tzD7YWWAh4OXm+36OPt7E7pEAjFzzD6vKU
/zJ+oLurryCO6hNVj7nM2nX+uyeHpkqEiJGEQ7w81qjkDZdOq23DpDqOBxIwRgi+IKKfHYB7uTov
Nhffoukq+wjz7rgAEUPYljtWtNtlS3SbhE7sxsY4t9ydyFznSXuEAPPvqCsUPm7oCqxD6dG0Vfru
xaTQrRN4rno25RHgYJmxJNcXHt8HG6dSAGM6gJr/l3+PoJdO7BkLDWL9v0Sfdx5aO+Co0SdPzw+C
+CTMg5rJEk+eA9QBA4UpteOgI1oP8MLRVeHzOtx2kQbmD3dphKONZ5qc31iKzHDua01IL/bb3U1n
B56I3JHZZqPNhaBEhK6gqMFs5Q76C/nKuBAN9MdlGDObIEMRTElkU7uiIU/hC1PCAYfkvynSzEqn
qh05ZzXXOEsk70U0Zb99xCKdoIlqk2zmKWBAVvt0ju9j3/VjesTv9lb+vKnIdxFXqFr3bcr5kcQQ
gC5dqCX0pnywp6Yv24JRPJTCQDXXENq+wzEWnfINPANDAcgu1QRHzp61O0m93k/6tdq7pZS+32Su
75BT7H3PdmnDx++qjQ+FhgJUe6+nfe10g36BheKtkWlK0ubX2aip9DnHKWVyqqKyxg8s0YctY9wq
qU7BJKwRTKbUfEP8V+onfsfLuC5SdmanFiK+V3kr6UqxKLOoO4uULXeNzuTYZI0dvopFroPwcilZ
uMS963jFRRr23bt5HTHjM9zMHOB9/rOIU3ujxANjeaVBz56rDY6tO3GelfL/W1kIAlvkK4nuv2qh
h0EOU93KL/ytY8gcAN5rMnCO9ZzJYeF9EGkGr9kfw4Z8lbKHRXawOeljn8WnmdG7j4f/kUX7KNOw
3h+TclSuBdF0Jjf+Vo5MkLiL+BvjMx8gHPdOGthRqNi9RPZmcgeKCXqiWyxpFW2IOoxNl6UtgZtL
5Sxn9Gk3B28QKRdi1WPOIhdzqCU/A3OzlMUsYSKWKPgfIFOjP64VOyH0vW9JnuR67BSgesCrUAz2
vjladuVyIEaPbdMfLIiIlKQRpeC2PkYLFJemgse0CuBfPPyMxRYpMCTK63OSc5d/KYRQ0zV6GmVV
1kA14IewBOOIRsh9GNLqif9sVylwFDYSKx3Vw+jGDjc4pgjDqCn9iryo0OpQso4YC3wXbgyg9xfT
RR3F7uBw0hxGdIrj4SmosB1CO7T8LuAPYHgl+qI2VVAQtHnyPVMcPcNgVXXz0qiV1C/1q+uPoQF2
xOu83Jv9lNRPXueC0YqxB9A6Btzi1pU/m349upu4HY4eNgSRDTPV1ySAAmSkGhbGSVQ96EQadMIT
JWCzr0qQNmT2Dsnu7tFBMJvnh88lJN/N118hWi/3I4kPMcQzq/vc8tpwb4et7i+tNe+pMbn+Ndac
FwfIRRJlMd07OCT7I3ndoGsxlau00Fzv5euEy095qqrmEXgX+w83OiZK0hBqbbCLL474ieuFnNqE
LAYZEtjyJLJeoIqbAcTfr93zQo01CdqilbZFQaDLAGhUCCjUC+HBU4xLJhHqOWuFZ/SErycPT8Nk
0yTw5qwJ8CCi/rf7lpbEUy2P9GARx12bC7pNJFoiB8qaMgRt8LfbQUiWp9/430MfdrQ8c0jemaRA
mxQcyreojRjWrjYjy6QwZ5W69+NjeJKk1f3svAsBpd6n1zhn8nQNMpN/7lDmSBO2veofQ6nG9hoR
fwd2oA2t/hC441lx5mu2eWPb9iNSyYOe/i8ny0MyZhgpJ50+BUPhAh+GR0tIjdVYnFL3hpu5ya21
YSkIVK19TkiaScK61ZgoM21EB0jc2i1j7BriVd5Dxx2y6vHepwnl3IhIaYgJPE1tLMbTJmAFcpeK
Oe1RcOJbwFBnRpBg4ncbhwK44r5tpkHmK7KqNJd3vWesMVWyQ9YwCEo9CUpycADhkWWT2T3V9BZm
DkiLJevdEcgh7UKiH/sZX6MexbDgY8QdQSXHPV2k7p753Y0NDEYSql+VxLCoD4iZPjNoGP5NQMHV
Yl32coDOjwt4JXd5IicfMcIY3byWaeWgdwxyPS9XHB9FFii2Hb4WVVKB5U0P1c4Fn+MsqCYgA46G
xDro+kj4aCTy/RVKsAQPFlWaXr/233UJ382DuQn0fF86ZEF4Ht1CxuZrEC+9Pqxq/0Gi4I3wBO9o
gkT2tJQooCqn2NF1LEMaw6IIn1ugSkVtG2wj/W4Wp/77Quu+8qtFTa/TWwfPseARB8+SxC1bwOaz
i+V9zwJJh8CtSu0rNMgnG9WUYDFG5tFskqDJdXnw+ZFHnd/SgnYEoOZXwbrh4sm9NnFQRgFO2n8s
58OVy1gWQLlu3xx1Vv02+ZFsM+7IwUIYXFZ73c96rLzUM/ojGCoIIjBWAdtCxNWy+Z0Uvy+BYeC8
Z8xsR59h0oStjY5dyO4mQA1hMT4zUlUNIvwqG0FVq57L8Relglsvh7yfxpzIHleHyhcZnKWza+21
qmpfLY4yY9MU1i9RtjXzHOt9a2ZwMZQ9/HKR8Qou+HSLYxbLxCHmpLtENwbWA3R7B3cn0M4GycGa
Sf6RuFsoJF/TVOEZueS5Deds9qlq2qBIGJQ12jbIBVKiJEw1Q0itMxHr9AB6GuUox2oIy1miBpKB
1bSPbUKWROQUcVnx+IvIlh4Uucai/g1hdSltNUwLFYt1YM+6Zte7sIBQw2FJ2GQWpRZdqagNJBCZ
VsnVKY1XuiX8w4YOuOL0fV2X1dYzsYEVKHt3xlI/OaRFCLvpCJk9TAXZGv6a0OmUlAdDDCu5Xa5c
5a0xtvtCWGNnvOxNaSlU5v6v9YGf2P4SNYLYvRDmGV3o3DSEdrpw94w4tuAMUOXE0GMBn+b+dhoN
YeBhUxyQMr2ppHQ+IUfZSxDYN9GvG++fkVSy8QYKck5D7LG7IQHKb7/zibiZcWQyfrNVMZ6P9IVY
lh4kRfRCTA2Yc12G0Wu0xooFeVpL6iSmv0gDIkjc2lYskx+VOwQLSHNcB/jKAQXmc0UkME8TWxbz
15pSEMtfPKVbpu1lPGth+aCZredBjrc7KGNm6UPCFiFTFF8lTorEt1NabWmDNOoL6DhvzltIPrN/
B8xW00kxqxKBW+jU1c8BoMrupLX9CpljYvahPNjwixws+T/6jsYMZgpr3pi1Amj99uWt22lIEXDF
ZKbu526cJ6dIyrlZ1Dkl82GGjb9t5qAHG/ljFvwkc7JqtJRnrCEArqrq/UGRYAymHVWvYFe7fq4w
yFzSAIR8bL/RV+kPODJ8PZ2d9izjvPvY0Pf/xSKzOPKjIS38x26+ob/JNN+Z+hafoQU7MG9AQAVH
YhXAYwlIczjQG/5tIzBRgVk1brtp9gVXOGHdqgPcyw+wWf6egt59DOxjZtxylk5c5LpvDugq3TGT
r1lUjg0fRqNoUbp4h1yHGMPrLOcge5tHsWwBkS49WSYljW3yXZShN6ne5xnpqBAziXJD1YX+Lo6M
IoY121AeRZUVLNdhM0Qyp7WcNnjyHMFQ9oH7pACouZUbCzjgCZHD4mp1Pz24LLJY8LO/vtxV4vlP
/L+TF+tocd2SjBcu6IUK3GUCuCQ5kHx+Iq871g299hMkqCYeuO29qauPqpX3tpobWg5F5CgwbXz1
ESYz9Mi51OcWy8k2EQJf0l2w1EU2hsQ6rVEyDvXMPjsEjHBH8ZpKHO02eeSGkxhXSi26mM8rYoz8
NQUzeG5Fjok1LxXvqLswDQ1I8D9mVHi6ir2o1lmj/kkcldWYy+ooVrh9KOUduJIOXAxc0qBH1f8v
PxC3GBjJCOPz+GPv9Sq6w38tzcENEKSa/mpCy3Ze/dWdvSpvaKdLCGN8NDZtqwu/4D6sen+AG28O
taj0fEwRuDPe+478H3RnpRM8wYNX9P5sV/ExwiDPkUeqvlZbioFIL2XO8QzdVh6bSjyeGaKcpOmf
RgQjIzn2c0uIxKGsmJKx6jiz0eKson3nLp3tvDfwkf2Yxfn8//kPFYQ2Ub8x6Nt2Bk2iuj6MhRjE
XxUXolHzJf8WF79jS3Rbm33HL0H/hP8eAwHsY5ry419JaNQ4yT5+llBQoLhqI0TpBvK/CkmPcJRg
uimOvlwC+OMM7zqiJ52uUrLwqKpcHY3F0B+AmfTvpNgqcF36HwWdBqHD6sKgDtUFIXgDPHVQ00h/
h/jaBnXCHqUFKdjSHjwaXd71KGaW204++5JBLkiw6B8C2Tw9d3L1ygmQwJbaZDpGtloBMfzf5PJR
AV0P+AdKZOn3FfEo9fkADmXBPt2f0PRfC8igjjcbN6hnYIAmmfD5aemB/n8yno29x0fuNN4x631Q
hru1Zg2byP2aa/iYNtEKu9YicF4Lb7shrq2Ob7ce4nQ8EDz0f1QH/aRcCzwOt8a2DLOX6CHk4uEE
t8dBkCRbEw0SX7844LZNOyM6juOxx8gCwRqi+NVKGjVjGWpEWJgA2q15vIu+GNafDTWeCh8nS2ZA
fq/Rbxas3+UiwEaR7xMuoc3xqMm3WBK1X+gDtd5Exu3A7IpuM5Z6krrccIpOVlqBhUDMX5yuuwak
cvfm2IbObAOU+mF1gXyeQNvy1iW1RYVQFMbDmwMZRnZM1SgZqlYRYjgjLXGR5O/rdIYh5d0PwFPE
pMhumVjt1zRvgtYeYgpPWAdxIRXBgXtMTO+7KcOA/0kNHczMneKz7PM/DiYVwfz469lhUY+qzTcP
K0WKO4GgfG4R53csF/QAi4E23HfIOXeIHwErqqUoySwGCXwN0o9G/KgJA9JC8LNOzarnixn8qhlo
+JYXRr1dJJj5umBpVJ30FS05wqVk+WpqT6fvp/PFyslcQXgOKn6ILwsktvfp4JO/DB7lIyLmJBIu
Vff3hKTGEbtztTrx6feroNxaMAFAGqwjy63aS+5kU9V9Rh8NJuGwpmsjM7R+HrwCcU0jH3W8gotR
oyp5ZqxGRqR2AaWQ21Egf6rOQ7zzFrLEKPJjROO1+OFzwWl2q95eHCqhde/WmJ5X4R372QJlYoj2
IiqYTrVZbei6yvHw23ihBC95V+CZ2yqlVR2aubyxwAixAoZW7RLvb+4QfhxpFdyorFqImvqoIrZa
OOyZg+xyQVcp3Hqo6ah3erCyXuZZdCAGMtsvwsIonb0v64xlbH0Pic7POlUdzDOPpEwi6RYeGq+P
hMmMn0NNoC0udnkmVzLqSoUYXAb4U7wq91kT5bvLN1tAyS3dlEwFpMefULABfzUlS/X8JTQME2UK
Way4tspa/ovCJk/Z9gRMf0E9ZM/Ljt3wTSxxueMWOrvI0FTRblb41QiLKiehNnuWxl9qGL+4asif
2bgdspDKD/J6k2XCVgOyQyB/mPtDiAqJHwIVAK+6foNpCLYtmBsJZ40bVfOCJilLp8BnDdlTrCKf
zzzcSXelZdYDNOc8QZF1v0rETJvGSUeKPmZFpbSGnnYaZBi94jB2XIIrWJEih+Z6BJNfCJ1eOID4
dRpSXVDqgFVWCOfhPvB60dVFnHE4626FfzO855NQ59rfEANuWeggZiGGRlOPFAGdhPe0LgYQ+GYa
nN2KMxajcQFFZ1CGRNd/BVYZXHTUcWwZXE43J0mUjfyT3LmoSw7eBIH3EnxBegXVnnRVTl/vFYBq
eSXVF0JWC/Zqlvd/zFDQY959V0afFxMcdMrUGlL02t4XqCSQsHxeKW+NHVjnLwDFJNmxAXpBSfjd
vY9Bd3uOrUeHfklvNIzJPGQ1uu7oZZeaqKyKXFxWCZ1I7YBBToRukM9j+GZ/gcGLP9dbau7T3Yhb
5RP4pWfX2PfTt0pwErPGxdORoeQtsoGi5+mkrCBAMUWylpKeiGuZWyvs4qOlOWq5or2efBM4i3sU
MZ7BAOpofn8BwYyY82OFY1RvMxY9ZJrc/UmPJSAMSOsug/GPdw4e8umDTJyPc8sHe9vZfYP8oXpi
/4qEMw8bGJypeDWAoJwjZUW6rfxT8klJYcxg5KedXBwt0BBUdFZT6qc0if469/KLDfYZMc6dQR8g
Gz244bVEu8TssPIlHHHafg6Ihojm6mxsYq0Oif7s2n2xaf/cceejnbuxIXICcL0ZKMiMLETjVRN8
SomkUIAx/dIRhd/N7HtXr5IDIiAJdBY+blI7bErocu524w0r+dU7lhO+izPBFIXRjE1jx3dFBg8V
rs3IQzcpwDYBX/IH5kY7e6UCYuhhTUO+znwL18tX964Txdj01ylYPIZywvB5D64rDFLOX09RWv0C
eQhUaK/roT3kjrXsdHPAiiG3axsv6Umtg1l/TQYpm02wMcJbm1gLkYeP/mYYPuCohZJcWt2f0xQ0
+rzIhrFDkCsHcb0cYkQB0apIlIwTAfkSXtmexeEcusySSMezFNm80LQisjX/+Hm168v2SAx4Y1gV
M6zRFQXR6T3zgPNtM+H4Ftru8f85EvudDcjI2iEHrGVAC3NNI1JXi90Is8LX9BLU7H8IhlTmiosW
Jcye2gXkoMwx8qEX4wBCPk3UJHOSI60bbh2gwIW8K5ozFTdTJoPjECDR4gwwiLE2Y/b7/VGqh+Rr
TzbxahYGHo4MLRbZwqP4ggilw/sj7Iue7qKgZMr9X2pJ1GbAAfDPBd0yCKuh36vCmDh+HlWkTprh
J2P37s5gaBMjc5meRX1b1rwm5lOBKjRKYFq90+IyQGtx3KNrzAYnRK2l1Q7PDVe8ov/XEvt3Aowf
OE1lSQCqjmn/+EjvfEMSNvOXUv1PJ4QK00AfmsuooX65luCrBcyXjZcOAFk/G+NoMzmG/Gvs897r
60TC6fWZtML08vjj7aoJ+01cwQU4xQQ3TQdLb8cLrBBVzDUstoprzxGpZCJg6078T9GZu6MQ/LzT
UwYGeBpQZuMIhcPUcbNBgdfoZP89zcxYu9/NunSIS9zuXbsSJ2gENreaI+ayPA0sGct0t5ezvlkI
5jUpieHWlvNr2CkT03wPUvL2TWkuTYOfPfAaFw577HbPGQ6CAd//RowTvRmUEm1cja3xseQqC1Qs
QxjotHcpghwQtgLr6x/AnieglGwbHzLA8IBjHxAIDfqzL/a9x2XsNMbrqqEETam5YZf69dj80Dca
xW1S7neTl8Dm0KjvAm5/yT7DMlz85PPlhrhfixhgXAzg34ulSY2YSQXKLFaVO7WCg5PZNhf2+XDl
aphHFhOnOzFZqN0NTQrQuwXO03tvqAM28ry9EXj2Tn3aaXtVWzlYh+3nZLea5+6j7zk1mI0v0iTW
PikOMFrxV5ojNLUPJDAx1ZQDjqWITW5wL/giBIiVCtdbr8Pqkth2uym5QAfcGdQYlgvbKPFu0rIq
6Zl/knvAK/Qy61JI0G7C8IHrKVGWxUDpdZ/prNPnXlsOyzXyL2TXI+MoBfexNQus2P4715SFNIT8
VK/i7vXULJ2TqofHCATKKDWdKzozzgVOB4wlH/B5rIOsQUhxmaV/yIFZu3LZzoFxXYPunLHWpQZU
pz8dOPBxi5mncvCoulTIchEyL6aBKoe265g+P8HGnFAZWbrLifq8Vf/X4jex80WcRdXp5dRJ3JQ8
U2c6XOpxitTjUfBKKm5TH87GOTXhIBX8uQ3vbsm9QHE5yKLJonCEeZgeyiwAyLd8qvEa64aFe8pE
9FTu1kL70joTOk+uNqg6rjRtLm6DjPLoo84CUsAw0MpaujUC8+7+pxt/pD2hwp4Qesvl8WJFuWP9
oFHPC4TBve4YKS95o7xXX0PovqS4q4oSYEdbwmtXPd6QZ+JATQGwrilpMrD0NHlT2dkq7LrK3j9N
yCHhjeFyBL3fwsKiUxSi4UEsXCCoQVrd/rwXdK1N7i/jZGGa8IG0yaGqTguaWBJbeHtg+qk5aiIu
qGRLITHsfCWjJ5i++2b4NABUs2U6HygcjZ5/cKwgVCu+D8a8FU6ZEW2JXa0oz9isYzr6V3lOhDjw
HhgtPLLdNgGg0/37QYYAV/9kKxux/ouVUQmB11twDrMd9vxjIvY2AsrpC0Z8aHT4kpJHni15y36D
+u9JAP101GMKTaKqpcvreX8CtY1wOpgowjOmqzgzyEWwMPYyPEgZwFxTs5K6fIp2f8rsnte2X5lR
6fhzDKcMcdSLReN0oQJ82imqGK9u0+IsfyPnLmojksNwVxXD/34LioJ6VfPsGmk5D5VXkxQZV8HA
EW5ewCzUjvF8Q9GQrCVfODj5RnNd8wdLPCFkifdHBqjC1p2FHw+/1VIr4kLd1LjFdV5tKZ3ZAOta
ajzKqO6fPuiy7vj4F26RpMRNC7nvBPW756IbkMYxziNZmnqyYNckaA7jmcHSQolDrJRZK1czq9KW
8gbF3elZUH0XyXTe7lcVD5+S7pzXkIfFbi1zQkU5MKvctoENKdfU6KnGaJC2mNaJIRxPBCkIt7fT
ol9wXXHe6rCBr6vD6EzRRGfGIXeqb5719mvMIKYJTYj8i1R9gj1j0egkEV+9n/HDufPjHIsmZDEY
siZnMReO7gfbexRwXFxSrpafPaPEU1P4xCQccVQjdTR+8zlegUx/kSYg065XHWbNIWX+bYJRIh7X
1NBdQCEx/BIIrvju2GBYAAJPYNUIJeHYzAGH73fLJyWfP77HmDcwOz9qci4XnI3Qd10/5kS11I2Y
c58uXEmsMxat7FVdYOvM+O8jfKVInjg8m4avDpuZ6CT8QVPA+gW9WpqoWOHVtSUjw9YJFLMNk874
0WFTheUj2SnZb1GYNtmysztTzYSP37Fe+Bsi0RHFlBIfppkm8DToxCOLreg2hqmZ9LI7N4/5gTGS
qJXx7dQMSHvRMecW9KdjYNW2wU42F4lctSfiFAzu3Q4gy/8But4RVeWTbSuwlzuoPtRDpKBbP5U4
rrQTWU5S1m3PGIsUJbL3llnx/jQLyD6Z6+GQBIw+xn9pYWW4DHoS2e8RATJFQcmLaov6bAOqs53S
u7fvTJ6ESvXTmFYpLm8xIsNNGUB2mhiihIsAQx0MwRkODXXMvh46Q564cSLzl0hVpv/NL4MwpuP9
epE/glzh5arKblO52yZ3TvTqV5ifMD1BY8oIhQBjXU+4I+HaZTn8Pt1ZPRIFgJT70UrFyWhPQfu4
U9BDRUvQWg63yg2oyUpZS5QtPAoa9iQYeojbDWSjji41IxNXbdF/wsS4CREKJy18BdunkFgsZkVA
wO4njACDNMC3CG6zg5IHSPr9Zyl3vyoJFOdFBt/eKru2OIbWemODhNH8QVRNPJlfdDngMoZJHQDe
URvUPgVOL2jNeh/9FA5iDkSlKtExlH4EYhoLk0s9TnHrLtfrW8rmP7vx1hnQZ3vCPBD7McZrQjBd
OarnTYqpBN9arFwyFVf9QIBp/mXmFDGA1s1IxpBH5O3JS2opBqIVGbduzms8ka37wxuaXEwk59sh
i9Buw43f0HkcbGZV2xj3P/iW96MvukBjkvfFO1zg8G/+U7GOmBnhXHTOb0cHsliRdY1ue+TNL8mI
dmFsGcXOdZzCKJ9SxDmKc2BDHtp2sZosV2+Ir9/K4wJ2j7MmZUlud6cwvq5w1zNz7OkYTbAfXVtt
lq5Pq4LNPhDXLD8XaQOF4eiFnAFAcpDRgnRpUb3tFeMX7to8pQ/O5sSou7++nbeUCDt+Y1EqqHUB
5BMmGdpd+Ilh94E1eWx9VlXH1YJfBgjHUPNuGIleZRaX4bl8g6jkwPbj4pI7njzjMEDY5o9dDPfX
CibcC8J+Mmf0rVrSEidqdrasY6FWWrkG87OqJsw9thzNyCOHNPbxu8y9xTmWVY7cETPYaQv+lMwn
ERd+q+058eqhCASa83zXvhOKojykshUCTTYOpTXZnSWOCWSfZyn10DdwfAdTxS0TkdYdyaadjLIk
O3VgDmqm3Hg22N4LfVR/fHa9mObfmUVNIm2nUVIENFk/rhBoLqx4HkJH+RcyXoGoVkmy1RBrO48k
Tr1A+IciPvzxk8W5PQe3CP2cfw44CEfffjKNKwp4Mme6KLXFDn0xJPDYbPjTQfX9J/NVcvDF/PVe
7qeF83dQNztlhndsNDQLPlkggb4v+kehQ4KS6KM2E9RWMRvhGHinus7/u6Sjk59kRnt0ejMEy6nI
rpABAylLPqhf5XyC1ffruuXUeew9tN3pq1QH2Oxg3Ha5B5TgTtf+OkyCW/uifVLUuhCtWisbnv4O
wpoLFxRx5JnrDtADzWeFdTGezHM1MQN/NPaOEnWkZViI0J0d07PfYlELrb8y3i5X4yE2ksTAw5Iy
FMwfQTPmXBWnYVd3qeMGyvdgilOwzaAOn2H78jNHl4SGPTWIvWO4JTL4SRhS6DkksVTOTNCyppRa
EnHEp/3nh6mCqMLjUjoigVp0vQcmg90aBhhCbWYwQ/I9T5hQljTyPFB5lo6/5XU58xeaVReYClYu
nbYEk1U/RRUSDqIXX5Do9zsmDQ2WoL1+fcygoZN+lw3pmbAkB8yMGRyXmXOydnnCR6K2+IFrdULy
sbUvm4bFuJB5aR6tygfELo4/Umybo+2aQSsCHpGhkMgL66Xbq9DPjJ3m6gVPV7zapZyBYDbcMNOE
rbgfIccBZYnmSKOt/f04ZPVNYTNwH/JZcPIbFvymEZuBpPk4V9tj2oRyyRpGkLX5gOGNWHVXBG17
gne7PIZtMKqVmlGAU04GgdbZgrG6xsGwAIcl4pyzGKZarY0cLvEejEVgy9m+4/BJRPfsAyqJ/B65
8ARfUk36zso9dQsJOHVeEeyAL4DmpielZz5mKFAP4dftsfT1Dhtu0EXZBCYyGl9ivKgbOQAN6Go9
gE4TNXOmtT/7CeL2yikeZKEyeWFt9PC9RAQMGAcaiPVqtNGMWXagwvELkPY3JWeiir92DrmHBWm5
oc4DRnp+rhnfJCfaSNeWW4b2b0MZmvh2IoTz6C4h2+Xnll9x/aJ4UtSvD1mjtS0oNrze/Pc/8/hf
SFopMdPwo4ZK0Y/hOOFQDb5f/nrLeQ+D9jILdVDOYksqQo2oEGtuz/rbUCcHCXc/iOFXDNDyI8xV
iTtWS0516YpBo/jM1CFG0slv+CvgC1m7sV2X2zEr4waFWAyk9fGZpWi+ijBW7jzi6jg+fjygyfYr
NGu8LRDoJ8cY4d+BdKBWrPLzLSB0jO+n7337Ue6LGYLmxu+MbcKSiDzyB0oLGDbFTMybBDg8pleE
JxNdXihOTM9OO4oYVuhl7ofcVozyuQ/VpAUuboJi6gNRUeT61XgLrKuN6VjesK92ADjZZn5LC0uf
slQrXLGjBF3gluZ+yUMbWpFSXaJ++CbHehjuMi2wFxkDL8MnawjCCw2VawcDHBDEM5z7LLhQZrpZ
aI4QZdKlHz2uuivSAX7LdiED1K2ormKTJE9F0lqgKHVbMBJ5eWhi9RXfcrqzYwUun/jkxzewlO5B
Zm+CP7RoxxHtYMyJNSf42ddBGJAbEaugIAjSxHiVek7lj5Sa1ukdVXnao/bMI+uMuXFm+ymbFZHv
cuuDaTHbolfbBX3GrVURcHWtHfDl8F1RCTgHe/A3wyXCLcYsxac7jQxPlrbdC4klTmchPjKC/ksl
rh+rXlmoLuwbzjJ7gl0W68hMDnOOOmP+vY/Ubx3fTNQW4jXBdFrFZD6ZBKf8uNpDClnSZlnK9zdK
+sFZ8d3cunyoEEDyU/lVTw5+XSNHrefWqGDQWkr2LNYaMcHPBC010XGDqRc5am1a5qsG0YsbtLax
t1NsIFzfbzARnz8/5JrkJZeHB8Ywhkyeh77gyPVREzLsHNcnDSCDlH+0GPql4rqqlRCkRAc+yiiz
RJQZZ02l3GQKSdoxDp1TxV2evxR+vKznJwLyrZBpV3/Y88DNcxy76Xp59a7q448wOrzlKVqeqn7K
MWPOcoTyhoZNJNXX0iPtjqN7/it9A3r+3Xbp5gzg5k49qPfbx5vuVmKcA5xpfGvSCT+N0yn1aqxa
+ciAt0VQt8TC9m5a7iNFXJgscJZg2Y0iL0KhwzhhZy9XYmoDJlmYdEuWiHf/VO0ZkVlrhsry1Dqk
Qhk73uijpFNNUiUyjjPp6lGfHA3dsR0e6dQxOfBF+9367b9oXDiwILe98CM11bmipUxu7cNUB+qR
IvDWyXGgoRf/UjXMIGqDYO4xiJtKEeVoIcYO3YkJbViLuPpCh0dSpuZAejhxYMlvLggfw8zPTCXX
LpUlZwcEwUl5wisRohPvKlLa2Dc9ndlPZBKObnJmejiWHJHyIZkOA3lILY0alL1uiTK4UZacvAdD
iYTDWxmzloYkanZzfycgmEPYGx5/6KXyFdP4qGnZtX1DhaDjef0d0vrlDYSzL/aLx7v//eECXoQ8
9y7NFSoqPKSGGTFDkLlWbiLiLpe9C4IpKDFfNll9ehlNkTbnD+4LoZncd0sYELFf1kn8ViF7yH7r
TYtLu1NRGOCN1DYPlJ6nB4iiOM5w8FOAQguerrHYgH4rvGZ32V3eJPFTMdXzr6J3Kd1kqApMo0+t
olbdnqKykfVHcvfdxB5dqikS276HygrCb2kvj/TX/2IlSH8+3FgsO662MJy00hOaGqVHilLvly7d
9uSH4uuu5mzm97TXKPTc+j+n7bcJ3qS4SbXy0IChMB2ktqGHYa0TDseJn0wSG/pFsqjro0j9AZrz
NUvjWIsnaIBx/AZJwQRfswbYrJsMS5Y1yOF97GOE+P0UuZxdo8n0UVYpaeYH0/qUAIY1BauEDcnN
xX0cpmIUa01wKIHfZ45dkDcf6H1d5gWkAwEsw48UF/cTzqscDWW3JYeo3GFnVuxbdv65+jjpUMdt
oJGLECCt/ayaXMfOy2YBJl1awwjK+SkHXUdhV6P/dKamhSsGOMVO4PILQQ29M8PTpBYYFEicDe2g
wdsbXk4ae+SBHIE1AX+y7NRu93FJb0YRGYWbJ9lTGe/3BOeB+7AAYiZntlOlbutsb/XILvWWAy1c
oVaKA2iJT4RmudFAcdWAVu3QWqQdNPvAQNRpNdjAnj0yFjxp/NyGP64KJqytcsZtirAsfmWyJ7P6
Vj8NUWjNCtJmZKsoNsBwlDMyEt3lWY1aSmYXs2NwXB43bDOSVTSH6H747fUJRwS6B+6M3haSnJFX
h5TsZCajvlkbJOQetkNhymQhY2o/pU8BtMs2W6vypvq1iL54oVWeoV3GH0WReZCArxJ0RuAQsL7f
DVf9rf7yGsko0H0fpaq12tbrhJ3g2TpsQsXUXyO5X553uUKspX20TzfZBwXC1UCu/U++CwYGicGy
FM1d+DbZQF2r7OWxX0kR0zTrie1pYXMsOzdtlXtVf4Yswz855Wx/4Gbn+XwphN2OxMVKskUDTWkE
mHjKp0FhYmAm09f1ik1692A9qqkuoyo3W+DwRstbDVihZqQ6ZhyAXAtRW9N0v/EG2ZPG7YAhjNzh
T8ogGNDmpoGl/nvi+SrcBQ+gd2lJKKWJP/ehP/yyR3Htd3UVVZ5nwgA117f3tZlbJ0QGn+LMruY9
MiBPRgRavXYxC3VC2GGWbiGJ2RPpI3aZgg5w9YWRBs2RMvVPZoSA6ai1oslq0+y+hznqXm2EbhWJ
DgmCKgqMX4i9SMexmV70bQ2hjKPZ/Yn7t5uWyXCrp4ZciEnuz4ctlCuzLaS0i+Yllx1SNP7GGyjn
tj/SB4IDJnET9N57T55foav2X/vw9UrATnvZ6uk4njwjHxAKE3GHyiYz3ILMa7/5d/OtgzbsVjrM
WHgtXsI3u6X1yz+lZSJM9okfcvBNBkVQr9+0wrZCFl272DkdzNn6cmlPvGHBpEqXAYAo+u8R7XW5
/UdmoS7gopUl8lcI4ym8qmr3as52MT9s1MyjzX1VSRdP6OrhTRxay/EcpknIgBhVOhP03Mfug63F
4ueV5X+YwR3RAgj+s04JduckKPFskgeu4ZEVxAl2LRQv6WOjg/dZPdWvyGl8RiBYdjlWvgKdLey1
38yFShc0cmE2kVMNeDBKjHxP1VVVndeGwEX8s60zoLMtLTFFUucmuV4qrHdUtMZxGicQ2oSeJgTZ
o6D/aVAWOyy+1bDJjiRCd66QuP0cSohGZMP0gkhD4AfsJX6AoGlqFLgotFV88EWJmIJhDDc+D0Fc
XFtitElXQqpzcEaE8UBtCHhXYUdVHVE3h7AD0O1bGQh7kFxhYgBIqUKrOsinQ/L5DAZj0tlNa+Ry
jPlOEdp6rysUGlSXAfBehUTDaBUAaVZSSpLgiz+ZjUE6k8OhN6Vt0qldzXAQDSbEP+8N5FHNRsE2
3RdHQMOOXiYwnovwcLNOdLyJATYDxgt3oGiqTjq3+QWKOfICRRuKeH1EyvdSfoSLyVzO20z42YXn
D8QCstImaVbZm6+4Myw0LORjloiRCGsvU33P8/dk5/MfDTdv8e/fweXH6A+XEVLOw3v/hiD1CRVg
sC7jxLy0BG5/bq2qQEpxUQZrS4HeFouKDZ+jQVy4/gHLKhK3K/BHBfak46OfGxddD4RdkhhdrqYd
mWtZdoSop+iuEemqqERqQCXsqEYSUtK+3JB9sR1atxBENqvtNXGWfG1Ie6EIo6bed8I7loQuV8PR
qJuyCqA/Fmd5gniiG25FM894w2zu0R1uM2bLt5lhlx2bsps+nhYQ4+fxdYjYHOVWFmEVVRGnJwJn
49IQnSAwTMTpF4VEgY8E4gwxx93lm9+bdw+8NMBtCL8Oorr0+7mezshKl17LwOpt/L7bAG2NjPU5
g+E4PdzopwAVmuCzsc2euBt5Cd7TrXN+u/Kybm72ba6FdRt0cKZB5BuP3/267W/rZM7Q09U0i4Lt
ZFicy6d7WJvZWyeKo0tk3v798qHCxqAR9DAD7qbXL3qe/FS9WrVas9bI4gPr1Laog9NEg5QzkXdu
EY4ycpKWTnO7kn8ReRn8lvOqkx6QaGeJzmJCopCPfsHcOGeql5ypjbmKoynTVGMLhZhyh2pXVTUN
YAlO88FrrD5GZiepPI7DG3amMql9ACO2IKf3rWUJ0VQO4U7UV4yTCanXLeRkMdIjILUqID8X7dgS
7ielJL9x1HAR3bCaLwPwIWvnr55P/RndqDHEATHP3F8DzZ0FrquH8bS8OHM7boKA9/m81zTEk/rB
2qRAPD6KRBmvKd9O62IJsVvki0BRJfCkmxXa0uMVRK+RcRvB885hGvzgv69ZKAsnM2memrRt2+eD
ljorHwP0VmahY/9xnMHk490pbba4y06KMfkVOlXiURnDiZUNmmuNHot62ctTS4oaBFtWEsTvjEBT
14Ow2hP9oJfXOzz4p3S2CY4aHCW8nDsvlUDq2vB7mR0fK2WEa9dV4ydnoAqVXiEMBcGfgxFB/sAt
oRDY8i2a/ZHV1YLCiWwqi2s3EOnM1zi7YoTlA7bbL41+s3F1fciruCCVJZXm723J5Qk1GDwsiLXq
+DppgPMeP/F4ETST5+ziq03RRNvnA8mdC4rfUDhi7LkOoO4lRzbwRKBvAgvXVcnDVF/du6y1cvip
upYgD0bShKMfibfCyOT65t69OpiUXq+buMmfTsGtGjjm5SY5A2eztBaTHQLlE/Qiv4uHNsPruVKr
vE64ynwGtPE81uKPlfoo8Ednpjt3uMwBlRdseOHllFbayLdylwN0HTR8YbGEH06TE264tXTaAejK
CsulThQLLW6wgj70f9/GukMsl1hjJ42XnNCB9EU4YKRrDYfDxwcsTAm/c+pJvuH7JzKS1QoXybjb
HWddYbPmnT65UfEaWN9JASJGu8tHAF5dRUb/MVQj/CIIRobJgaT3VTaV/3j/U4QV4MVcbEAMFbYh
1t4Ta5qQwgOYR/tz+VwW7lb/HIs5iKCB2Zc5DQtmfxaWtBvqok9SfPFktN8EtwF9IOdL4Y6Lfu2d
WW8MSf+UumiNzujWzk32zFhTYiQuQZKCnKaujusx2Y+fwTEo4YQPGdf6Pq/hCrRh4x2i9YBpNQuP
11D1U9nuJM44dPgRe8DzvDeIyEglZvnSeB+KPaRzXbXwX/nYTf4855SP+tOBZ1lytyw0nXvLqU4T
jSxSqa/uLHav/l54Fcl0xNABnbcvfrazGTS5C36OCNi9fRWoXTws5im9iWb23MiCWNpXoNYCFdmb
aGqvkyXTni3lFXeXlMCT+tFKlJiLIYlYk0zJNrUPC2nH5we4EjmJNdp7dTSl7uGFcslOzy9Ko8Iu
lgOR4CXe/ZgJaHoyj6d22RBTKbBtZ9FpL/EyeixS+PEnrzqpNfVFQZzdCJInr7Xf8Bn9/KE3/B5s
9y2jvM/Se7R2bQpoRArNWI/2J56vye6jPQ+m93K9gR+tFC/3xLlmXgiDy3Gf7Vj45uHZcqKbikPr
T3O7aLFV5bENeHzhr6Fq1jTxVb7587RF01wzfFgQPIUeuhP7bBuSha7dkV81EPaicqWPnQR60A/d
OGK3BJ9C7e5xNRyq8RRMrtTg36c7zdmaDNTWUslSZeHzbChD+HcU3ZAp3Emz1luUaCC7EaOt/mUr
uzYDjHn7a++5zVbVutQq7Z/x0g0xSmtbgrAM43vfGPPW432YeNwDFO58Oa5wsaLUHaCPXi4Wyybb
jfszxBdo1bo1SxjcM608Ah1xu6B0ZJYFpY+m6jqJRWPGuWCu7T0K1QTw6QwQkbestNR6m0IjAFzE
ilVtEV2AI9EoinuTekFaPZH6/ttbFehfN3qPQPMKtbw4gygOaYxeZnkeA8v8qB9ru2w4HBtF4xac
W1uObrx5ilzmb9M66lC4u/4cyehSiH7aKU3joFzAyks70Nw6KE+m59XbNwHYqsdUts0fsUKTEz0p
YXhcZGFgZAmPT35ux56+r+adkcrUiSjOnXc0oxSNnneSSgjZEOvjqtHU5q1BFg97ftFMWUjPoxWT
m1VYvQQdkm16O3fK3vaMBSiDn1Ct8ymipaw1daMQ/iAbfS8rDbQV35ewzETYnykh9nzraI6U+4un
znv5de1eW48ukDDu9CVNGmzqZ5C2dtOkND1zeTRuToY35VvGtXcdpNKuntgcjRYo6laGBl952yqc
weX5GO0By1N40SXf5dg03EOffTmz9T82H393Rd2TqvkpHzHhp9g1UjNmN5matGqW/sQKI5L8LnEU
vaGznl2mV4QvpFAPy7sep+20Ahh83NBQT2GBQgZrnBb+M5TgpWQgE+W1sAz+V6nHTa38SyFJxACO
3YCrzd7xTYvxXIqi6D+qWRcoyWPX19j4qljLyTrzzGTbnXwF0GoZ0fUQGVBELZCo6IFy5GtMWfoC
v4bUjOp2cmBcMmgqNBs3BNage0I4+lqmDJ59YMYeRee4xTGPeNTPHC/hW27egb+MrouLoVvSu7xn
DhsIZP/Zjh/LgbKQpejr6WpJmx0QhsTdg+lToheDjEylgptWHjvFLN3FYl+5BERkeX3tMMQUQFyR
2/Xs2TLfLSEZmOtXyIN5kO8Z3rJHkjsy7jISM5FHyNDcMmU6nTBaCQyEUHLbRzeWLgjM+zyRNl87
8TuI9k4F5uXq4Z0FKoHwc+wEBRdeIo0Er354qh9csf7L1vciir6ivMhyhoC0ONoMv2NEFInYaaYz
h2ybt6disC59sUR8a5sVilJcuipXoDMGY6JWqCqIL257Y7pthyvlYxOqDmGYm5qvPQQKWwfG0MNw
Gw99U7dlhp39ExbplBEj7AUlDMz5O9ttIiU5q4DSCEZpCL8JhggQLA70HvBBXkvfli+OeZEL0juI
5l2pcuU5gjsuqwieRCO8tgPRqUtoFIheB1rcEGkTv1QhOFLDD6xw3JHuVaL5a/iVOlguloXCGUXn
T0DPBGZwGMLazvRPXyoW4mMG/6SYZnShSbvFn6L6wL+A5x8xxbW0a6xdA0nL66z1lJ5bEjhxBuRg
+BhS5MjbBKkmXgYlA+mEEYHx1oEEeO8MuJ+T6zLY8EFzdhBuT/nwmwq5QProtzKF68VACJxRU9Io
WY7E4SfLWEM8+Cnj00tif5iFC4w03DO5lTeVwTvQ8nSTAjcPFa0ekLKgjSjXsG/8bBo7S1gPhsj5
MkjL91T+5+7rZ63Po4CuSvbXPHIhJ1UJuzrsA54O0XPBfwn8Dr+asr/e5bV+eg8gHqsgssIfWbt+
5eYjvvqBiiss3Q8d9qZzVnzP23OgJE/+AyHf/GSB8whkbvrq7oCFK+mA9fEXb8gKsv2w2Ig/7iM4
FjoVdjknHznhAGlZr4bdgqo29idAJwAoeSJZtiMTJQJsfdaO04eu1CazphxkYDRyRY2xLQM0UmwW
+D2XdW2tB3l5qc14cfxp4MSrHSSxR/wG11M8tvAM/TU8yHckn2LjvhaqAEcBaY9wfzxSzhGcVTyg
FkwNlkarmP90A0uI8UKLlHN+tCEAlqkY/bYucVEshyZDypTp/yCrCnQtpc5JWrgezxXU5F1Luaos
7DdToXhTGmexLatWMylhirlBKaa2Q+rrNyEtRj9oNNVYfDW8EgxQA1TVg5VQ0niVQHkvMuq63VvO
lYXHRmOuyxpakti7Tvx4pB4IGSB5A77xEa9V+H1KJGcSwGZb02FsBVLrSIVbsJLPTcA/uo/Ja10+
slAY42UD7u1MO7y+vOz6/miXMShgpUrzumzpUFvY1/SOrJhzpTw2xSTBuScRI46VoLdxUtSK2LdS
I95oUqD/23DUYK4FEPGcCHvP18dyMobYOeUyfYuDYmg7DCk1PmSEZFViOkp9hxbzGxNmtKYvQ9Mq
siAnPvIAohUh6pMmGLhJdR4beXPidlABbcghKUJxkjFt86lTloLBWe78q4eBMq2PaAEhQxPlb0ib
Tub8Ti9l0xjC9HCRqmXfxBwBp4fLT7y91HH6PIZCRz39zq6sl8/d1WMsGRpnBISSa63Ltmy/A/dM
JwO6Qih4F5z10vuLL2Kr88ml4O1W0TbMQh+Q4XBIR1LJ9GnKtw+Vhm8MMxBRDnfvWGLcNIhKdyCp
F9DBYkIHvGv1PmwELNXKXK605WfxfgvbmfEK3JPl84odoFPMmHRGGxhsviMpzbqxpAgaFygLeGrP
D6t87eYphyRp+2l/3GgO9Ivz/gH4yx6Sj5GgXB9x49hFbXob9olOZr8Vv2o36E34XJY3RRiyf6/L
J066I1o7M7XZe4LU3n27W0FEfQnljBAJDDx4VyR5dcu+UKcIbDzm+TtG6cz1GoCSdYOZXwXi5f2+
4ICM7qEqnwiUdZuNLI45B+A5lxP7fznublhyiIUdy6WvCvnHGEIMevkdZdlsjEUFggRPLQ65ka+j
6euoRcieeI2In/Cjc5T77O5J4MlkjpM++7IM59gBY73dEICeqIAhj8C08QQxeuV/A3JmYCYe1nQ8
G8hznhVSXOv4bWWvgOnXqTsvKEaPYiXsBWMVkjN3X6hEWgY8DOkLj8UOj5VY25S4EQlh7kVdTk2m
+C5pNdEMuFhxZy5hGQGyY6ap8ExxWhY4gpRqLONQXmMOlW9rktKnCelSmH2hipQUL1rg7USSYHft
WbPgIaIpKBQdrGngQrBYSAPpHUeb2mtqIgaZgRezObrQvbA4lgQjvCnuSM7t7hFjk7ZZGoILBEvY
M2kn6P2cDt2tLfksQo2ejUUsQgBsXCGMNHGC965vVzf2BYxzsL5vNE6cTf44lbIrpc8nxs0P67jx
1sLV4DjX7GeNzfCGYWmwxD/IQwytO8ocX82BTFKOOcXJgj3546pZhbbTk4Iy5Upv5NllZAXHkfRQ
zNRfE3fLrdahwKZXQ08Wk256BQ9DAjTgUvaAcLK22sCwH62glAuXbLZ3pm0lTHwaX3Hdg+A7NDh+
Y+zE9l0LBwELhDxUemLa7o0XA/RW9gAZS/Uu8judkMOpGXIjHFSe95eBTKky6VzhxJtecXTBZ4rk
suwNGIjUND6JkGo+EbH+d3DHQxbiYfHUYgtaoUT9+PLdJApxDqYZXWbt/YqtsPSas9Xs94G6HNC+
O3EU0qGyY135fzx70iyRx4FDPMDu3GBO5mXaJVxOhyIU8OI+Ave/gqRY8KqqH2lI8evLh1BB9AyC
MRaHTPKhqWGwvov2c+T/QfKxZgqoMiWn7EhH2uOWIbd+z2z407hat6Nqfzb48nHCzm4HaLzkijOp
0KBUPkKwIoHw5aAdZDT8CEIf3hwnG5n202ukLXiGjIHOdjiAtS9+DugFE6vKa5T4Q0E0oiKuqgek
W/LNCIAICAuO4R63Jmuj/gIZIw8i1ikvH3KekfKX/O6+6/MWN8rQOp3ZT70Rznhfs+oR4wJ9oj19
8fS8v5oHjfFN9O52scAM6+lhTVRg73jE5BZ1IrirNN3ZJvwtkmwUPkhTYP8terL/03RlHXr6wb5k
wz0gRwIW35fUZK81dkN5GtafcJD3po/TuJlDQBjhBusot9NxWR0a1PNYdQ8LeNmBhehHiYcSfrh1
5RifCnaUcw7O/1+XorNwHsFC4v/l2dvmGx6ZHESC4CeYBJNL+6ZM+idHN1NWxqla3yHrdYob+WfY
DVoD3VYu9pE3gjbZjweBbvrstWsG+qkQj2VkAzvcB97LOZNjKOnmXWkQSJ4BiC0urOYKMaMgSVJK
AzYJJe57s1B6CV0vSxbvBqz3SY0uqYfg+SZN07WiTZZ+sd6reI0gncUZAWIFF36BG/MRPL0cA+Vc
b3ed9hsi9x4IeRCd5DEEIHtqx1JILUT3skXbrwqUkMPaIPv1qiNovEqskuOnsn7pdWY8cCEYsQZI
FKW4p+SbRuruLZqmSjzW/pDRLq13jZc85ETxvhlie8vQYGp+C+Q5EGVhdgVEciaTsz1avRGzWJyD
lYDt2bATNj/+t+iv05W7S2w74RjrnA2QpKR57MCqdr5qYs0GuK6ruV7VIl/x3KuVJjn+fc+CLFHs
pMptueZbidbMMQY1cbEJISlWYW7qDgIONCFIbBAC62qCFPaJKzfj+OT9hZTurM3cTWbIC6am9JDL
Hh+5W1C8aVa5sFykFv72gVlVs4dLDlthHX1bShf7eWVdKYO9WGHBtHqcIqj3aVQQoiKyRpRvzHWF
JcWKACbbDDkl6EeiolxjZ4CaKspQ7guRyXnLeGin3A+/A+2uWiBJY828pOCXz+YBWea05V6xJ0nl
oQuqNzA281CY1hZQND8lzE88cNcT5XUa3EuKsrhKJrQGd7jevDjGgcPD1NGNdCChnFX9LB1bTx9U
fdGKRVsFJ5mo2Ur/orDXp79FF1ZWpP9oZ4wOyLQqFsqLhOQanvD7SFhgeNtVshGebX4PaaOBQlrU
zvX8bGf+FtxRgE/y69NFdfGo6nFCGEBSjfEAVRA3WjGbXwaHMnE+9eCl+xhthIAzYkkNOA3G7qVz
/IB0+SwN3zl4MWYbImKSIt/mcAo6OqUa0S+2VAnvDb5990QEE1kmBZyrRaWQxC/LSRhdQWbFv41O
cwwEIhbr5nFaYqChwOiX7zkNTC9zbOKoiX++ne3KUpRKxYHQ6wcKTJEMitdtJOddhAUd4XULYd5z
V66EhxPSuEohFmTsLpG2478PLOaehldGXhbptfiItOld8roY86mDhoOoFG4bsz/bM6WSk9GCO2sI
ewphyplLY87vddDfARyXWyVQbDNdU2vOSeb/5lyxUeuDm47sVi6IQBjMIoGu+bIwbsmMlX/iq6yj
PJs6TEk3QggQQfzrTFY/cTSoLwejVXHTyTs5iBON5K4H5NugAs241tjg8OsmGe0LD71tQ7Tdi5Ro
SYf1J508EaaJE6bVVrun6OsZlc2HQlZzUmZ43pdnYFeQF2iKJIDUf6SroEnbKbgZFOZzY1BJWxi8
ks60/WH7G2jznabXQ5ivq01jAa2KeW/NY8W/MkfL9ldUQqO6ANyom7uGSBskxRfZZceFQ/AZvzXW
ba45HyQBjl7pFzyuAE01CUNYy4g/8BKqlMUKJIxAS3Xc0UKGwgOSZWs8YCkNV7ERSLiq3tTuymJA
4EemVSrGNE/72ET6NJzqrDZC9jMfoBYLmhCYrUaKxmn1m3gDovabcd+ACO6Czx4JcqLObG3xV8EX
wiNzFhdPZrDa00Kzwz/XjirRbQU7A3q+q8PMKu9UO6OQhvrIlh5tvojgU0SIJ3DSiu2yXCCIE6Pe
KdAwC4+1owIhgvcja4ixU0jXDQ4YICAVfTfFrszDe2zcc1WTtbiSIUYlZIm3pboov0FkB6f9ObZr
t7UWt2RAp77Fmv2IUbfHURCuMawGAa0pwsbfW4p1jc95HSPdl74RoKeopMQyiQQsT6Rsw8BkEyrT
tccYCfkgtmKwl8b0g8um0z3fAP+URxukT/+6FbBqdteTTzWytbtWUkhJQi3lPyt+yP+ooX5UylA4
enPwcmYus5bKQlFt6Q6BAn0haLbYtpZca2GUpY72QiTwvsiGhBFoT5bDcPhvd+YGnIYLJxLbPoiP
d4vJvdm1ee/l0hrrPTHMKvovs72SuzNQSpF0CTD1gKYMwDihUbqULpMJ0oN808AP9RLr6rKoDClq
Kpc/ziQvARty69lD6NR5vhOWHGTL0NawWDxIliLYdVuVBkpaiK2tUOWAeDeiKxBwIWotk3WCOO/v
xdo5NwMLrF4OmgvQPp/RANtMpPaSL/0woZDNG9WCvUZqL0g0fmlWunYsMF5qK0SliJmZpbqVhDKn
aqjk1jySsSilYLxWz6VlRwEuSLQywjt8/LVE7gc/vO+s+cFZd751tsoAXGtfAvM5O5fIXnP8FGpu
xePiVkDvbAWv6sWl3w/T/nCx/FQFUQys/XxLnPH2R3C1qM2F7SXV0OELFniwvVl3HhlkIimi7imw
ahLTXw2FalUV1h/bbn/eakjDc8ksYAX677jVmwgTbidMrTpLcjLETdo+2S5B8lLn5QZxiT5OwiUj
3vKz5cWwA/qPIcyqT7NUyvARJ0k93DoQNdpbd5WmAm4+Olk8jHx0fM0KRbIY/fO386HL/UElEq52
3e3bsKM7n2WMwXxKIKmSZs9c7m/iX8Fq8XOdzTSrQVgFb8R5B/WK1+akEBxBkBLxoE2Y9MYNOxkd
93XcOQSL6Vv0LlwZJzX0cKIh1AtMk0He7y8Ihz9N8nAKqpMYsgVxSOMvwxwSR3Oz3Dsge9u5fQkb
MA8LAt759O458BqrVwgdIohiQUJMXRMJ3dFxVg2cuE+ilU76hpnUnD8QXuJmJucRmx52fzqqwmJ0
nfapZmE0vd3FrdAjar+6kPYym3T/ulkJxFm73mZa6PcfG6hyUi1dgeegtHCZgcFb8oS34wY44y7I
+8Rm7gOZzICYtb6ImMgWsGekab4QhMuO0b2vWdBa9fGOkfQLenDVBfrdPe4X5qItx8xp59092lpl
2+gEjUNT0VGy9rApyeMqSlv7/nW8aH8WgXCjcClPWgrPU+YikNl3Ex2hvfVD+D4A4Z1K+jBQKftG
9dV3vxfvJ6oSD4N/64pLfpwPlXmHVxR9m200pc09I5RuMEFs7t/SMnfIMkS8Ny50+Hg8ewzZUH4a
Bti/OwylKW3zCNpWJl2XX3AJx7zJ82tTh1xKs0mRbVsja/j8dJfmRrj2DpW8RKNFfQJnj8CgwfRn
AYjxSPdMGr2f+rlo5j0Lan1dFYWMr65I8gcnCvdogNwrDowKhQT7/Q1xZY2c1fwl/4PHhigMkrvL
PeaDlIiH8DjJBvnTWTcUstcUb+Wp94Mu+btgGL9vjWV/6k6b3ct42MFGAZ8DwgqenXF2A+Gpkbfu
RpxNip43cBvEKiN5CSD7AsQd5JF2vg9XTWU9K+VyuwgNMtVr0VxCbbLm3/gDxC6WaeAJnHO0VRvX
bow5gpmvW5bqfUamn92xP1UPVrAbg8vwMjEgzh3HJksypWslx4fTfDpf1cwTmLRgQcAacHZnzF4K
Ym12rqDhSB83UbtK3h9VF6Q3osT0oN3AxlI3AWHM7k+tKFfeE6BYrGnJ7puhfi0/dlgIqs2QA1XY
CWDIu952otv8TR1QAX8557OjBSIFnmaGz8X4UEKk8XM7k+8ZIOh2NkxbhaW7WZt4wPpGcLO4i+UQ
0IYq2U5CEQp9i4xFR+xptWc3wSZ8uo5d3N1z4XlByrKFWJvLHlw2bL49Au8MaF5+gGLlh2OQWT21
Njwgzv3AdN/mnmXoLN9EWsrndfHDnFB6iyFTy3rENJ9Er25p1BQ66748FEfbY9ZyKZ3r/Ty/ltZZ
aDChQG9gBugdxHEaVBEHrPqwgd3w1ECfes9ZwDLQOOFXniH8+yk1ipRvXmSXIqMD2FnC3yGcWDgj
7aYGp/U/oEaSlc+lhCmCSOn5jjKAR411XvkHOZuQjI6IxnVjKmnChuauQ500vIfVYzbEImlcj+Ka
o4TB/qqY+p1J90WqocVVL0iNP/td0E82D3L0PeDFMTVAcJRWufzotcQpXdE+AttazhzzM9rve7Yq
jYt0YUpkSQ4mVQEz05OanSZbEIPeNyCAPzTG0Lkqf7VUKCzaEPN4CdQgoNFYk/VC9aYD5jo0hoc8
j+ydg31Av7yagH9N67JNgRsVBPYzYb9IellfxJxgPv4wbKIMYSYaw529xc95fsw4mdlKHs/xFIAt
D/CNsFaS+a8BX7fgGJ0h+f616mwquoYdu/AuwTJRrN5MksI5aulXA94LjOe7Oup89OhXjM7PwugW
UWpCu48J62KoBOhWVOR063JjNu25TRmT1EwGSr4Viih3BNptQLNvjhOYa62y9Td8/oGYh3xfs/1T
S/KgZfABkJ7S9nV/X7tZePl9E6vayw+oy8aPT/VoyioILdDrv2tHCYZXHDyHeR2YcpdsHFX1ofyi
Y0dUGajMIHKCHyjdNhlhI3/GPMQT3sJVmQLF2hQoa8tNzhTaRbNhhSS44a8izPB4I9LaMB27OA8k
S1SvUXAWcZISIFcl8D7uTctl2xjRQb4po8QI01/VaNYfidp3JPkEjQ0I2tzMh6K/9vCAi9rQVRQj
p1QOXpsfgEcv5qrQTUEe93NQJ9U3d8Gp3eNEVQxOVXwik6DvKDrUbcmcyfem4nMH1T+sn9gXcexm
en2DxoRNPN8KiH6RRHUt7W5rKRQVMb2NYzEGSI7QDOuNhOmyGR3IERevkSnAFYSX6GTvsAaOELv3
EvpyD/GolDHRsZmW4qfArF8j3XhVITxe6x5IwMSZ67tZQ/3ROKv5nRQgKpFOYLCJjZnXjdM3zkqn
jIql3hVSLgopyVBV71tuw0ZYngPNsBEB8Qj+20t32X7g+GcOFjdKObXUwPslpTK+kqoy3coDjY8r
QNnAASqkReYzxEXsTbSCMQtBzWV8UUguMoRcL0OR9KMJq56jHYJZ94rCRcsCubLkfFT8UZYaFTak
EmJ98jbD9qi75ueGFYrR9pnb4/03j0EVEM9GzSjrhyQcXVe8XiqSdcPJHt+hjZIFWigiU9uEUjjU
LcCo3/v0YTFwYPV6bO2/Mi/TinjNs5u2BDaHOhE3tkbdhseuNfygqBYjGYFYfAnYBoNFWppNop8/
WXx2afZ6yuHveFh9EJ99fQz/HNPL1MIbVoi/1mm/ACdjWHq2YvVERylagK8KenM2B7g7ANcELRe8
FAD5fXAqzD1TNzThSPZbB3l1ENMTGq8j7YA1gbsKTmO4rfA3NfH900g+DtMssT9p+jyrS+7T+7F6
fZDKib6NUnCbY1h0cIHA+5a/kGpjmKCTrpuj6sapuqIByo6ObBfcYz3Vv0iBvJIdwMBk2sGsdNpY
cOJXeQB81Ww2ZvRNKtsSwmE01dPiwuPp4xuUD4TH7dM6xNGf39UwSl8YXacBgQ5U7z74zSs+lgNc
zFiTLTiaAVIIvNtow2RrdMKE715lUGwPvHdIBnhb3acj8NKmRhuVz2yIBp5xci446xwmWQEA3Aqy
Wm0h5AI5pj8bORnrwWJhjHkdqAPYYBT4F0thGONjGMRdAN7LK97WhtPi52xfVTGfUNDgR6vycmd5
ZjZVOzwxpiE4gxt0tcHOYc4Xp5460BKBG0ZSnW6OQb+JT4iNqQBmGZB4DHZuyqpeItqerlfkJUnW
T1CkRbmuSMIQ268unfvPXExwtZ/D83AMKs5MjzDwMe+6OfUlVhh9xIIdD6kYHOpPw2vMXV2VfEJA
UbEc1T/voLaw0gey/bkO2ZLWt3dxeDYL5wGwYt0AYJfUXBf3DWBwIgrXKPMlMScXtqUwjLJc8ptB
RgtuRvR8Eulf6kly6Mr+yK/10Cx3P4+wcGAS25G73PuYBhQrYG4+gT4u1NO4Fh0G5Dlb2SjUCKz/
HgxM5sl7hgVYS/FhWYpKCRSVmPhtwifaAgmrGzBSFzHAJU+keFlWkVK/Jwa09q24TLqZR+coMqdz
/5zHOmMDNETCRJwnDf7Rx7ygDbklL9UOcbRF/cg/tswnFLNO3ayO3YDMAQG0qr0a8Prsj5X27ZT9
qvjAXPLQWu91sLghYWNGPrw5ifXmRR7qKtpnpY8L/08QPRyfGaHiUxriNu3s8wwhKdC0jVdw3SdG
Gmmh19QhZBt7fAew+7AZ9zcfKxUoVEHqCdBgJFgs0HylrGaceKOvuGIO8H5wD7yhqv9PQpFnhagB
RniF8wBp0QNZl9Z5ufqeoyMCtt7fLW/C2BuBv2bGUlD0hN6UgnLLuTFFvieMazX1GMXqugQnE6op
i/vzm1z9bTnaTS6k/fFy4qVQ8z/kbk1l3qJt6ppfNQ5fXx/sOhBhPoOaKfn7v7HxEXIpdCrE6pOG
wNPJJmU4YorXmg9JB44xPLlFAa2rhXb3ady4NxzPd0WNPI9SktttTfIetC54CfoHPP48LlCOf0+o
kANCVXjY233MxgQPdmL3u/MUudLH0Q3ekFcYWubbwsYlJ2gtI4M+TEgxrFYxDWeh9btvAVZFYUfD
jca2VD9A89bnG84IY0GFEM2LsubnN4vaR1NTOshShxv7ssdrzPzswMAsvaSzkkzkvpAH4LOqRJym
o2y1RGA5CvX2lOEVKXHo24qb6pan6L9JJ4n5W2oiDbDgKlxnFWScv/L/W1GFBLlexsKWnHKOIxYw
gucb1sgVWT8slEc8abbVF1Xb+0j4hfI32TskhevQok/5om6ME+YIwYz5mvKiWzX8iDWx6mvApqp0
q0LNVMYYwfGNHPz2jZJcGPWsO/b5ydv38JqGopsLLbxp8z9VSY43u503caAikiubPKZfot9Tb+H0
SxTc8zpw2jkMpVHrsdilehQ+/tbh72U0LNbURqLGm2LY92Rp3UrDs8Vbq3t6claMNrSLfE9FrWGD
cWThVmlpw8hlHxEaaMl1XUQgTzDjuPXxHapLAjL9P771aQlmtneeh3xbROGgc/ZlIXPBDEhS7dr0
kZOM1azcDmSKfDLktQvV3hFlX1MLORbC4MEgXsBWhj1MsA4DVUIEoXCmK+I3nhZSUoBCg3S9zpOH
SUBT0K1/Tc4q+29uigzc9EgtHFRKjUqzobGeFvZq+TkwBGE5q4FGkGU0iYFBXazFFmWspT313Zyj
lBKqm0n/ni4FrZ6KRmQet0zF+whA9UjKrv4p0OqukXtIjhOcKWVUJWgjP3edkagpUMfD9aaqDKTL
fZ+4cJ9+VDZkrF8K7U/n0pms5uPanQs0mMt/aKdbaSEuYq+C4845AbSXSD+gFqyn4n3Fm3098tAQ
ewHO7CxZeQWf6ykwUX0SF2d89KaKaXajtM/059dNGzDXvrpchbY00V2MCoenyuX883odUXUgmiEC
RG9T3U56VLG73gpJmhLJQ5CyxUQWbWkt9cHCeWil1rnPIfGSfCdbfppLstElwYVQmejoBnLlhA1Q
H/cYS9/WhCGmhagjWBlRbxUwpAs1xSWQfNTDZDDg4FTnxayIlinEzejw1HFAglUhoyvIgfycm12Q
6HwuUL9tQCTfQI4y6k+3qsJPMmP/uj4GtqZ2fMmqHxiclrPjeD9xhqYONWjCMiWa4gBHjuxjnigs
igkR6vAtIemeTmrNQRB0Z4tj7FceDF2gTyUwRDVXCNb/FOofDxAvfv9k3GuBS1bQulFFZaPtsqNH
s3VE7luRJ3KxINMsME7+GnlAbea1AVrfE8a2ERHCn4tA9u1T++75HCpltovoS24b3C9R2Hf51/YW
Cb9OGkVWIlQ3qRZHsMJWIFOBocIAI7cV9Ko8U7W/UldqlX8QTRonP6vvd4LfV8FRdtDMCqXg4bhm
HFy86PAtRwX43S/cXf3T6sdlNo4HF97iDstsCMuDACV7ilecA93GZnuaR7f8Z1sfx58J86Y8POuF
fvi0w5OBtrKcwvnqEONXT4hTV7GAagA+waX1xrJ+AUsz9TY+OxhpLxGVR+lRyP1wgDr6ZrIuz94x
TfrwcpEDiVWhZYDrrZhc09OaYkJ9JsIuChzB0FBqVvtKbFWIjGUmpgZZ0rppFt7W2BIzyCTbqiPt
7AEk6MS5QqqNCmz+CZVHfeGqXymYJjfGAD8CH0Rot3NkU2lbMob3ztLxmj+1++VDhooMEdUHWc5G
to7lwiMAWew7Y7CTnG6ggjxgZ+xygN3AtQJ2WLEpjLi3SlZbpwJiCKIqKoXrmj6H2wSuK90MLB8K
I+YyvLb9FXrye4TF6bsqZrXPC9VImsAnaOKGKrLITPTAvXqMezzOAVIQPSdd9O3/Qk7QPjwC7GoE
UqqYOc8jokIDMiQFKoowtszVigCwflosJfiVAtQEe12z6Wt/ULORaaixCoErxIE9Ig1Ej2EX6RuV
NyvOLmFgfG6hk0G/j3fSGxv9Drx7qBWdNmWBqFjOlrC/nQZF+/uxIuOBQLQgVadUBr/tsTDDkVZj
F3HCa2Skk9OCDDZPMptmS4SkhLnZQL4w4NUvGqKOHYkp7SOgJ7rXoHxQLjJwJ/A2jDAvHqIvHpvk
X5eKvQtpxnsCf9sLY1zdTmSonBbjWmW+8V8oHDcCeGeW2WI63s8wgTIw/VmJTeYQ4tKhqGWg+UtH
aO/KJtbRCHk6VwOhpv5wuSU3L5Y75h9Rgyy0bdLo/O3p2bL2nDoZ/MYR7Lkiwg9UvWy0tmsvhtBU
c3oMuA+Kr6ulA719ZLNj89pZ37Hmh/uLlAlDdBp1w3yP9fZ2glzf3IqhD7OlqdiCZ47o1rLMb+36
ZaKQO5jB231jRKzJZ4HgukSF1tcnpKtyGn5dgga9DSffaOiw3jTbxEPArazEMnURGw74KkCBlPG2
T7rmgybxl5z7iSTYBUZwgXFg5L8beBv6KoFQ2J5XyPK57m6ntOVcgKkjmYPmWbg0BCPUxLN9ewxG
r2QGTGW11rgRI9pwumz/3tkmqe+bnJSgsRIUm66sgp6UB2aJMcqTgzInhBRmej4qjHamFj15kuJo
ljVtO0uEp2aYrizLh1ATvudi/40jxRJxQ34k37LkRkK6lWyp6MaCb/WBdwxUSI3X6M3BTKO0/1Uy
Tgo3Nft9kwQeel6psCSFVP39rO33ioFiVRKr107eDaS47QfZKYVedr8326Z9kRtR74IXUO3gqzIr
RwagsSacB4D6YmbqENLDEP9PDyFg4E2JWfsImbNvV0Rtz+BuPnFQXpiM4qdO1NUKL3iCpfuMq8hr
YbLl4TJmav38/TnqTT1XQG9iWLSOaA56szApK4c6k0UMlI56aM11UUj7itnI6rMQcQKWh294a7tF
jczevHIxP8bt0H4COlVJHwG5jZ3jHTHU9wgE8fD3FNDwa54fGiMjlFxvv6NhjpqzJ61DXKR8gTTr
IpbJJLFL7NQ4X6PNDkS40Yyfk2HGzdWQvNdlLSzA/2d3KE6VfWPSNNOGjVzKEQYV1VTbt9c+sVE0
UT683yPPPcYx7TmDHdLbocMspjQumPCFC4DYk1pZARPfXGiOhE1zfRAA2jFOhIz6mzesHTDkvD6Z
Ytj7uKS95lWWCyl7ZrmwOaO63VfP7A/4iRm8LTODis6j0zw5EDMU+ZHIo6Y4azIlk4QxiivI+EES
2AV4QJPZuTBO0nKQqmlaSG4XhmhJE7OgrIjIV9weeNIqlf9c7CwHYGQJTWRYOuCWOtcQk97nZVLr
IuijfUMT6UKB9BPz2txSq4G10+a3GAhEXCYe9EZA1qLiGz9GxB7PIfVdkihefZiLyljHCRAf0pO+
9llXSJrvfgyBc32NE8zvOgsC7gTi7vo/lF62tqM57aS6pZZGtmPH5xokIvRnG0WXCY65R/f2VCsi
HVYanFelRfH4uq2PO4GC9q3CMl+Pj9IWCk5zTJ+V8TIayDK8mtPWQ3E5l/DD0hhZGDdin2sBv/k9
zxQOzBnMrHLV45kRRctcHl4ZTx0p0jOp6CWIv7XxwP29DK67sk4GxFx1VlsXoQTT48V9gWO4ZhPj
gtt7WuckpVgaOKmeEWa/Ccb0BFkKojcIMr5fxASnlkGn6Ry9jGuMC88RjSgqQYSvM0tY7TgRCPK2
uVZjqjgdUoIki/DeZtklHv1jhltBgDJ9Y4WeFray6yZ2n2+ntWfLoYrwV5OAyXj7Oekv09z8Yu2h
VGuKuMps8kzrdvPsc1bQv/V1uO/XX3DnwFXJxYy/Cd98FzBI/bPXDL7Ct1+Pv09DdNoh0Lnd4rOa
AKT1QEu/k7WnQQlxmd/S2luTtuLCoUII4TW4ugZX7VT14lG8NtbYVAbMQ9o6t+7AWPGFwRBvNSRw
j1HnLR36lpr3ZLH3PvDztX3BlIYR9QO44sQbdjYwfEsdkx0g/0RMwAreGnIjJfaAiu366a8B1lQf
HaGMAogl5ilqSMofSonS7HkRN5NqQrAG/wuZ8C9GrLN1QnES61kDT4xZ8XZF7EBGhhFkrZyXh3w3
ovi5LDf4pQZRgHTBCVf0YHFL+vs3RYcHqK6uW9E1Wwme0IoVk2HX1YuPEbl3TsMsBxS52MvFAqYE
jEt+tQkfWR8lw9mTaJG6FQ5guhvagLWW20suon7bfOWIB9kJdgMlE7cfgbkgvO2wRpuGSNiTR0gs
4A/qqRHNfYusHzrpbX5PK8kOO1cYda22B3Xw+unPpfxRLCMpdk4BpcofMnPrGS/ODCiA6dcmsmuE
yz/DCFq1FvUelanLoswquNnHrruoHqZZ0+BmRKcsh2zsS98nVlzlKvEQVJfgGf9cLEFI5JIZKG6W
wrcZGO5WhKk2W65vPAzD8ppAANl+B+7ip/3koOlJ/0Zg3vBnP4tkDrZbeg5nknEr1vKNH9zs1SIu
f0lqeQadhNvLmwdf3h/uLPGJ3V2PAG/JQxl3RhOgvqr6eeH3Jvem7qHdtnQBuZwbxnUcADw3PBTH
y4uctTnPuM7JOxu+3lRtcJnp6wt/nPZ8Lg/UpALNTODtcVU1IvNIoHWUUjNfJuibRTzTNPi7hb4H
adp+BgBBxqqegAmCKIyZkPlMtBly9iyxdrIUoCbpQfPaoChQ+DCY5ZzSxJCHohQNbhIaFZ4U1N20
hl13MAnQpoWa0JHsY2PxRgwNea5xthlTj5fWOza5BdBRzbYS7nwsBa2LhJL8wih+NsmqZXJdODM+
DiOvwuDCE/NZdbeivE0jeRpzGnQXhaSdy2yZI9KgAPHWOVdi25t6xb6msS5wkD2joJ7TuWXdg3Cn
yKxsEwz1svs1MTmud++TWavmPYR1xmhj1T8llbOu+9qrcoD3jYhhEugort8dwSnkakfo9xrjU7LX
PP5Y7HhywySuMhDDhIeS8zfL9PgfUCs94gJpNnKpIEtPGBi902KFlioR8xvv/4Mwp91GUd2/cyvc
FTiBVpTlSOxLnhQsbbVp1n3ePR49ZaXjazWlHaf4eS0ZnC+jwPdse1eegCTjRivJO6f1dfbyGm4y
rl4TQR77pskzaRGw67iVod/xbpfBUl+UIaneof64lxhYcMilLqT40Xx05dQOPTmtYUog44MobmHY
o8e2h8VGPpmm4q1AAnxn7n/uJRa0ksHYT43nGvx6RrU1goA+H5dZjXM202hJ7ZclWY7JvsOlAyXG
j0sNVKUeeQUIVNW/TeHJHOtk2Qg8eXD25TJJcUot/jEhUx8rbYVqO8dGof2SVJ6Z+WIn92qkWpBv
rjqXKkNytkepI12fUDzRtY1EKJsCGijY59bORUSObGgDhCdWFsUpuE9JARwPhSKTRrYXJi+ogjae
uDSC/AkPJE1gdoaE8S+3WuxJRSpaTzoPqjZMDUVfiM+NXri+n+6CX0LOV+iSfoyFbB/zY3EiHiuw
gXiIJ+2L4a/VuoQFX8nF6b21P7yMbceP8eW/swaBMw+117a2XO/Dliv3pCiZb3tvCc2D8uwoY6pO
UJ8mo/JMKqpgviAZFC+bDdQvHmBDPy1QGjzduDtX11RmJhf8lMGe156bNExAD4n1TBaFXTj4G8d2
WA6U+GnfUEyNqbPBA0NlSL77hLKC40NcT22dK/tjaIVq78EnwpkXpHRl9SGbRJWOtrCA5+JBVcS0
K53842gENIvxkrfbaRfNo1CkALHPyIuHjsYKR+ikSgfRtThILVGwaP03CiczaBJilwcLakvGR7o6
1EnXyn3sVeeoiuOfKazUi1/hwWRRWJEBUQUtyCpUxuHOtat12GXDzwSfZn35rtz0KmFC7artA0sK
vpJHmQU05Hq3E1Dp5J9wGLPp8mUtGZ1mU0WkJ6NPB4Luu3U/FfAgOHBEBwsMIh4Vf6kzNZ7RwyyB
2HKQB+s4ZuMkeXVJ2zW6RtQm4A83rT4dlyDkHmb5O73xiYGw7P5xeUBEojhDwOuvbS9ZmGrEcoUa
yvnzV2iW2wYTfz6fdyxMzh9drzqOUjWJj2oPyCRDBI3Bl0yQSGVBnbS+c6PhT5CtuMBDyGUdaL+I
yjzksOpkqKweo2dQln/7Tkc+KRv/qIyolG8fwICIT/ritGBoaI1rtrQZPaIkJ9DIruf78Dd4tdo+
ZIyEsydLZv48YZpRzdKWBwKaz112wT3VCP7M/rmGkD/rFmxmu7cUjWGCmYvUIMHKLYmWk73FuD6v
dWJ04FqvBHrldiSRBZLS39zCtZgHtPlkfZ2WDXvJLImLVkZMDYOSHL1gxrfPczLd3Kr+ifFHTQs8
99wC/0DfgpWaPYfn5N9OGuEMZ8u6dNd+dHJRdGLLzWkyNdJuRdIJ86Ez0avaXCkJFBHpdptOtIHr
yOgV9AGCQZXUE3PvVclVL90stZcjCtLGtbji3nOvttZo4YNKOcYz/HjBihc0Q/Ray5KTZ9GjZahb
Vf0DhPpL4fOGtwAP3dbeW3kfTd3HrE2hZFsPCLjjb6Sj2Kap9r46de92OClAtfOv2RulKe+UZBuq
s3Kwx2yyF+XnCqD+MYh1RPNy9U2T++GBC51D7AyIsbQxG1KAZxXH4ao1XLtYrt58Vfc9WqTYu4og
eat13MtWFMq/HOOOw48PqYDqovR9+4IeXSChd2KR2QBRq0mjR9P6Hto+mGl4VOel7T8AfCMJHmvH
c+jiciR2Q33lQIxdOCQh1hbn911ZzQjtpCP8Gyi8xAi6QMsAw13ry/NhrkmQ2gelXVYGcMiLe0DM
QF/f/3ncI5goneIIPYYYzs5x4s5AcRymbFtxHsJ2DpjzUfLjKfL2Uxb0YE1s5PIB0lWj4F/SCvAC
9dMUbrfC279cGPR5S2b0FFz6i1QtPUI7/wrI1ckvUrsja5Xfj5tQyP3YkUAd0U7UXRYg6lX8jLqF
1SX8jE7/XZhU2H9zLV3LSBFc+0nAfDsdFY33zOJqbqn/022IfqBSvLD1KJzkun+V8V5MfF9AXTZi
idj10IVBysXV/L/c9wJKd4aSIa4znpXS1QGQYWaw9JJRIEB0FhTB5BnWAuKZgE2nebrO9lQlOV6w
Bupue+vb6r+8lClmen6ux4f0KrKI80CLb1mslD5QbdvYrESw4OVjGMPPGTxJboVORFuXNF4eJm4/
QL9YbEWj+SBzbRkyLrMKJ1cDbh8/Gn11kYpFolbIjdv9h/KDPGTN3Aa+sm3fp+Fj4SiT3blYMrCV
wDPBqBg1x481Funu94dsVwQLZNNN7tVVj/qNHRKit0tdRPtKwhppknldrkBEafsMnBmTO9oMjphN
kvmQjvb9HUVhb1ZSwsEK3jVA6fj+IGUziJOhEQIn0VtWO6xZv6U/golJAp+zmX4sQg0EAbqDQWen
q6xDfw5eiWBzzvFdG3uOiWBconwm7mPhShtryTlqNUVcVawhAjEjs8X7oDWSvEXlJcY7ObQNUGg3
HPCX0JHM/oO6juqkRmemLN2pcqSODMkkxyi400UI9NdQ+p21+ffN+4R+A5eH6M3X9GkvhEZlG/Pe
76E0cwmQETGahB9mtKjO8EVe/+c6wcV4idZDXaFXn9xCgAiMMMXIrbM+cERKU8qXcObF5pv3BG98
qfxiR0fcKnUcCsZ9mxrK6NjGe8wIL4x2gBgD/w3WuDJUmVz4V55+OZDDVvv/LXwUbUVPkAJ5EaRJ
UH0v5GOcHyg5Wh1s3nW8yZv7SGfgas8B2ktAUEVvJNVsevx0tSE10tpJGgrsvFUoc2/IJlZQVoPD
pfpwPgCChCKBhrkHmmwEwvFAAgrpGLb0KDYEhOlyMofrRWQd68czzrbyTzkxGeeQvvIrbUru1jQL
U/gQ6p5CWP01qk+vYLzrpUpCO2YvIrihd+Jliio1Xn0Muw0oyWsi2qyPeH0g4qIdpt5bgWWON1hm
aScC8qqPjnpyAinCrBsZbZp9SNNjp5it68Z5diItaEBfydH0ZwgLizdWro0HvOP9UoWHiefJOxwg
lzKtUyS3aCAOWc7LnEbeieXSTc87XRiNnjq4N8hBcSZjq99i3cYOFmQeT+Ln5wNihN88BVJyO7F9
nJALElvshkL0ojg9lWaMRgiIZT6EeOO7rFTsltBurqw0O2JckrGxR1KxNNuCZQ5tIZmc+o7Zl69B
sAdOMxq8x7n0nvcFzdXJPu0JF2JgvCRih7i3RIJfj9r5nSOQKxmKTzd4/SPPGc+lR8sO6za8zkmQ
ReNQ2papdHLUAerBh6stwnwC87kOU0kMbR0yyHZu/uOw4vs/vYvOYAgkAqo08ERfBY9afg82qdiG
kyIzXTLlAaNnYE0DRLCt5a1vtc8VZp4cMj6x9Ti5fTFElNZLtu0pIWKgoW3DO4gSzfKVu3eim5L9
OmXqDdBAx6ZlFWIuFtVd/EYgUSoZWvaLNrlBTypA+tvskiL5/Pxt9LG7Zb7mxot4um1zjhHkh/CA
p+N+eJXuAp+guFVvRNT+h3NzCbtYyD2BxMz9hnCrE8GHMtZTl6OufIJGIz17IJ3Yh8Ex+ZibOXMP
9KCOWSXZmaWBn1MF1C8ODlIAIKQZR6aYqcecIQAK6P77qMBQID08VAynrLfsw6o7VV5ZAyo7nJCo
aNrAW8xK5xL3e5cYo9uBn43xTIfwRZM/7NKSc2JmWV92iUan+klcv1boQm68yKArBb28qNC6RceW
PUp4CT6uih6S7MV5pgMq68KzdubCfZkrynYCc6T6k3OJx1Qtdfy/p6A9eYjQ6mM3Vju6AxWIJl8a
90dVNDAuzI5kogQ9y62ZzNGqdMSLEMYQx/VTvwQA0dKiROQf1TkfP/L3731S3p21WeqQMabxz3Fu
8Deu25KwUhRnYRDv3iB9gKvk8Tyw5ctXhdTjQKB9cP9gyWBv9fjy2gOom1lsoz3KbtPIs1rOSYaK
jpjNnyZ93MKcSp+/MrO/IdH8T4I2Prn6JnTJfF+eBK3QiCK2r87NoAlTMPIblBYV/XZtI/+MVskK
n6Jj4iaCmzHnj2CFQjr9sS2YhXizQTv+LLePpFNSLOL76Yopdkkl4nwTcm30Y4ZVdOQXDGRFWm/K
9JREIhDhZCnwFx2of0bWRtIxqs0IFfF1AeiYqQLpM3TThmX85n0bsQgs75dP4YvxfCmPxUVPzAfF
XVzsYk5O9RWKKgO4YicTgI8EZICvCmQ9/WDQEdU+/aaQb8q37EgAGJfPMZ9qsIshTXHHVkyQkKaH
nVLUV6u5Enib7Nd5sDQUbBOd6fOyA/dL6BMBWIPq3rdmjsCmNhOuoIlpN6smaMM2q9s27XbYVoSn
KBdTaRblwWiHuwBsPARNIGcHxM9h/mFA6iBvjheLl0oe9E4wVC8km/fu2wlaSNqgKulqCCHEdNc2
whSRK7emA6339qjucW4b7Sapj74j+xASnTl/bodqK9l8dFZuINRd6lST1rcD3q9/NOMjP/wLRT1i
W1sew/Fs+pk7stNUANf4nVMbHtvV28VU+mlgCJvZunPkZV741lcr1QBcmItA2e5Sh0E+qEgGTHg1
YkrPXFyxGd2v6UmU8S47MlRIZN46k7pppFo1LS8lshtfXg0jI13MdFyztMHDK/sddkNPnIBpsY+Y
XsIjwMbJOz7sTCt8nJHbliGrVSH4IRWPebSPzUQS1A+PniiBA8w8ZoKd/Gbgbt1kwTC45ehxO9gT
OZHmHEYUgIpdinV1jrDZhoUoaM7ujNNxo95u1xoyv/H0lGMTe0NwJCW3x/gZtryWbkUBK4zObqus
jZnIZRISRU+qUyQc00yw6dUP/AM0CqUDj/sBPT5mXa4fQ5rmOatWvxsp7a+AEHFugRq1Y+JsL47g
ojG2JcUyCEE3tlejjgOWhjf4elPqtrTmo78DTfPEEmkPaIHbIfStcw4Sr8ZwWhTJBoCbfbvMc2XX
ODkms3Vqt5oDeQ0AaxacbdjEW5jDiiHdfhpJpXt4oFgeA1S1ZZAxHo0wwk9Vta9/B5fGPU9lng5j
eNdPd+ie8ehq1GL69jCqGO6t9Gdk7Pd5+HOXYJVXdHMd+Xarx+jEbduW3DyB7jUhTKgx+Di1i1FI
RVeVbMegLJ+0YdL5xU9AVlfhMaakvOPB532+i83vu4NggZM0mJKmRWrRnoNS4VErrEXR56tNMbSl
iq4RAMIj70axjuLY0AHG6/jdp3dG4QfV8UKzB2Qv58+KzNU7XkA6mNq0WOas+d4lfzm+ZQhHbIr7
a5MFMJCPVRKVQEsFFw/JKewMFxoNWxPX1v78l3JJKW50UWvWHTyhgrJ997x0UOS+xN3KTQGEuIov
FU1Re3oDk6O2Vm0ZrQZBSI6yq5U/GILuehndLcs5iCnGxeBEIaAusgZozm6dsOYu198zGp822hku
CmfTdseS38sxQNu3TAmocuHvw0oXnOA24OgMANbPt63bWGkWlfVqdO8IpYSSOZ3S3I5QevRPyfAf
sC4Qbzcc0kBTyuEiGQOIIeoy1Sw1iZhTdOTZWa9BqwdYOI24Qd5aAt2Wq+hfo8Sh3mu+Tm2b197O
Q7Ywul7tCVXdze1YkFevwGLaDwBBnVTGUtfy7N8Ki8ZJlMVL/IFqqACJzGVSjemLbOrImywGhj19
56lCmLQza3iz5DKrbJewWxdLczKWnu80bgDFrNsQu5JRlijPyyCeVWBXy6NShiR/UqYxq21hjm8J
sljDLwR3PDHlfIGqhCS3CQreY2stxBAxwEsa1Ukjkh0fSprWKVHL0ZBCEegrb3TPRP+mu6c8nrLj
CWAsY2KXNhUVIyKW3QJt2W4rAfZGzzNDtQquV/9getogAdTmYFE9O26FF/1ywZ4WEp9zPOUQrfr3
UHWtJyDFqtIZC/bP9z6xpdlUkwqswhTLkyyZdyNhKJlgWB3oKudOket1KSNa+xgFdLsTkrT28KnI
DGL/qcPr49tKTZ1tTKbvuORfrWc5LZFLrA/5Zcj+R34UD9HFKdEkwKdCwr5SkarebRi92g8Iw9at
pqvApTK6hQn4As9aYVV79nc/njOpUAPkVcKPnttUV0M6o2y/eHYFC9aYWTVP/sxEVIgpwCyncceP
z9XPJYLSfHfIs5wxLfSGCekDni2GDMPSfPe6963o4whMAu6Jdk45tfsjbx7xCCCGaFcaewTsgM3v
do+FRVI8xRSZ/5yIWllOyKbRM+jkVcH6mH2a4RiFH0GK9zkTY7Ut/5OXCBu8RHWwMrwnu5xvwhQD
tU0M9qK+UnmA6gIugus+A0mDsL1BjOn6Bj3bY70ls5S6t4Q1gDBQlBABgVsVhmtkGPpwSDL4NZ0H
D7VNs9ue6f737vaiNRSbzrWGvW9l9VCaEFgbfTAbZirW4Qt7a6GHKim1ho/+mIpRwrxUgaiQN89r
OzXqjHv7/qZ2Y4+6ZwJybqsiNZCjuBJ52mxLO20ZSukV4ZOh0EP+3lnzpiJ2aPwSJQQ2F645YDRV
kxK9C9aDgtqRh8mr9GDzrWC18alZ8UGUKHq8SLNvwpVIm2jktOk6XkiBvq0s+IClLRjZAIfODVZC
u237wZDxLElsUTp1f3r6bk3dxGVnmunpbQVyF9JmEHUA0rI+a66jgg5YQDY3HQA1/Ox1HWVV4qq3
aIwBDkCKTvcBdVexvX7hbL9G32wAi57wW4epc3ENzSzNnofqRAyYDS5vFd9BhUz9/K/382MdxcHA
eqyqMvvPeHcvixztvIh+fbbKNp6nXrPkmwwO/5frGDqm5T8lDDWjGRXP3uEbZhIWHRSjXdAHAj7U
xhYCmN3Hk+wVAx5IzCtFk+ZbRRRHuoEhAgHyPCU/dYYQLDapniIS16l9Ib9h7/RPvMfxjX/N99T9
NVOcNft4+g7+k6EkgpmeT+MGleVk7huS+6D2drHWnTAHSXPpbbWzkDszeFLh0ePOF0VUakKHNYlu
JCY/1tUpHe5BPn8O4wnEMdPvXSDISgYVErMtB9HXeL6qYeD2hB3q4YvM0DY73vByqJuU93zqXEOL
6nXxx1YLjqUcSbB2pg02qgAJNX5QpY7OwNO/E6NK8dgf73MgY8aEGX67qN/lvLz3gmnYLxtNYRm3
QRn1esdjrpKl5y6gaicDK9iSv2GmDxbItvH+HEllaOID3IlGCnHZ2JjzZ7qpFHQgxRZySqnRYb8G
JePgFO3H1ch/kVGoy0j5gkKsiWUIprr12JHey1hZG2hJ9Xtk9u15bXqeuXNPHTRCZgDk2KbHmbVv
933istnvqd6jfGLDm6dKdVzsPUY/5A38Yz8GqNSKLy4d7yNXRIAGRjaE19u0UT//ctY6em5hpxEY
3GMFsnBtCalRoZmf1H7zuUKX+g3oMNOTntkcWQOICfHVFMeG46XYXP671W5E81Q5kY5LM7hIe0Co
HxfUtikSmAk45ZOo9jn3iWTOog3+iLYLFfW+JQva731FRDZLqC73YlOJ3lebB65MHE8h1RpVLFX7
G2+vZkPcrQB6cWDtxGubRaHSkrEmum1e/dwqNslwxGP4yY0FJwUl5lfGQ25B22ptThZ7FzGrVcvg
YwTzwxrDRZB3uhYq+fRkJFVN1vuIU597eeubUt5fTBAXlkVz9dQSQEA9O+PxmzWJ9GXfrmHI2EmL
DrexrIRA8iWWJwGOo2gbZlblyZ7Lnij9aMYVYURl+ZIGbt1SThIVh38n2eo0tvEfAh+NM8LCynVA
GCgfFRWygjQfDDM3RA24mRlpGMW1kaociqabDZeppz7SN5SIufD3jR4LXfHxsJ619miItDRaamc2
XRtBwaopwPFbbX3C1j9c/aHB2bitzVoeB7SUI/V7HV8JQIvGlYcRL84VEFXS3mAqzYSj5KuuGJoq
xnAl0yaN6mUteioOjyYbprt9RyF10xxxYwfpFSbxIDKQ+ejCl6S0zn6mbw0mOyN81VK4+lSpevT5
bSWWtv0wVJ2sMaB/CwZpWdiN7tBtIfPiUr8xn/6AgURv4C6h4QODNOjy6d5F/Tz1//5hAmuFWEt1
27eo3wrv1ewFphhBf4pbGj9vzF6+aWRt1btP6SQ/C5qVWrKbeQTyp6Z14QC/X1mZqfiF28hCSiBa
PM2TDCr5qnMGo742sMWEztjahDGxyMpiJltpv8LdowIl/oBh23UopCv2oPshIP01uE0TqmCsPS3X
xaAWu7G/h9i92vUY5OrYswE2dyS+oWHM2J0wjle/n7ZpUdE3kEuy5laGwaYlEnKrwl9KgiCeyvWf
GbYtnIUITRQJhI+j+3MaTyHhqkIzjB1ZbV6A2Oc7Ou6UTy7XlbUx3KSAiKtDTg3ggE2qCH+UO1Dw
x9JiY9jF0L95KDeJpNj5eWnVPxZOwUniQCSFcNZ7kbqVcRebkXK+Shjmbb1NhM9eg62GakIVhtK6
l6clgmR6KL6ieJUcp3bz3Z4447w60MlBhudD6s6mwze5N5ERR8GavIdiGjRguiqJnjMZU2XAzrSh
Fx9/6I6bUrLT6J875mGQ6NYavxc1lHMl1Ra8SLzdoiNq7uQI2RhotEzVdaH5fgWNgGttPEonDnW6
L7Ea0H9f/TJlBdt2lBQMXEoN5ktojqFHKbn35xhpLGu2Ub1Ieh9uSKEaDCoyiQ152eUjJg2Z8Ir5
1t6soesba2lXZbx0nfhEVO40cvafdZD1OzAzqVSQ4OEejGSL12//tZYLdY4+WbjT9nZt5o4HfZ6I
N1map33SIzxZH+rum6rCsfY6l8INDlkK4GMeiNB535Z3k0maNDfbzZFn+KoHuUXV44sp9w8U0NWS
sh6y9wl3S4DGCoPW9Kfa62QbHKEPrRfX50tH4IeYxrABMwwHrPe2fEvlZB2Ycz8FI+IlUJelhG4D
cCaoeuOlUrLZy0escO+58hAm48cyJw6n1BQLPUwTsjh+Hd4CMDOrnT41dRwaE07owIQ3glA2s1Xl
Lu5z5E3EUwuYldwKPK1BUPGNqWLi1qJSHoCqTWRLHAZTpkh5lREBIroXI7QFnu46QCIqksbh8i3/
MoMKHGampwLKr6GM801W66YWGekK1f9IfAlw4FwNE2L+kMWz/TOzhMVwMP+chugswc3uTAt0RG+G
2l/9HbqVkxzE6iic7i7hTmdd1259bzEjbfw+76HkW3xdAilyI6Fh5NfsITkdCjPMnvIeecIl5Io0
+H9nsQ+NcRwfVCj4E6g5H+9/Kho96F0/5NzbpIfSxuW45aRFXyFs4XeJFB9JxtavEl4hG17m9UlY
KNSlTHQYIgx+lm8gVQUeCOyjGikWjgpLbKJ03WLMOEHBTslOHdkJSN03/jeT0bjWTbC98pIlwWCq
UEB2yD3JJhi1y+JkEoYsKKc020/hHvLPBJo+sjC3P1JCG1wDb9mHhMcKim3aLtrFPIwa9ivCNbr0
Ji5CNTeKXgu1wyXvkFJAscNVAZ8PL+CxSd5BgyLDFWk0hOd3C8sjL0yYJlsuIoPEd2dUoT82XwFo
RK3CXuI3rVENcmSd2rBWQIa1lDgITjGu/FnVl/ejrbGKZZKljAWhsZBS1ASTPQgKrSaEaBiLXJZN
p1QhuM1UggQWDwTlXyfpYfyu7KwN8j2TUDZ1qszUIC7bvILZluSgby58QjoXZOWxm2z5nH7Igf4g
x/+z6LKZAhBIDcXpRfU8LmzutsvJiJbJXAYC0i6Rtx+RFzOf6tVtdBeChoONOXoNfYPgixD0ycEP
n1qxf/s1IqyOc3uWkK8cTBKGjLUXHVw2yuSqPpDjKA7tRXeND0WO2eJBiVoxYVzjsq2CVBK7jOfc
XkV6HRimotOVENttvj8Cqr3WsRycNKmeKspoilxNJSILPcXT0Y1A9o0iQM0LXyf9kZMd4GZV/gl+
4PF5LESmebvJROm3OZqWI9uVdeSByibJ0QhD43wDH66Pju7/oykPAXl3s2XIay1Pey1UjmXguaL9
9NkEB97ZVNLG9mLRe0jNPSGV3c2M5X8b+/sLZ5UDuKl0YPgcRppWEDCE7cLNN99w3e0wDkNqhMoO
WcAIvF4cP5MM9PCwky3hFxBK02Fr0vXiUwthlQRdPzIfRb4vOptbwYL6lT5l9fxEIVRdxx2ulc2C
So8QEapS3t5lVci/CWadq4Fm1K2SNP/ZHShbIZid7uoDsJFEGCHDsA6SkW+lhJQxvAe15SHOwPBX
P8MresNxdsVNx1e/ZGn9xVoPHX+sM6wRVW0QnwkWtxqi7g/HU1vH8pA3liwoVGAVVcej87NgbREW
XOQROVXXDHojCPkSHaoLe+amCh81yC80ChchDuF0Q2baJbulkOn2VrdTbjfBT/If0yTssZGUpOwF
vwgVBs83P6GfuXjWrlntUPbK6C2UB9n0MG+8msjpFrTTosJpmYOMZex8sK/V+9mbWSXRx9M9VQuc
rICy9BAITIGHEhs7jTsAGwRl3jzVxWKYYf3ymiGBez8UmH9mLuHhiBl6mKWCXUMuuAn4JDYhOphR
engFBuCme0eLQSpPS4FVC2GFm3SH3i9LkHpPW6NVNT/ffjDhTHmUkkwCUxG9UpdWWZufx4LBAYDg
OkK/h8ltNqAtAsRVLdGC+SKgaLKnr0s9WsTKKkBAjk6hA2YOxuzkZdNyykSkBaDKTaANBvKNjXa3
9p359TSYwzRP2rAeZbDVqOW61+4oFb7kAqKw8i5r/Qn0Uu3J3PKPs7p0ldCao0pNbuv8rzyeCvFe
rj7hLJCCoeHZZLKfReNd0sb8x/ZdkFAjfYRTy31ejLtkOsok3QRg6zh+YD5FAByc36mVs08h9dDo
64oFx2/AYkO4LsQvVHmw1XM6Gq9mqHBZlFlt+v5YRYfzuccOYquEEKP/saw+oIlQ/5OK7+xTBgk1
fITNKePHg3bBt1043hxUMD2yp+oJS9wakNfmRLYaItzOdNXcQj7V+Q2ncKX3wdDp23PQnlEyqiQQ
zSOuAaWx5be86FxYwTY36MR9VuV7HY6hQOwBKPJw8QpRho+wwLXmU1deRNAFYjNkw4GDy+27KIqW
FWQiQ19Y2DMGxlH7MiLknhcsjUYF2AHYej3SdMfghwEebkv89DbF7w9xL9k6zuLelMxOvGJL0RmC
y2PuvEDI+xPpSPdDI7hkV4Ur3xMPik1r87JJRIRH6s2GaWA369lLRFArCLNHbn8K5QTSzZ7ScqsQ
x5uhza7gMJZ3zWCpuwGaXyTUF6IZ9yEg/nqMWeNpj5gOQwoimXIk9iL8V1SNamxOQOc4TrVME8i8
cE9XsDGqMiFrh1MmPehwrmfSt5c+bc7sV5IUAucrFWQqKro5YSN+aWw8TTYZAy8He76SphKlLwcd
D0wP9E6aswy8AACQuwma6vOgLCREMgKWG9zoOLdwxm3KDXvnH7BciypNr0m1f4s8FdJpL+hUMrMe
h+gcS0FaMo3S+GQB/w0eWqnc5+8x6+igz+lAiYkXgXRkgP6GQ7r3bOipC6kbqxLmdmV+LeKjHbUw
3IkvwpKE0EYKDtt08naHYGFpGeT+SNqaxewG3dgk+ZTWYHMpZMDV3cJa5niemnI5Kx+SMCzZbSgX
AnZ5z7LqWyB2/sOKvo8+8QqwiFNBJd7reBbUuqLSdGRfWIJB4GFYyWQQ6qNt4jircxl7KavXATSR
qyoPj6aVfqBlM10Q6drO+BBNaqUURzCLb2uy1rskPZ67+bBDKnohYLCiw1DOROgoxZd92kImrN70
KnNMtunqILMo9YQiMTa6pnLQBYpHYIESj9OCNlxMacpoAYHgUx60HbKQe2Wkx3rnOtkHVAgBsf/i
/CULKLPH32UrnK6ZZIeu70Udc5Z1CLQGxAKLprIlJj/w/pnZdzJM69ixfb1BLGXdMBB4WLuCIK0f
FMDuz7JDcMpIdKomk/cbU3Iv6/JxqiMjaExSzEhe77DKbqrlXuBT4aiGaHJsopSkmhGeDUWU9ejn
6PTl2ji2S96OiMc2iuCyvGk07j2ombKVapsCM0SxK9MLeb/OnLPGZDo7X2ifpPaNR+2/NFXA2m+B
fGu09pyGAK06mE/d9QUv+EYpCL079VfAc15c8tiZMWRLgFI6UIRG/sN6yA0D0e3f7SN5RwbA0/E+
YaSd7iFLRofkwhtGcwj6+mWKh+GNqwvcNXuEShDs5MIhoNPE9bhaJbGA3j7cONmVB7myK+8OdZRO
JU+SXXR+ohQmB6K7zv8Nz4JYdtgBTiDfuAMEtC8W9IFWWJSHiuljYsP6FyPHr8EnJWJ7GFbRm4Tz
4xLExP0lz5/7jXobp9M9gKbRNYMJUwGF90H9ktGy5bhhl2h6KjS3wD+X5a96w65ONXIX0REjEi88
NxoPB1xrD71TWNP025McexGd8mZzwN6i+6D4MRYRIorEqiGgS7RZWPaX8nmOEbekhD4YdSbRXDW/
M6tOgmjLvnCFzZ9GsUdPYuDpM4I3qEudjDO3zPtjhjAZEq5mIo7WVuTNgqXLCCI6gsZl21JVN5Om
YVKTIV7YLrmu56kvTwP5RpRhZLs4X/1n5aVohqO41tX1Yglm5WxNnq1Mr0joemaYUHi57iAqud12
GdOEawp5jnG1HFV1h5ZfretnFOKTqTl+i77WA8h84Y1/fFJX2O5KsWPX0i0WKiAnoflTAd/h7bUG
AMCH9y5ftgmrZAsEBWGjJU+AWgVfplvPBX/fn7lMiGl9J7kx/xNHtyFY3Wfpato9D4WvQfcU5bhP
pGbztDT1mO8n3HDwNnluRihWCXgr3rKzyieAj6cV0NOmooWDXMYR4d2D5YMDmjHKHRiRHDm40ra0
rtaZaX774s4lokDBUzIwCvby4cnA4DbsUxrZRtoSNTTqRjj5DgoQMv3tEw9zSP96U80xexD4Izqn
u7zLm9wVNIHnX117MBS2VaAl7qiih8Kxs5nEIzg6UHAhdrZkVp0SIBrEen2yyLg37QG7qUYy9skc
qe903osXB6tczq86bVm5ht95u/WoREpatUfaG55tmx++A0w4rNrEwvXWSsXiJRkOUQXL5ZafmtlG
NZ8zWXK1zbDs3nGkOg1lDZy2ytEnMyyXZhtZBSFseyefB8huJfvAeKSV3lpIL9N7RpsnhmIt942p
fefvzCvBB43du3R0+L0tgMhcutfmVsmTtnCQZjXVcwKWE6zTRYKIVLyW5Z3w1qzBPfWcMY7fdrB0
21PutajiQOSqOB8mul7Vt07EkqtA+3B2ahTpghDo9Bgqi8d8GA2SuXtxkjHlsxydH6RE5MDjhgdp
vyN8Yph8HJAxJwubqunFKVPQmcCa/KSNn8/wkkvsg8LMwJmoUqKmdDHYipprWcb8+PNaeG9v1Nay
rRXNGlztUuRaEBghxRjJTbuwus24ZPrl3U61VjqiVPPLns9EAN4jchYRx35QkdLwELUjmfCcvKdw
476+tTkjPoRsfy9tKSYDAV9rwkV6SNaLk9ACiCXIxW9fGVTvUdYkpneADyv7EP+sVmCb3l0Gzxv4
jG8MPua3oXK4EQ9KsMLCScg4bw4Vt9w5e66kfN865IMcEErxFO6YV0RPgrZyqvSVdpYI0Vw0GRQy
7kAGSzSesC7HdBcNDyXGVEDGnHel6TwqSL+49+aSroYnyITz85ch9tH+VnV8wcUPL4fGxg96Tl2R
k5qeJUZw8YbAWHhix6sQ0dphZQerutrpNxmtv+HA9pWwj2Xz6mkm/JLhTtWCJGvP116wohtLhoTo
VrejFLZAL9dRUEAVVDyII9tEoIZnpq2Oo7itrlwwn95z6xbtsVZbrtLChJJuB378V8Oq+9fjUGzm
Gy/zfwKJArwPuWSAL99E0WZ9Cnoo4q17YzudMvY2qgpVfN81BcWK2XVTgbFxmcmXguu5ReGGJ7QQ
KudJfuuuBW/ujQ/YprzfTAxdo5sFc+ztyGTPDnRY4+C/aRfmGpYIdXj6LyXgnD4xw7F3RLeSKWO1
t7opRRvlA4naJ0642dBlhb21jwyIIhMR5x3Mi8k7meh/enirLndMC8F3T9UG2wDKpew19rrRLwJ5
PPiU4CXnh3zp6HufVmmq9KRhJO5f5Iewfp+HX6gHB/L5YMJbCIbor1qweImD2O8n/XQpGUfQq4ii
xXni4SBjSJs45Qzbjpv896zQrnBTKn8HRPSDh6m8YtaWYPIlzGr1+KwmXUGy3zqnNGfXrtsQj12e
XNAYfJ/TVlfULrUJRXc0IBBUpPwcOwXZxZ7QjLVJ/8HFXf5OsaTCz9RKDkyOZkmLlzEaWOxzvKKi
ljte2Jxu8K0zap2r6yFfrntYOvLwwt5CNrTIYcjPxq6jZRHCfZtqLOv2OUDM4wdBIxVy45mUGHaD
DGvdI539/LIqB9vpYsZHyYkUTJymxe5w4XXnLU/zRmEpjuqdxttknM2rdu0mbgZalkNQySkPHLLi
YZbqvUUb5QBeXf9nx66yW10LPOeuefWeM9MG4LefwEKsTThLRPGV98qK7U9+esUUANQ4OJ6Et3BT
jctDlrImHHG77wIFat9sjD7OlXQkdJXQFJyJfwD9avIXBg2Q9w44AgLstIGd7hwc0B+eZs8IU0S0
UJJo9ZIIACskXv2xeasPm29ejWrWJmGJGkfUC2Tgi3Ndq/7Drem5EK2eJgEmlHk1bDkigHhOERGm
YhtoDIjEh/OZ+5WdkE3Dn8awKG4CT8K3IbO8sKalKKwMZCzUbbd+W/mJy05vVmBh6B619O8zcSMT
IgqrDJPrVKVIk24PDUpoAUK+8Cu2KzQFR3wDJ+wszCOrz5fYqLkgxvS5dBg7aFw3DZ2ijXoZcp3W
T5g1/gr8KGiLMG7wKTQimSOLO8pOTu9VbwZ90oXj56TOQ89QzSfSNCqvgFmEa/Zqn0cLKNTjJ8gx
sb7nK5tuEW34jtghCZ/V3JvTGUcK21mGEXEOscz3Ng3xTl1fUkcKXkjWyalgyGZIz1NlLqAv5Ve3
cnpxvEW+plZhSNi4faAoFkmIjfnCp2ZuwAQri5eqAFajK4sBwh/rYXrAF823gLo62wOT54P6GMjS
wplkKp7i2MTYBylrAaIZqdI9SJqp55DLncJ1rCCaYmso7phBSqK9eurMd8VFdPKjehkVqEbTOF+W
x6BofW1s9RkomR2foEyeuzaA/DQ4p15XMOE+aPqxKa8NF247/OMMKeV0eb1gktZiwX3YuADY+Go1
b+DypEavPsscgL2Gu3INdPNcMxDRkktZioUbd6XkNcz3lunCln4FTktEllqWE0B8VyNLLPxiA1HM
GQ1iD3a7JzeY3p+m2yXD03eQgOGvKbHZhhNv9DoaGjo134KtlRHYxyrd2hWK6FF8tcTBDEA9lXo0
9cUE4Hf2u8AbkVtiyCOGGZaJYkXfG1zt0v1K/ZexaImZgFUrBqfsjkZKS6EQPhAAuwaaY2TocO1m
2SYSBODIUqJcBYW9zCUvrMpR36kxQsFMZNyb39GClo6HIluvXz8fDuvjLlSc/80fa4XxML5WUG13
dHrId4m3ude5pOQm8ub+NzodPrL3pUjwVVhlY7P5HyW2DzcNlZ2WMDdd+VmVBP+bwn9r+s38R2Q8
SdXP0FhcDEw/z/5ZyAwaaKv8Y2IKaOIKNWI0bMAO19qvH7LVgqZ8GHcTPTOitmqCPB3eb+Iyl2px
eE0Ifn1O+z3X+b2Ojq4UDgaff6itvoUgLZOAAzmd/4PtBfPRVkFG+gvr5eQrZO330wY1RC3oZ2wS
oPPwNvJqHbdis9e3XVFcCss5t+wXuRqhe0XpoyrBoj6cKcXEEMncpbsGwClukaazXfpz1eVV0UA1
Mw1t0SHjDjVXEI+VlF7hm7HCPGNdvmMo6X6s7UMi1DmNKcqHVrZJRqkhVIfG8fd0UnYYmsvH/VG3
LmHv6XUtzTqT5ILHqAx2evjnCAVpH79mq+6OoNc00kJaBj9+oYkQZ7/KuzLq43XC7u8sylS8JaAN
fBye2B2gZAmBWasE9E6+3Zdp+e1ag/EF77tfxW4L+pGqRhh6otBOM0cPuJEFuLa4OZg7Y0AuoqcH
/GIq+7bMitcqphzKAT3X+fZ9diPYsXMnqFncF+jkVoeCUhR/2dxMJI2HHUSPGRuiPOUNP3DpII72
UzkAmq2eiCHfjipBqiujK0eYyZw80qXY3isq+vJy/5vz0ORntJEFtaQq1D+8dHa5YKpsn7F3zL3O
suqOw5RKn0gA/g440U+Ovwkbywq/QYdgph0y3HWhIr0LtClNHbteSBRlajdvFN3G22hAl/MT4md6
8XVGjSOMfRA0gCgkdLSEQnzLzte+PB5bTMQFNMux+/EWguLTJnCYtPI9lhg+HT0HeHKwkXFviXUE
LsA0rzzXSgAnDlRI0UTrdUr+2Fdshc4JHA65SP5q3Iu15FERvDWvOWEYhdaMgB2BLrTp+8hGaR59
Zx+0XhcGHSEQ2MqFCXqUuJQVb9TY5B2sPZn4Nx/kk3r/lE0ZJj4eUvp350xos5VMEbdokIlb0uyX
6zcrSrU595r7vhsmT92AoxH1EkIbCPMmHnBwKOiaV7sc7r+uXFNVO/Ba6pIOZAerRpkJiL5B9/Zd
mSqjOinOTtlh4A/jR9QHNxLRhVZhWsQcS5ORN+ce2UoYOFmjDhgSyZrhkeW2xFwCKUD6Essf+OvL
gS5Vy4gwaOEO0TlXF1PAAWKwgUNIYKqbvr9gfpoalGYKk2UdAhQoDhmxTcGJvrN74/J7LlvhmrLr
f1t4sHhCY3d7LeUFLYriD7Ys/qOjzmqitzfZEX2KY8BsdxhkJ6SQDBkFmClbGdyATvLgzR4p2hHY
/q7wriiIwJeH8OEsbBelDL+t2kA2AMatfoisN+cmQcmkF127kLezp/55b7jrVLFE2D4456VGwKqt
F2bRrjaoHo+va9eikHUFethPc/vkJVuDXOvJPEyFd/RnL2vY8VbD6vk7esHuod9GcG/jEgpSaWQ7
6xZzqAvampuZZW0OgHXSKFAC/AuCm4DxODANPfxTjSHW1gZFpznTyjthF+SwhLEBFmirDkeSae3t
NC0t4h/h65S/3DlVsCvYxxsiCr9Ljpl3XhC+2xFY4ikLUqt5O4TVgI0PzkWzVnQu12Edl51FiRCW
2nibHCasmEPS8fo2Gh68xrXkHeUtwQlCXwpNaTzWAKLdOKCTMywnRVz6umMZj7DPjjPFHclykaZm
rDq4BgzdCPdL6jcGfj5LnBE3sH50el3qWEHIUad/89Kp4ieVh4Q2mh5/cN/MIy13IgMALH5823HP
UtsG9SCpyijZMzVyeDQABBFYnU51lkD6BebxAYUQK199HDzQw09Mj1HaOG2waQxHqO1fabxjk4V3
BbP0WqkzY+YlQDR4/iYkWTS+6mifkRbH8iS+tFUg9lhSlqI60ATBciVblT+Lb4HfBopTg+WthW+u
OW/NdRuqRY+1kydRGFzorwOah96cyY8/UL7ud8izbYFFE8/ue8NM6MgJLh31f/Y6e2qIiN0YtfR1
oWSDtjsHAmQqonA9NfDV2aPOTFqTXpeoOTwzwiIbglyKKltYKsfbCZ/nTJkEqriYm2GiPts+8Ow2
PHutDvtyouBWFbF5cuScQeevxSykgzCsLovKs/LQYsI+EAArK9dAfsKXGLcHv78k56sJPtiNlRdI
IbLr/RWydqkBEV4cUl5d6YlhZHLCdCDgZG20lGC4VY3Ey+IZ0cIZsJZIkxoWxlwHnz9LQgCRcd6p
rC5RDms/vCHESDQh7H/e1U7tpeqkKGDWTJb5/1Y44I8IXuZXud85n0xF1NAC8EypEKpMdhb0YAtm
iAdtBYtw85Is6fDf79Y2UTciP7xK78D3xok/sV0Ofgn2tsT4DHDhYnRC/1DZySMFJWLo2PRECUz/
GHYzW55OZ+389cxVbhzAvwjkOEmM53KbN+iF27ApBEv54wFzDK3OnTzE91dt2b41zVYPGiP7QSCE
A5tJfJr/6Ktru5G+8LOtuAN7nFvEUu52oiOswlK9iSulS6PJuWPnJ/BhRXAQFm1U3ZzgVfDdmIQX
y4M5+2MwXPb815VkUboOa80rNScISasu0fdBNITLs2IHlf6R9atu8XTIKtia9JuHFJl/XpMxdX47
42oeiJCDRSzqXcRdYaAJh96661vv28+PYp5GPN0D9iGKWpqmEqkhgHxml7RAs3PsUd3LQuRAKfhG
iyTmMr9Tv4QhzuyydiZ1r6iCkR3r89suZ4E+VI0NDokIpf8I7UjjiHhYF23MmpztlKisD63ZIPLe
mqSr9iowKAleBvAsGfQD4tOuHI7u4zbwQnT+RTsl7CSXUD++Re8kh2wK983gAKfjlIKYj+blkqHR
diy5hTNKqBAQA7wEoENYVJpFLR2rX8/QRGnNYuEyeWsaDCqp0fbtD5QUDLbKWo8iQW5xciK0gDjz
31lFp0Km8lciihSvC88L57GGuaMmn+mkW1RE+XZ7jW0SHRbcEc8FRdi1qqB2OYTMjV7JlGdwYUte
rWd7pYt7CCUeQqLnpN9tJH6oOjxw5l0jmbqU3AYcIaUVBb+zbOcWdd4qHutUByITDDDr1nLMJ3T7
EUlYNcoQShYYfYFm+TqwyoyStcSaWu1o22k3BvVZs4nyVgT7KpBEX22DR9lFt0QudWBdRR5/OOL6
usuS1+vYMeYDnsvmbDBEKgjiRsbqkW3VyJ0qBm9mAyFhLTvuNNx4oCFO4yrYSGBSjVQcnKo1rnkE
Ms3+oI3gYOM4SzXyGyUpQK09hxeocZC3eKa/grjGQB4fBPf8+gEURtQRQUNmgQHMgUphV5EL2Pha
3UuXJTXYLLC+a/LcypieuVc/mcLSepeCaAyw94mqhba1A7SrqdOHP8g69LQmn95qIEH9YJNy91Cv
rzZV6SNayMtaa0RwyzdRvVqzIMqs85QTVHdsglwHf3m+ksGYVCZP4sBPvNpQgg9aoU54NoTbC84p
HhwtEJsht+OY7O+NrH/N5MYTo4m5Yqsyp+qiLGDVVib2Njdt0MWFe2fapzAPdok0r4kw9iv+dFXB
JHAhaz9sA8YzTSubyfAfvYcKlUslx5whBO4WXonCGyFCwhaW063DlVRTnG71+inKLLwN3q9ckcBA
L5rTUsDTT4BMjJazK4OnroLfMXJ0n0PJuj59QsdjGJWJxHR9Ap/gjRxGVwjQIYUdDTuYdKw3OTV5
Jws1cpXjAIFtBYbNu4pA+R2GOj2AGoQDGP4xidwgzXsHF0AxMtkmUeMuoHTP3T4+++jrukRwIQbQ
Ga/cbfGGH2n7D3J39pHVdwIJ++9xyQk/F6Tya4toXkdc4K1gNgCa+bimReqFbwYfXKiewSF5jMGd
M+DGh0vxhuy6DkOikmkWdUTpnBurkWw7VHavc4RnkE7NMfzIn7VBs3Zos5QjRvGeChfzlLaxa4bi
Om4xf4f3MNeIrYTnvJ3yKGxyDRSSd0cDiyp40pvfvjAQanPKn7KDghXwswig6Cl2n9nh5eSBcpeu
E6jFswKCydNsO2iJxEthKrilX5SdWo+TZ+KUJ+tyTXr1ZMRZjNS2ANnDO0aKBnGEZ5iOjGMoEOpy
fHTOoZvdkAsMo3VMwV0ZyGPpLKwVOGcpsU76KqmeMh2pBX1OI7AE2XD6OYJgy9Xd/WPtC4vDH34R
thpicWH2IVa7HImsFQXqosBcQES+S5GbjJCjiJvyAMdV6ekwiTrn68eF0JD1vIJlc+Wt0sVARi1t
jGae8aMY7lnSu1+iaCx0KWPfOoPantIr5Cc2N8ChcFZ7YPBIDXqBbKJ8ol/Ok6tcXE+/pJ2hCp5e
/4Be98Gq2ujEqzqX2CL1u3WBqITDd3eVGc/O5IWTF6S3lAwt0xETo4U2iMlCir4o/3Y8APhlS+nD
46j340y7KZI7/Iuuf1aMvHvzq9TnJYPqEQh/9eOr0HKo4Zgp7bT1fAgT4HNtShgXdMhcUJwtaBWB
q/hxu6XjszsSxT9y39x/tS3mEFxIimQ0776n7Vav2pV7OP+fIG4qr7b04COCs66DgvZEIjO6LENq
8cFtKPxeL8DRvhLcv/hmDmEn2yMQHMU/2yVG/RR2PULa5gry+7QlonmSXwb/jhBF4exlWPlMN+VJ
7a8hTTbtooGBeeLlf6KK52RricTH4FLMfpNjJxPozSAkt9l9JhoTYfXDpgTmLY8HwWWZzPxyrFit
ytHMMNpbtZ9R7qf/yNxJzV9x7BSRXKHeT0HYYiaBfYbbc1mMU85So9mdiCjLUhyWkZ0zWUUxW/4J
Ybo0D1lbyRJb+apfwDctYgFFgpbZ78bj7DGfHU3ntBGEm+jZDGA9jKBYR+5wDs0kkpHFbZ2bZQMr
Oyxx4HU8Sa3g/Qo0EGRSM16iy+sf5X3Yzo9b94RBuyINix5h/sB7CqiOZ1cWBk453PFFcwFQG47h
uFzwjKXUW/gQyPCvAh0zbn40vvHwivnayAoBPLWADeG3lwLLbKefkZvfzZGN/Yp5mf1MZxCOvQBl
/nQUcMLup20NI2f58frg4i6X/rni74acIUz6EPEXSC1ZiPFgFUlkKxa798hDmqs2gXHQjoLBQ8bL
1h5GCUzOqFQZALdKGQ0XFMVFyBIJBvbC8qywhTinwP/WlNmdYPErjtXLTUpywdtQbnmi/nIJGyhb
hOTul2ZoiAXbEZefyjUacto7sas2vcPbMzjEep9eoBKs2BUYPaebvpLAKcl8GF0/u57vdkYWYjv7
7kwAYA1UrltWI+Fm5QOPk9Rmjz5FIH5c0bbV0WubkYfbA4LG1prFi/3SLI5RRcXUer1EWlBqtvfM
54BbG4f3xwswCoiCbt7k2XDxohiRxcuWrigA3AQG1uMVZ3YuKWLbaGTi70vym/EqZf+ezseI70PF
16lThZpOXILu/Mza3b3y0WoA6MvXZX9EQnj/nlVJ5CKBjNYgJkZUZ1ElmcSyf9DAJPZdi0gTZAja
Iut35nEKM/jnlya2jDlUIc79Sz8tUQNOfoL1ktDxRY5vVDoQYzQ+Uqq4gq+zm4zwag2oVSmTbf1c
dr/tnuBNUd5aZF/fd1qZ8b4tHh8E/5B1JTxWBATJRwo1nOGtrD+Cz8SIQ5eiECYW63AIQ3JeuJxd
cRca9zp6vmZRL/zWkuuwyaWWX5nT6e2QXigoceXjnToFl4qTluvG8EFxjHquOoB36ZcBNORR32XT
pgI0tlM6X3urwOrQElWf/Astqf+TQHq1G40SDbXatn6YQsU+LxokWneoMX5pwWZlsetcmmSUtdor
8zJsFFNOhQFI+sHG7FKQ3isHZTtymqrjHFEzcV92bAcJrfIf9KYU7X13CQ3mOV/E5gUuzVXCECPF
Sxr9Pi34T4+vF3GqvVl2VTW6LtV+YfoUu4FBc+vtJ6P09h0YXzWuZMvFqQWGll+QO+SHDAd+hoJ8
chcwGzwWAOnhBiQso6mBEv4Vo7/1h0C8yrX28/CZeMSwKygN2WJCN4sYtzaKbSlc5o1c+3WisPGY
XtOQ65qKcy7q2CwsgY9y7jdLcRGl7frv/ACkwA9f4ULXYs6qJh6fH522SepFzsBcaZA5ydL8Z6GI
LDv9WY5lNfFvmKH0OkwjQMO0vSvqizjxSwAGwq2qnNmQvGxbSm4wzFTqOhyjxNF2oUQDDExC6sBq
87F2Fl/pNlQwbn+bZgjsZXmDoMwawn4DZo/Z9egRYYbj0hfvKjZfGcL6+qM93Q6p8SSTixg2NYUJ
WF2GKhG6Na9aR8qvaYZUNgwh29mtAyB082DqUjS9hrGojGvGmTXkJN+sFSzbsclYEdlxKkJO03JR
PhIHtSR85BkXpU7p5iOwvgw7+fQdY6irpdSjUJU83lrSFN+Hxc8kVmvTfR4z9ZoB43w+cpzKzGu9
+KDYUnBMfNVYRxHpdDilWpm09K1niC3T6fkT4i82sT83sfQR3KNMcXSm4k35duE0JuFEzr63paSD
FMpca6Av6OSKBgifcjR1jhE6/Cbnd3VSzmKv5pdV+t2AhFvGdt+eywUI48RtTlRYTpuX+AhFvuPN
cGMuZFQPn2dwUg1VGm5aQcF7hDoZwIrX8eTBsVjO74rrcF5p3woGhYu2k1eDMj9ukBSGDBioV+j7
uEqBsLhqhUs80Ogy6G4lhj6uEGvJdFRYmf2cN1NWSLoGdi6C+lmVvdsyPxiu7dXqVPEFl/iO3rcy
aPWwbDmltlGkC0g+hysfpVt1Nw5Khi8vo/nnl7pqxym+rWhCep1h7qDhm8IxNguG3to5f3w+ssWR
YvRFRDpW9oH7Ssyk1sqrorJIiDlVRSMmTjl03gp+NXFAjqzc9ZFikFRnVqH9qLFYTAWpxSzlLcfY
z5sO9+/X50GyJMh9tY6O9VPU8Vt9YP2mRoYgBTI8KJGC9zWLnaYHEKYdVPe/uX064IuSbdpyIQdR
rrGsvZKLOGpO69+11m/GTysEdR+jEKqZI/CnY16L16ZNNJ387WsBngXPVz5pjMbt1n9LsVM5sMgY
/uScZs0V1inz1D/wHH+dC79VqKylmi/Teub6wznx89FixWVgk9Iiha1RK+wzrEJvbi61z+0bpaqP
jLI3pHt5riUCdVsFGmz4009c78ODVsEq6qhQNETuAoNj7dpZFFTRa/7Odr+ZPaZV/W6kxfoEYGfK
0H2s2LZPjzty6VI0o1p4TOd9sOGgcLfeouFa9yutq5PgGBexGuMkBasGQOCl+Lkn/HhU3kLqzUPl
FFSxfyTbq7q2F+y6CcbP7wOOZW1o5EqBlKnj1RVV9WAAAqaXCoZ9THrS4B1DX4A5isfzGJDp+fBn
9FECJnaLjZMeaKJn5z2Y9IM7wO6baTSobDLT57r19T5xLB5VgAvkvx97I7WxD5nkvj1lWvSHkwLg
uDXx+pg2w8d/c2P6RUiLAewQV0LM3fTtkeMyO3Of6rngmO3mVlDHSBH5nH3cL25LD4lgiVVO9AMa
9i5KneMAx+fXlfK2PDsfBXFW73d8VuEP8yTDv+x7RfZyFYkfaTsjm4ThWii51ZNtsDz7C3HV2iC8
N0YJ+9vqjHnF1hBwH3M5fsKhvWJEPEwXQO2196axg/830uUS3WAf0FxvPLVH8nCry8kK8kUKwYW7
HtN3KO5oCwjoq2EYa5K0XfdooB9KhjlHUCtkaoR5kK0thgHEXcibMyLNu4YRBVgO2WovXqaGNBGs
aUr+M2XFVzgBD840+AmkQSquZcDCA6L1feo5E+OuR0iYTARsWrq6y8W1lOry6TJSOJ8n/GhBPvln
w85vqcTilFjsJuuxH5Jv5ZQX3JT3KmNZ9Y7rP/0bOjySlAWy9FFn3Se2EsaHisjyhn1U/rgqiLgI
JDlJSWjpEv6JzrG+yQJv8lTi4o/e0e8RkHXo8yQUQ8LFdhbHlAzMnNKeVdpu/WZ6/V9NrtGaRQwd
u13S8aRGRp/u1yb0TaK6jXgpvEpt5Usas9nI3VIJYdh4W2194eIuwEMRp5HrHX3klmQ1zPa7vsPC
u5hOpQJSY/tqP4TlZWIDWHCOvUl4j1n0/AtiPJvaykI0xu69yEb35isJ+LkIylnM5PPtXWcsjMJa
W4bB7lk7fKlb2+P9fQr58en7cwpE2zk9UJ1FXsCmwqgGWmAEbXH1nVEOjNwRxmSb0gfZsxaja/3v
rANlCnwMAMHkZOBf+5Z/62pL0tS65rrM49DTmnQuOhzYCZ5xWFUmmQL73huGVwe4RJrKBodWoOig
KVEVrlZV1kSzfhzjeJCe0kZZj2jkBxBoRPdxQoF2yNuR9Am/HBUIBS6PpWylagCMDrdJSmIcqTm3
8L8ZsNzJcQZLKaBWMGbbvITgCkjM86I/40Uwtou5zjMpvmr7F+/l9jK3A8dUuXhLZIm5ty+3q/6n
1/Cg2S+Mz6YJWJs1CSUaVnugUV9YC+bF+3YkBM6RTxSeiAAjvHVYAG/EX9otN3VXSqs7mu60ShZL
nJOoWOlcQoZaND+0eERCCVMQoxUXO9aNDUpfllpHrjThdbaTx5yirQTgugNwFoK93sCeBccMK9Zx
tNJ9qJ9sLxZNOHzq0w8yg9nP0c14t1HPQoSLmvJzNPLhwL0PVqq23oiFfMJuCr2jLxF33FbDcNFM
2Wc9LAMaBfRMbOI0m9nDhvw4pFAof6M2IPwLlHzuEQUIuaLiIN1zJ0+Z14FSMn6QeS7E+qI64o4l
qQ2v4x5PT93+vIHPm8cANZUGNtJ/Ir/5x6DCfJ4Goo8oJKDYsvLFkuthwNHyTgr4c/a0wN4zEUU5
+uabDwB45nOkQD2KIVJMshTeFjYkXouqxpRshiU0zVCQIhgfeWG1f8lFUY8uHANdLQj5SVqOOhZu
Jitx7vdhKyctJN8GM2/yeSuc70WoeilxJspdjSaF+NL/qi1EzyG9zC8aCFXVTfifsfBK1fwCjf3F
OtThIEmqZdlKXb+Lc5zs/IT13kWQ15eEPpTIjDNUI70XFsWxiCPQhjaw6z74rOpL9S8V/vbNQwC/
WV9ZkF3HSF23XGDT3dpA0Rxzb1e0XJD5F2OXqYEbxFunty8wIdjOD7JcbYk6D7EL14Keg/Q+LWvn
ErZW7woAMM/MmhIBrjPs5xhvR804wv2v8QG4L8NPlBssOXADDetiBwRIsgIRu1zucUhpsXTxrjaR
D/uWjdPzxUQpZGYP3iIyDgehtn7WeZJFZ/BZvk0R4iSsKAu0p1m65XvXQyH/VlgiQWzQbqRpDyAh
67XBPOX/tPMILsvgJE8t60/FPicMDbOESV5V3XYBTw0plIO4U0DIZfzGuJYZ/Xl8WvRCIEfBIBrX
94N0dEnsDeV4T1fdvfhPHER3kmVfGRXZPxeTBf9OtKOACLyz/8nd2SOBWH6smIoajW8TBxmVES6p
DNSq1mUNQLSe4x2OCHbVvYCUSi4FJa4aU/zWL6RKkt7P8NoJRUIif2KbGiMiHbpCmDqwCqnvrj3l
+ZkVdxm4Ooa5aDpXXC3L5fhzK/iO3hNRAfyUXrbMBNdzCY8gGj/BRS0CTcBFc5Op6C2DOhUGCJqS
emNWRZRR9qgh5ltQRMa+9YuxfedoZYOqe/DoyqGarfpFuIPTQ5OshfIw4JYm2tXQ5B/20XmUgYQL
JMJRc25+33SmVFqyfdCiUsIkwcV/sGqotqUqmEw9kJomwAOBYWuk88GMzLyo4/uz1RHBNVQxzpTq
8y7MeB0F8VCpYAQGPW47YhMZzFBTBdvO3hQpQH+F6N2WnY4cbb9rYOLBiYzVLw/6F3tyZBLDDr/P
Jk2G7dOGk44ulFA03h718uSX7znTuLq2G1gYNzAWZtR5WHfpJxvm0tpkqKl4+sDUM6UYNpp0ya+0
uwRow/wNicPBAQO/xS0h001UrBVq1QeZJrQ/yCrSJxqv5pRHIMcGPI3G2T8jhnShMJ5vTstpP8Cr
O3fkZaOF5FxyhIos23FIJ+U9Hv12kzmlg4Om2cT/BQW2yLcwa1NpsOT9TElqp79HbHtr2r5w5Dox
7jY5haOLX53yKWs3YDmEDxBz/TlMcME2EoBu7RWEi7mmcgCJ/eWeWqQO4p3g4cInsLPpanb4VUf2
EkNjJbSWvEUbTtXXfYEFLAa3zZtu6Hg6gJx2wynyDjeYqmmeOTUhWcKQc2SuIVaFJiLH6yRKQ3Vp
wwLAdyOUlrre+sTDpSBasS/F2dTFPIz8Pbs4buOg/EJvOK2VRGWWwNTjEo+wdFo1JC72dqiA0uPg
H/7pQM7+LAiPSerglheCrdeB9jVcxBF/hWbcR7R6AsvIkzROMgsZ0SbyNjtnmVaXRCn5Se7EEub2
EK+uJRsvNFSFTofoKNhIi1SyJt5vEFfOjy8gLgdGg/kFdInuiYgH063oCuHda0YAimRYM3SmyUS5
2ZBFHZjNorzyOUscOKt4D8gK1q1oT8ekI2/PbZawHUAG2xTjAG3k2UTyPFdhwIXsCsJ2J9bP+3eu
M8LNH/7pmb18RWsXVDoonGW1YZg/GBQ4VfdO+RXyU3nv22vYfIp18hp58j88KL/j4CBU1xipWed7
lQgTT/mIfk7VJsPZk9om4dYoO9a1fPCIjdn5HwOwclhpOXiSsZ7JGZaSkcbP4n77pAndE9YGyYYw
yFM7Yq7qvByClDsH+OmXHDJoqZ9rL1nC6XShcQoMQqtq/wHWjHvEEHc40s3KFeNsgjBOcX5+6xHA
HumOYJN0vXC/HFoYznpE4lflsaMbkn21i1zPthvLJXMkng8By91AIUTKwJMegrmCNck5XvWKElv1
xrSR8ojKIvx6R7HuyeiM9ip2raIwt4r7yLqYDINwu+irrVYxlxcYpyykrD+OJGPa2xAAWqHIYK2G
FEzeD3kwxGV9vNIizZFLt6YH9JzbNL4H21KE68L11XqaZ218YryP0nQKGE66W+mqXETB/OcmVPPF
e2Noq4FsXo1GoKhNfI1NzFXaSONGm74N3Dhc6e6BaaQLG89QDeuDExTe9aQlc/RY+nAd7SlPSN6g
teWa2avVRP3AB6KB/GHN+KTz2vrjapLf34+M/bNqVcooyMWMoVXv8UzlsKLJQP2mrXrCU5DVzhSO
AqlW7204MXC+BN5TTkf6myxdq8zdIeu0IUBkkX8YaIvikXPEd/TudmwF0S6Bv26/fT8wBgUT1tXe
jVogTWspYhZdwsbvxhRnE/amj7f8+WrdU+Kzqj4OWAFRpV25IhamYwchTOYSHXmKB7rauLP3+wZD
90Q6vPtEqt/InnaI/0wLV5j50rdciYkuM4ahgGgwNMDHXg/AS0WCueV73ufSPQiHcOyw6Bc7EzlS
rFT+oQmNzpuZAjYWhDRPTMI8N5+qoHb7Ecs88rxgPrsyazzfUqxyFKcvDUjR+6+Z7XLMDDsLFJXg
SGS9o77hYI+UP+gopBfvv+7EnkTCfOWYlcV46g8MyNDjfcEPVVWizEWjD7hXI6YkvYsOP1w99S1r
HfZvga9KxlTcVHpe6Bfp5+knm83hTuoJBNF74kIfUIpMy2d7g9pYZ6wQXPi3zR+HkuGIbiXTv5gn
5zmELunV1PMJlBC7opInCia9PK0gr/B+vIkbdmcKJge20zM6KwGzF/m8fyDnypmXsOCAnYs7b0UY
VpeyGsuPggKQMywleKWzUkqcrErAVOZQ9bI5PoAU69sxG27dCf9bf6+E72BEbu5Det1gi3/y1g75
wTEnEhQbrcW/+WloCLvI+9K9egPd7Q82aCZ77NW4DXy4enRBsSlZdKDQnW4MFd0zHobP0cj4i4Ji
kYtL4Ux4ODhFSaMS2IeWdNJSduxPGEVLHpen55J1ogj7MIyz/xBWx+oVMbm/03oLdtuoz8Y7thr1
4TqlKqgSoj+qGY30PeJsdqQmK7lnSVADmZEbGiCbRJT8fH8mZdm/mpSZ4EaCXGen5e6AVw3jhxjf
eFjxYiMSDztgfq4oewMooPcPIpS42TZP/yulzYE3aRLyLrlmUJOfjMsab0pM2pta9esVgBBFIJHt
ymJWXSf3XKQg36MU7pw1O6QkqPzZm/Zhwxq+wBBjR9twW194vBpRCtpyL5U02jQgmrjR1S+62T+K
0iSnLFgi0OIM0YW5cX8yqMKl+BOUdKjvEUJMbf7Z1lYN2x1faqEEcNFsq/MWXkN2jVvV0DoQXSj1
BRDdhf6sfDiK1r7eNIUWPZoHWuEEC3RtR2XuaPF5jEXVBai/bRn/d0IbLHARuelH7FZ6+D8MW/xN
3Lg50sFl0EOw99U2T/SMmXn4hbhMYEjVXd4a2DufOBZslT6xF7GPgY1SeKzG8O07iLAFXNYHSuPW
ElPO3Cv/dpu03e4ML3nLwt2NAO8xSpxbXeB7yEX7v51A6St+NnJvfCyYhp6F/qQEscYQj+DRnzL4
8K9lvzNaK+4liaB3qZpmSidbGsNoO4ogl3UCGrFCTmJXHUNTg1k8upxICieJNDqCDjM82CKq1uiD
hM/132ZVZFL92SK1K9baCeY+SOGI8Yh7vgo71bGdam7+dnbs0oo65xULFuvzHZyYwVxe48epqLFd
sMekC9+lrlGmoG7uUJGn91u6dgs32hkeG03pNcALnyn0qUs8bEp632MHgd+Vtuyb6CQCh7IM/7jh
vzV1ZPQJsVxl3BMTIU77NJiYjz+rBTuDUez93Ri7qD3LSaeTjOKc9Efmflw8mQcgjmZJeGjudtsO
AFiJXYweHvYQVVLNhCnn+jI4TTqNuLBhWWF3uevD2jE0CTdVjQC3vtrT6d6NFVwUkIv0UrPJjcE8
0rw383yoBwN9lxTfxFgqTN2iY6tJySImGrJjO6AUeMcXMfLrH0DevXNpK6WN/EwWNZ9/pO+nuxdA
s8Fl/bzTP4ciJrrcCoGBMfSkwccd8jS0MCfW3EE+wglNPqxv56/8aSmtGg/7seT6jLvjqlhbGsVX
waABfjKHg7kfbz3z7Ya3qh5AVxPVsEi5TZQBxp45t+SWDpMblTJjXIoDbV71q8j5ijaRKX30Wd4i
10s6KTLjXaCqHr3e9059I9QJak/HKG+h5RUt5RKUFeUrIH5x4diuJ1ZBYKZZuP00Zo2xXY+N5TiF
AYpp4nf1TXdscat2lutBGHtTr9FVNmPHzlCRG8ynUoq+mtOax7KAxJGdwDH0F661BMryzKNbogJb
gPAWUzwoXr1cjM2bGOsWqEjnpRvsK37aLqN3SxNepQflonOGjoRPycZqeJsPCRAh2zHOX/5ql4pU
5g9M+DB2o1peITK0grNE40aokUejr5lorsSSnHB0qCUWntCb4s5kkkr7GJql8cYVwnFupErGWSLP
9QxFMQbJiXBDD39REST5mfb9R0CTiIc6cAatADiI7HVD1k1KTrWcIhvieid3G0Nb1v0KuuRpZMRs
mIJmdVt+1nZIbA2yScUac03EuSlggQ763NlrLB3OWnCxdG2pxhM7kXQMgoxTPfheSKld5ji2mssw
j3GPXACKywwMoLLO40rjS87LA/6+cl88MIxKgOFUlJhcTExgcEKutOTm1MMGdVUTWTLG5mJkdca6
9x3ftM5ULassx3nhnJl2oAuR8Yz26dBwTh5FQmV8meUT5HodlywXj/KpmE4cdDoK9AlES3un+I7B
Iza29uFauup7o6S3PzlOSnR6TiUsyfBk3eZ0JB9ojVB/G5I2JhttttqaKa0/bZ/EJQLTqK+qS0ql
6k3TsuLlGTrhstT7ECxuxPCgTjAucW4vNSZbXl+RoFJI1V36VK3LS5ygoVZU5tRQ9nwR8KLcVV/e
PRNvabGyj4plpdDuvyXWj8gMCwNxfMliJpjs1YjSiIwfB37j+T0X8ZkZNlFlVT6+AbsKMoCkO56r
MxxVCuSM6P9B372H6CMNJldYrKbNRwvBn3WKs2EMyHd0mVv1MVjaByhSSCyAfXJGO1F+FbrAsWPG
GwAnlIowhYlnA5GoOfnhJHADdsMFIn54hrmVsng3V/2xjid/yXGU5z+BOCgAdBUVUitcmv62hZyk
E6UnzzHDSn9oDrnB6mihsacQP94dXDsv/xDe3JhOlB1AsKq1S3O2JWtGjSexOda0TLkRgDq8GNro
vv7GhmMSTgvY6r2tWGgtvlPmUa8TNRyv3Trob/SHJnDw30ltaoULQ3LdHmf5X5lQDn5Jo2Pngp1f
AHjPRWqANCsyhtyyvFmfyIO5OFTQCFGHd+UDMxgT9pOlVJQ/YfG5rUIzjm5VpTMh7BGHZfiXWKog
lRrK02R/djiVI8Wj97dgFzrPkaXXDGk5p31+K7JIkwUL2L5dvZMm5NM+KGwLehU2pgcQIyZxOgs+
2SXCtSknrIo5/Cd4KnSSjS5MHLeYJJ7U2p2O/05tl3l+1uQw/MVGb2dU0cUOSM4OiFZx1p25BO01
ylkOOmQ3rHhNYsPWFbX1u1/OvLOxnzVnBek+hEWuSFLVZw0RHH23czrk0V2GX/Yw4khS47VUM2zH
EfAn3Lk+iuJBsGS8+xKmHOXvdAlHUpjMRsps84q2jdTTatK02Ff06ONLT9pV3jlTsk+1xt921Un2
dwhFxizSmKokoY2hXqUuBNlbAePcHh8drm4gPfZPN4D4kvEoh0azL2SgHvD1K3vjn0zM9jozLneh
0CIPwCzyxdqiowHrqgh+6FMEfCGFxV2gYNZuPD4k+DIRnZ+eaatMWmHb9Hs/LJd0mjLwo1M4f0wq
0xcR74+0LPlX/GjmmGTY+V7YTDaDHIDN9efzSv2LdweLSlrCBi720lg2H2nhTvuJ9ZM/ag1jzUXl
3Cjvxho/eZJsm/SHyimO9kxfVA/TocTz0PQLBH5uzLCYPxih6jQ2eEZWjsLfcfbHMRMmE8G/jinV
+ShpTmcfpFHR5Jh03I3HobGfOivh7hgxfT5gkNTDHRTSwBo/WiShbba75mPvPCLQ2TFGsGtVaQEa
M3dU3C9fBfxGodh2Dt4QtMpk2LNgLBWAE4MoJQGrDaOhMInJ77SorrJQ0JX7tZAB8ryR5V7EA0Ib
qsG4dX4B8Bhj+tPnkZm7cIPLBRNhDwBzBRYYLpD54Zgp5Em+D4Ejxvrx679Mtp7JwKZXMhELKs3l
8Zd0eVz83UAe7I+D//VXtvg3X0J2oMxPDwKlFuR/ZTRPcudSiSvNJOOCtGszi4N/4qzKDFxV3+ZL
hjxq2CfOHC3EX9otEq/VzO0wolusk42G3wUFrtUy4YYFCusJsUFAdox/nsmwldlJocnNiC8pOGYQ
tLUNw0FHTEyx592Ulk8wMWe2M1MMuDGfPHf7VFCPEhHydgz2pGz9LDpLtgZNeWPEp4KnqO5x0DVq
rFRB+ejcgA7jCVPvjJeOQCt6306bJXIKtZQf+y4QaVLGttgzhDR5fbDFIlaNsMAPb4lfnACmu+49
kS+tfRSjWhcbqIBE2QZeDg1HfmLfShdJuiXcsll9WLUUyOPXMjbO9IXl6dtHRMmOFb/FK9Ba19Cm
uIv8t3i/qnONSd1q0tcOFBBOFy9XuPTIqrliEB8WAT7vaXKAIZAV/ihmN5pCgzmLTbsj6P8wivJM
eeSVQhusrnxmM+ZIY85f5XrYgNJtzh41mS6MoQAfSWSAOWx4XPnbw4HFwDBPjIU0v8OJ9M1zUvng
Zy5ZvFVqUGLfeepG+Q+QxF/dCO2EEUGAEqZrw5GdlzaAFJ1UXRJyfVtp3KDFvoJFnm9OqasA1z9r
1eXaKbQPoABpRSpKrC/jvOIAkkYyM57hKe6Zlu+3zY2uRyueHtMYrW56a37jv+t4aenJBeSUA/Fv
9Xv0MSyhgeTDAxUMBsRbKn4jeVI6rNYz17zg78N57AgbuMDH/JfU2j5YP6xMp1JPmElFZRIq2LWc
jsWS9nThEqTL6USgl9b3pY1TjCQlTqDP8Hv/3xkfbgKGIe1aGd4albqQhUJkJ+3oMoGKuyjfLzEc
5+Z9GETvi6tb56DQngDsWc9fulNCUjLtbvSFTSNgXLnEqNRUN475pBdYW52MH6t3j+x6UhLeUcs6
dkKV5KkjEQiqq55Dn73QrxnaSVUfEqfidiAWvmGOQ70GA9pmzuDWkUV9rp2wKuCBx00trnmKmHrn
CRGJHbIq2LiD0FkULLosUD7TpLcwSbZJY/ktIxmBPtJ2La/vhb8tiI6HvN/ib86uaBf69/yKw0vQ
0KMSQbK0ZTVKbUqyHZrJ7M/VXfEgcl0NkiEaybbl8kKJYj+xhW4yKOlND/0sPq9dxY3YQV59ZfBy
FM7hrd4pShaTtwZ7nk4pOSnb3rVpcK3f2+XvR3abaPJBMrdXQYCz5iwfZfPoOXUT4sg3yRpc2Ap7
RpLCAkuGQERZqsNgfiyUak4YiAVlHYTWvCyIj0Ejs8IC00mYdvTGqGCWQy377Zo/9KPPIxJDgkeW
X/pwD9DxOLSyth6xFW/2OIqxbxDGbjjiOzXRvsvjLR61EwfPwK4se87SGVSGXb4dEcPgWmYKpNd1
SRkZZtlCNnjQwSOa4aFXW+Jsm43BgQG3czhr7zEKs/wjQgqGTh7KW3k56bRfQVDBWNNqNEQ/rO0i
MFUQSuZRP8/qRQFsLTuOdInFfTuMyeWtmFx7+ezj7o41XNhaH//zfgJuxJT7+rdd6pc2RRaWecQd
P7/ZfAESrPRLadEayxpIX6POHw219HuRB+in7ZWslqwe8bBno8icyTVkxUHxU+E19DZIOkjB0ZMU
mDTdGmWgiCehMRsDvBUK6Ug8svDvK9qVqBj54HLiNSn5JunJBEprtqGFmck0xTLAcS389UQI+W/P
vPQ6zcsCAVIIwP7UZoujq1KXuamIavYO9wSUYVBXCPKCjTrvj+SwX+q9MvWCQWlt8vGuZ4sqz1RD
8qVaIz7MfHFlSha1Y1s0Nzc3adlCbN7EoUXAgBv3hrEvfEeC2QTUSdvXMg+2Bh5yDGODmQCKe3wd
FC8HeZgctSWULaiBTHEgGxD03cCR9byZy6whBrMm/rLLy3ggaMdneRXCCGac9R+PX2icJ85calBK
ByN3AO3vBdsOCeBuJ9sA3q1voTkAbUjfML0fIa/0TKFRtp6ifFvbBNURaPC0RQ8bXyV3JwwQsIts
R2d+EdgX8JGUvud6UtK2IrWR7NS36bi33P1qpwDokeYBdaQh/kWJ1EkGrjpVn3hezUWMQrPePFhN
WyB/Tbsr9imT/jtrpLmloYpThRxXmSG0Enmo9Ie6W3R/RU3hQI+K4CobK0FPREyy2AGuvCqO1nES
pdMNHb+ArH4m7mj8ble15VIx8Bomw+hKrl6MBMvaXV7Tf7g1kMUVIRqjZEMyEIEn3PkKGgvIiRIk
Slw7HOM/vlDxxdR2cXiWZ8WCK/UFt1bUvCi11aq2RChRbJz7/EnDMhKJQ0CSuRjZ3h6RiCjhjcL/
ktG11d+9mYMl4Q+9ukm5BwsQu9fwYo38gkQ134zL61Cs7WaPfU7I3/5/7n9uG33h88xQbdSaoEcK
Zgm+SRkF+VtDbvSyR+k96ojUBbOBMR+LJaKr/r/FOwce0u8q1pjSYDnR1SvlZtRcF3ILZX6ZMoOX
oezxiC9EWZMu+vh8LTPwlql4MfsAlLyHlmu/4OfSmrO9uyuIjMv54NKrgqmQv2Hct+U7NinvLY7T
VsfyXKLW2bFKech70466obm+2WzvA0oBlj0gwaaVjPVLRGetUy8nePKQx7xntUaNJw+JXl8X2RZD
yG+jmQAKwYaFOG6X6OEic0R4prtHJn7b0WrDd9FNYRdyxl6cTEofY6YZ0/Mi/GgSzmSAMBX6blCp
1l+EJRQg7WfcsCDZ76uNjTt3Ys2vkFgGMkVpFQ1SxwQvlQNj7/7c33bg3LCZpVIObUiJyiq6+Y1+
XClz4N7SEPKcn8oI97mdq0gxsk/gGDadgHiqOajN2QLHj2S+gcXa7JIxaxbtnhlJHrwUSFuxZcJd
nk+3B2zhIySx3RVtYxgmQxOtUIx5bWI0uOu0kkXtuTLsX29/D9Z5UaqDr5EBHEdJg8pT4vdYfczG
4ijR+6xrYSIlHFoBJnJ6aonxlixAQMQizpKlRbuNu6ASY0/pSnkgeVd37gj8Zzh7h4tz1LUXNth+
VlDnGVowHr4jGG9XVPWBN+2R7wGPA5ZqRPOMT9a+Z9dw127PDh+nIHQV0+GLTdHd44mkh/wRcqYz
M5Wk5CScddGnMQi14zIlZuhrtwRCmQztlNbvfUCHJEJEjic4bVk++G1blkO0XFjgmQUWyxKzrH5Z
yLj++MNxyOuNmkFNPAie7WNRJLDRF1myB+JM3w5+33KXV/Eneu2l0BeiFhMFs0y6u4STWwyUu2be
z8QcKmf5MsQf/LOg+yOZJd8FnxZyjOHNQBXFy/gBPJr3L6ngVSm6hy1eSmE/wSjctKqzmGnkiiD6
K+6Ab+1t45jdIN1GUsgzRSp2YVVEAIhGZlbMddJxP3uerTJUNThn62fA65duvFCID0Q2D/qXYDu1
aKqTG3Mm62RpTTD6Wq/9ciH1nfb4Mzi94AF3LGZIv7mGLdbSyYn7BygEPGRvEdbxHi0DwRUPAOb7
FBj2+UKUI6ZwEmThxNdl2gHU2ksceYOnkALp6v8DvQq8Pp/qwr8DckmX8/ouI14qVGNY/McOWpFS
pk9lw8HzOm3x5ELHN6nF5Prooevd8MXkkJ9onx9EsRXDWl1SAMSBTUiFKRcuW8hO/LUM+FNOEBGz
aQJTs8pZtqeemlHOA1+1l/tpS9W4LMbfTrXmbrdHXlGzeAVuGXcqL9lNKLDhTwYJr/JS7/Zu7ZIW
nQ86zru2ZkpAVMTPzFXLkLwkk6gU+vw+TqlE2Sh+kB+19nLF7rnQ30tWJ29alQqyg7JWDeIeBEru
ZhemILKlIuy4GTyQRG8Zae1llrN/JHyMp05GzSdJjUpi9aq+a0AZ/toITciyz3LtpSIZNqVSKh9b
pFcgcdtteUABF2ega60kTEYnC+GNLCTQmNfn+IMcfdZBbg7X8WAfZy/CRjqum4A/BHr5cV4zI0Yn
sylyRi3vn5FGhjUltLrpr+xJpHbF7Vks8saMn/dWbzosa3OGn2N4IrZrD5t6T3fCKeXd5cykNuXh
I2adfrEdYRRaill73IUqNnwpawz91uY88vLQWvApsTOwS0kXy9g/UlqCyV77ZkSrBID5qRszWDWq
LuSU9pa2OEDD20sdQzyusVRGgHuQpuKIPkAq8OJ9cvETrV2rKBAL2yqgpjJsXMCDKo4RRcFl9MYo
+rbKVP7nEfbMTDmoE/M8gxBxN2Mm81Miplu1DqFpH48vAXCwFsnHD+BYzLMzz0vcb49FK4PyURyz
0b6qynDjh07BVoOB+D193GtuQIizgmEUJiGa1tUVzWmJeNtkiE9TYl4ejXw5yjn6naUuruWxCIT1
kug8cHHB9AuKT+lMvUXvXdcc8jU8eXJYMU5p0i5M6YC5QKWMMxfjwAfdVQv39vbSVZDWduIF5R1v
pS8dnqnOMqgwyKMtSA7OckzzdjiK2SxzU46VGxDi97mTWLWzzVL5HwBHf6b0+tBvmMTUEVH2rdZ6
VLbyCHI93A9LOcn6VG1p9fdNUY2p0ZJ4bQ9Yit/7iLQ8oSahxJY5lPepbbC3Ccg64ebc/jtSsoeJ
sy6wSbAlVM2L3A8p7inEV6gNrPKdFaX5cNIkzeIFJsZSGHELFbmQr3wtG+LzmOchwZaMhzy77RL0
YZqSBgGBJR/jyAWCWPvd8rlysn1bFFZw5McYjMVpXiMcLbEDeZZoSJbWOH1tFAxvwUCoqXJPzai/
qgKpg4DGYUPDvLLIuKAarqs3qMmwCelksecIqhr/q3gjQRvLwqFuVPNiicj7zVClrzwzEMBejJI/
9hBmEbka3qfGCuDX32jqZlaTENTgINce9f3ibpPl+TobG22GrgvC3NQxvAuWod8xTFQu4Kn+93ja
y9hJ0NpxELdKk85kYkKvgom7X/LqRez/EP7XYMEUP1C2H5AOu/fWlfD9kIHgoW6RchgcJT1KHtVc
SY7tBHAdcXDdd7lkO+vXQbi6nLEBaZ/5/+Zr1Ew7bQJ/Ch0LUYWOd3bNMthkmBertalgRPfWczaM
2nwLy9kYOVH03TQtWw4zuQeTQ2NcJtq39/l2Lx/QTB0YWIku4MSuSFRtcEwzIJIl/1+FhKbEZYtR
nFK+EDISGJO/Ohw86az1Bceb7Iu9Mde2gsemRKh+GIb5smSilvxgD7/w3AwKqRz49tv+1eBQgL1R
wwtPie7Aq3y9BbuV0BAUbr/4gjkWA4d5TqjKb+qQ3FIQQA2tMrxosU2ty0tp5k3pgN0LWL++eRLX
T7XTwD16JIZX1CiAFhGMkjikRwJDH2MtNTOkq9r+NJ7jMclj5to85KloN5iF02R3rfzx+KUGWas4
o2VflYBx//7IODPjLjpbpaPjzUBae+eni4F7EqEJT8Dz3McUAdklgvgobTVCGCz9eAWbUQoweKJE
Z1o/wlzv8QDFx1w6YOoBnA9RuJUU4Fr4feJd+U2gT2LMxyd64PKzoSDvMI40jsSi3IgLYSXp8NOA
Fsqjy4EsF3npZvRxz4SkvGzt2o7nprIvSVP+3pPc4tAGP0XK1b8O1/B4leaF53rVOLkSUzxQo28x
q6lCXM5ulc+BDpDwgHoyVgdhryqa32QJGrEJ8C2VuEghUjSD5JrWcn000rmXEBPqT3CjtoNsQ5ej
Ipv6xwzSbRr/DV02rdHh00iXVnoJr6ZHhXUbqky7I1PsIdsdCwsD67pu04yxkZR0kiVFtTG/ksjj
gaGbNkEv1aAf3A5DnVHvD8km4F2LPAGNB5jNEee0TOCXh0zXyP3fY5bQ6cw+xqYzmaYXCDEsM9S3
AUeBj8l22jtjpcBDJwt4F4LwUG7Y1sDwm3rbmKyk+2Z8KuQrhFO7ckwZ7miynzBahGpzteAQlkKH
iQvilNStnHWNfkCUClB1iJkOsDsK1yizzs/KPLHr89gF20wBYbditq7a/4kZ9vEGUzDqiqJSHU3o
VWFiM/Z3iovsogdYgrwZoJmxkk6Km6kiIUIVQLWea0siCCeHzcL6nJcTXaCyPIZ6N0KgoD/Lc009
kUTtRvI0WRw+CLibqbjWesvg6NG6N/9v5cIfyVAjWlJR6USPAYqo8EzNhwk/FiLhadpnsvj/E/eR
JPJ9oTpCCLhmnW4BbVrK9KKs8vhWI/9p9SuQuqP7aUFNb8R8RRLdcCtfLt2KzWm0sqRfoBVM78Gq
T1Q/XgJX76ae4eYGtxQMf5+qfI+wYdd5axP+guol/ygbdpOIp08efyDhEBfxN2TF6t0qbeNyC/T0
/wLx3mHzwxFvrfN7O2l83mn05HlAxgD8oe0u9UpBZUXqldaqgYgCJZ4pIhL+W4MvpOyIMyDL9E3n
K0ae3z0lFRU1FhvE4oxutbw7EtOaqW9TTKJrc+QNsaI52acSsuSqBEXa9YdC9ELsYTLczVzJKg8X
QBiVkfbqpR5DAZFd82Z55ehhpxc9wdtHI8inPsmRnaxPFvs15YKDqB8azhTrihmPvzJr8r0g7fCb
knbQ2hs5Yr5NKSa1EajlKZif9SRBgflONxrIvrFBUi+Y/ozAoe+S52lJkDQ9ME6vGkJGlu7ankwT
27LEyXWkvd2aW2qM2oxWI66xFzAbENHkN8DZffaU2h98xvHZrBTY6r4/cugOPEviiIGYg+ghUFEC
stWeHrdANSvSBV+wsJwe8vUyfn0hCDWl7olSJJqN0kiiMA75+JIFTPPKtcPYs5lyQJmEOYzFDSAu
LKq+ho7zfUvs6qsC/CKN48sj4xZIOnkVyc7eNObSpSVr61FkkBJyNCm3Sa7CpMYnuJ3C1Q53u5YR
93p83toJCCtiypRuhwASf3J/dlWytt0kyVOVehVhu4Cdb/8ZVrPvfzpYty5IpNNyEum46o6DhhEL
sBzlKVU0W99Ma3mBSD8M6FelQ0yvh09qCuqT0xXkqoi6KBSf7xSAxcqgOnY9aqjmZQOYxvzVvWG9
ug6m0uqG0IvRfdx93ApHNwpM7PU5uSSGDefJpDtUpyhd/DMfzF1nc2eyugQb22Jim4fPya0DwLZI
jVNsUCmoAckgf0xgKie2tmp7Cz8hSUw2aZsKrRsEDWGTYiqHyJr2abQCSrFXo5mxZZ/lF6+49kwl
cnV4xOINJtHZ6Uj804D2PSOesXuzKm4Dsmj9Rq/lZBUlu5TH1qud0uJMqKnG4FJOvGZqJ88kUGgH
r8AQbH7C9fOijPIOhVfhUehqQmZ+clCU2JiFl9ykLPNZ4SUkrCpabvLsjlzwkuJA/i/Qd860BMnV
gwpnzFHmDRm5doYvs+PnRlaZT7dR7JtEfU6Zgz++iiXRblf1uzIIMnQxqdcwaYboSUTZOasR66Lf
gPYkzjKR5uhjSuZ9WSLzCBW33pncLr0wu5hP4LNxVWlJob+G+87XKi02YT+3XAWSqjl7kuGRa3/T
aVo9DQC05aQt7l68hDJunjuaIz18RiF2flPBSRhmx9AF96sGJxdBVLR38yC8MFjN2NWnl983ns2s
RlcjaAi7zqHxbS8Pe4rFH1fSz1bsC5iJdc9hG8jpdnHchlvnHExqZnAMJviflynwaQaNnMuCob4p
OSVQrpmf0w+EuhnNyDiI0/IVwgj80rrJ8EzxWGXpelD0ZdIsy8Y4AQsYZexiMemK+6vGHBGjDvLB
KQF/gJnEXqNReY+VDfH0OXekILkzhFzLsYzcZiKZYIEzCPxCokfPkuRzlNgN6kwi0NAFIpou8RRR
urs12YOpfS2AHkkluvP0IMNkvModiuUKT9ExDxH0NtsGWwdBKl++yvbYdlqhgHoVD8GiPJoEl1to
RF/gttV1w498OzP8F62lRGGabHHimAeDhtPfAeGh9fmKTUFoiqKG+VA4h8kbo6wuKonlBYjR9PAN
RHwyRstO8HbhpmgZb4+EY49JOkkPjIhhvZNasEPAubsE2AdwsdekrNU260lJks4A+vtAIdCcfmDG
TTidGYe4Xr862XUlDY91nab87shtDR+W2gcO1Akb32WHMYgucVaSDPPhCkQmwCFZ9HH7ACHs+T+l
57U3VYnrItua2Pqyw6BRbQNzPaCYsxNDt8rqlRACMbvhDHKZkVsNz+JTPsmtVCvG8CHEy3nuRmMB
hk8WaYlhDrNnv+Cg2uPWbBi/UOfov8kmUk6Z7xUEPVg8EQbrYPsdSkJfnwsmeW/+zZrzhFGpBl43
2z9m39+f4TQZ9jr6WgkrbOzevnua3PX1LFMmdub5IIpqr30a0fMBEOV/+0El61AC3a/fKCthJdGM
Y4Zq3nHiR4h8tmbT97QWeGP/1+az1O8sXimCTT6x8OtN0DCpJWjCLeaEHuU87tZvJzPwlZM1x0eE
dEKYGFTRxGO8PBuEE1r5EUylMs7GUVQnxveYle2Lla1iZxjsS0coJs+XJJI0aLMhLnJ3PR5vNZtV
dqtZQywn2hkFpq+RNk8gdSKTTC3rHDKt+PPt+HxoSvbxT0vTrkK0ift3vRaxRDGC6DfnZCkoLzjU
wjXJWIcrhnck+IAamdZzdis9JD45tI8Agfd3Y0u78AngWfd8Ggcm0wzscoVMnkSPLG/M8hkrh+pI
O6r/SEorGyGtt9AGc0wZwPj94cLZ/ftkguCEizj82MjoO6emLveodLAKCSGavc6v8wRlFfClu5eP
O+Goh84tSNyPG0WYtKHyATl95lBLm/HLd4Yz3ymuT8j7tC/SjiyUOBafmvGEbb+ejLZJHB/nImm8
pDVCUGLMwLWHsOQmmqWTJt8lN3Gn4xc6lAh6hnd0asRAjC4O+CyDrrrW/q10tFsVBH3RO/PmacP0
3UnpxEFAPLUvmpWpqg9044bgK6wRV6dP1dWkPNphCFN5gOV5lORuH50wuj3BQonknJe6YEM6HTxw
aL+iIM1qnT5BVtBnRzipVE41pH16REln1x3BjY9XpdCflQRqQoXIw68UKT6llikvJEqbuoA6OjGR
ljqWZqtn/zndGVJfMnNhvKcC7IIl7yHyt+74gukybGxOHiX8z4kbQSEqzZGOvfZpmcgosoOkaLqa
9zoy616zm6aQmiAkhYF7WcKC8E9VDj5k28EP92OmjpyCVc9Jq/AZ5pViwGYt2BIxRzwc4zOe2wWl
pZU5yfB3WZ6Z1hEZfBLxVA8mFewc/P3E9GkT+6KvPvfNVbJlVeK13V0jreEOAkp3B3XiPJ0NKr0u
1Ugrnci/oQfy8IDoHDJ5zxBlpTrOxv0vP224LiqnQg8j1jhUpx/4R9rq3eQojTw2tabh+2KyG4mW
TCuwLMqxPc9QqE9z2d/rz/IQEO5L6B2O9y8FMdSafB5QBiocdGnTPFpnUCKAAxTTpj9ntKKrlGeS
TbkYHWIaNwPMrgfJThFNI7uzjD+L4znD7ozxoqfQ6jxrzDEltSTKYhc/n9z/uSMg0jkF1oeneUUY
kVfJPOvA8yruk1Z1vsdL5KrWAj6V7LmwUSOdkrH6XiyrTR4F5fVGmHFSlq4DKiBStK1Uq8KrmU5h
vdj9JbVosKPhm/3+QMgIW5pDfEtRzVVNm78WbbdupHZtpmecvMrwulc1AlYjRee89EWXP92RpNn5
W8XytQpSU0nkTb6eUOqfGtZii9JEhC/W++Xh8MTz64xpDViSUH0AspV3tkEMM1c8d74A9ZDGF7PW
yuJriIq4qPwLvt4rWdqSh7cl7olUEbOtD3ljfHt1C9ZxfG0xdhToFaV7H0m+z6DwoQEuH0XmnWo8
8WM77lQKYuoZU1W3sqZ5o1T2nAI0jhNAef2I9lvYzB79D2+Yc7qIRwfIxMCuFmBmYjasAE59bJrs
Ycxa+1kYogHjBa8ilT+HmoaOc6D4Y0bqs6XmTpe3JAlyBVo0TWvmzHfWE3xqAT6GAAOAQNVUkSg6
klZwsLPoa7WxAcm6c3clRFhSmjAHiss9WAMhPKWTuzw2SGmXO3tNYlAm6AaG0pNvOBxNvZ71LmAF
U8QQLMhNFaJmC1BO+QKCgeOsqwG8HohOXcQgAwQXChwKt+sxPosMKie3amZP+SP2HPdZ1Ia3RLZc
cQM2HQrG1nUraQjV58TdeSq11g8XXCwocVH5Pw07lV2iEVkttKRSduL9MA0pXGbr68k99d+LhBMt
ioLNtjNFHkwaH0T5hUU1sQaH7g/W4hyZ1aBCQtzSPuTVTd9bwjH9nqnjGtHrJhJ8yZL0Xqr9Q6mY
Yc06sOG9dLAoaM4H6as/VKf6yuUKb+Ayzhsz2cTzbgQURKUgFh+jDao/vFyPYMTDX9efjc2u9luy
uR+Buk6zPWiTechBULIMAE32IU2v68192zV93d+tsKHdHDFE3jYcSu+StzpVWulrd2uGrB1sEs0X
kKds4qN/PKurs8UlWGGPylE4JjZq5sgg5yFyeFEE/2V9eHeECyc+jpGfDgJF+mMY5jFy3j6YbkLG
DjygoiEi62nd5zyWOrWX3IvyUHzfLNN3zYncd3Bnpd/rjC0zhH9DqyiFrkDNnVhPTIbE/QB0xYa7
RFciDdUapPI8hCHG130SRh7Ez7fnRLat0NC3zOZMXCjgRK948PhNhhNBi5Rv8JXEb5A9GCDMxcEf
2Uyc9F0MEaQhfjkzW4TheFXTqmo1EkhwBwcy1p1a95862/7lJBKBDPQwmbXhbHOkaJC/tBvOLEx2
CaIx5kjFyumqUIFYdTjKj2stmtKP0vkIfV7Q6BLws4z5BZwV6sUyDEDO233cAFkKvUj2rLO1DFXx
qqcXVrbY8n5dtsAApdb2y2HMKeBUSg4+zsX5T2xYSgtysHpu9r8sDgKjoSdzKEXEWKUMu3AJrRWv
PZFBXUXGFRI+/TZlswxhAV9E3lYT72/nCjdlXcG2qUrwpKxABk9vOeZI33gtmUXwkFcokvYCERaR
O3PsFCRW4t1vXBKH1mX6cCInAWqfgLBXuPsF6Dlg+nZ+jCiN5orfJkdaNNgagdnSQX7SxTM0aQXK
BPQcT+OmW8i7dUAxTJI5dLf744CxL2vvcQ4oSXV7j5uZeyyYM9TUPDMR9vvCsiM/9fUyFV84wWRP
bz9JAbV7t8cIkyJWw3VpS1MnLiEzehik0fBRt8WqrQzyXbFd0SoqZ9PexvgeuIabzA3g4zBkidBr
fiEnC7gV7IkuDzcdr5k6lOXHtx2jC5YHQRG3oOqQoyyis5KdykbAyIp0ie0ONB8jdB57tfH9w3wK
SQC56yArpFI6b5xyLpOtRZP4m3OvdODCbVxXvlLOttWyC68Cs/E1u9DKj8+nNvuCnsoiSNXV27be
Y1lVOPMtdQ2IHglI5bKcJhgl71W+aOMWqDseSjzB3OO08Yoe0Nr7DY6eXtf9l0x0OkxiQVv60OOC
pekH9cZEH8g3AbsriP+4VfGqZhpzFr4uvkedeDhpDmX3/dKoswXOWQLgv7puMkic/sG1mBbSJpgx
/Et75jUMIqMF3vsnXs0wlnHrHni3/TwA1pagS+taQxeUGs1YANrnelo+WRfHakAFBYZPxSQcgNG/
kzHrWLzhiN0P9hUAH1JqYzMN5P4bll7rN/PyGqpBHFYDV2UcBxoaPNRHo7qFMMbYT5wLhUx0Zckb
VSKxGjRwUTqDblbNAVryk1mbeHRgsrIR6anSjvvzXyDIjAfmA63/YcDZOYUT/E4z5i7afGonEToY
a8AFCaGMogUhirtpJ+bNt19DVMgviPs/opKBTGnkLURqrqqbeF9BXJbxSbx1UCOzsVLkZAAPFZOQ
s8Oth0oLenOT2NkBDgT5a8LfeD9kNnJ9SK0ku0moZRn6O9/iOOlM1gDzZaWVUmZYpiVaGvpirC4X
ejMHVduvJOQbs1asjeRmJcGsgp/+mEufR/OZTKi/2Ej1Gc7DvpLqmOgwqF42jq9+qIaxq0hZNuIX
S0dJr5IchJPMAM0BRERz6wC5vT6AkNuG3yGR2XfVIkG1krJGb2KE6EvhOtOTBozc14giystmt5Tf
wEdPAgRDjsjgW9pE9E6hUTEW6724zAJGETK8raV8eLLhlNWuu1F9OCPB2crvokTQuwsvY9KI4Pja
PiJeQQsHstx+uATr03zp/jSqjuTx8lk0qTLAI5Wo9aGm3MfWCWP9IzWZybNiRTFKJP94WRdYxP8V
dQ8bvZ6U2EDYieONh04TMEGfdT9rITWS+4yoj0uOBboXw2NsfhyNKZKc7EmfV3DooCe3i2RUSUJb
YhPqMGiIY02iW1nL7+yCEb81P8TBkynyB9nCvFBxqOIsSGSGf08yYm1QIA671KSCHETbASP9sM7c
L5H2tfoWTvQDFZGunhk1bxQ+b2A3lInMmj3uGvrQyzWSKMp5xBACjbqcyfMSnioBkbKoDniPBdAY
Jf2KMiInq5g/nT4qVNs/P820bgAqT+KAJF6UkvbKHFMM/fPa+PGeV8D1cn6I4e4RS1kxgrItMf5r
5GAckNd7+dWOBLG5eMJiJHtgZ/G+I1EokrXMrVJlhdxySuwqyvCWpNSxNd7TSVJMhOZQSUHiSZdg
ViiFu5iUOL2Dokoi2Syr1XgJsDghFvCRPzVx3yOAljs8EJ9but2s9pAv4t9HyR4gjpYXCcfn7hq3
i7pqj4o/9WCFO9y4WwejTeh/iQTvVBD9rrfg3WMrHeC+L2bnQehWpDkxfQgn44vrRXu81KgZogoN
TAgGxaoT0HPEJjQOhYz6w4OMcNZSZbUTLE2hyE6btEhjCG6CzSkDlEdwsxpj2In8BXljdOYqY8Y7
Hw0iSDfWNbUrO2cfT1fJ6JbunFKM4kxGIgJ9lhi3vYIz0eD9gWRnyeW1jv8xNRpa3s+4iz1xj+TP
YB6Mk4ZuaaBZIV60ABAtdWCw07JWPeCN0VmKzxGc3PC0OXdbxKCTdQHsuQZ/xuQUX7P+7R8/OeaK
2AJlWEQi1x36OVHA6jpapxBgMObUWKa7HaZDMUl281oh0ozKg78Lybz5nUkUjw3FwaIy2mY487Jl
HTucaLf3kY9f4ZpR5HcqKnLa01Jegu5zAcUc/SsCbgV6AsHcN6JR/WVGuphS33X749wyByFCSWtX
yjvhEmpPnZH/qjRlPys9KVC9xQcWSx5FxD/aGe2A76g1pUZEz8kLGTKz+Nr9nmMFcwyRFeZhf6XI
/FMneO/X22Nb4kgXC7jypWQHz9n38LDYHHsA6KLctuRxn/RkJMl5eJu09ehnXGx70M9CNCqs94Zy
AUG5dX6EX6Jag3WgwLefjLA4KkE+mCLWWmqGCU+XJEcTa38HCJQC5+7NbPLz0OautYZ9NDC4wHt4
L4isXn5foD6BMDmkC3YX8qJhDM6kXze62fPMFvehpQfsOzVMpRIIUCh1QGcBDk0b8383QOhW3cBp
vYyLCYX7AXpY8rxw6l0s9jozhEgWCA3mSG2CL9TQcDBqZPli8KN1TZvLAklTgP0ntoOk61/ia32d
IzC4AXnZs4uPYW3ajburgJKCBrKv+DJDMmgyvmV+CBI7jBsXIF4RrBkK1j+IKlf3JPkqv1CXu/IF
4xerAFLoRKu+ekpX2Y7c0ZXZ+ju1Yahs6/aS+YUgAkJ3N3I8D6Da93AHkKtMXRF6I+7AvjKEK9M0
GcFTVpuIi1JuIelVyJD0B50uEbpFS5Ptcg5/UQH+8szsatjbIZdHHoNi6DGbDlJJOayOVuPRoHuz
+gHsYUKQUV6msvYPwWgi7BmhpK14ewjZ0TWx9ZyiK4Yg9yZMnseuOoNTzlNJUzsrollWppkbY7ys
FLXdXpXgUrHP3izy75tzujfFLdPxKLLSgzpy4XVDDKpwFtKkgSe+CZVQmZqBvn9S2G2IduElhrF/
EBOBE2O5a8VRlIpMj7BHpAB41d56jmJeJ2d2wwMZ0/d8nKonhfVI3Sg1TpSg2hMM4tvX0cJOapVT
1xiuvh301C6z6EidD0+M/oXVAnkzFxUCP2PeN+eTZIV86ZGTZEX7aA8msKp8+WrLWPoLlSgc7SFH
YzFhffG5+gYkRse50MvILNy+oBEkjfgrqHyL4SYQilBMVC538KGjP3mWOtdhFqdXSpqmIggm8KGl
JtsjeXBUTM0Va/cnTp4/oaFHNj0r1+dJ8K9dfaielJiOZFRQ9Q3ge2EqBgc1hveSE6PDAU9pFp7s
rzvY15tJNcjsnfh0MmLzRp1JtWbRArOos818t/krniwqXXH241MRzLtYSWrr7gA6RAwD3wT6UCt4
UFBmS49hCWSUiDM0hID0TDi12uCwM18y54CQzuzTnVKv+5xJtOthvlIaWQ8HwCXEA8H4gkhCOXbH
LoqnUspDswCbCPXhY8acDldtCk05LJnTb2G2NwQyY3dy3HBrnLOmLdBS8IYrrUlMb+7NkJ7oLWaQ
OqQ9d7PfJe1K89j8pwq57hOfTa/1Q6EaAB7hfU2Glx2MYN+4l4Bbba7EZvpWOP9ssR1h5MyAK1YC
teOtI68s2g1r29msB3HsNddNLm8x8w5YAa072QVwKvmCDeBQjqYAHK4m87w4QAaWgiPpmhNurH1F
nAiYSE2rjogPh19s7/W9PK4HUKmonG1eZrnWv8Yzcl4rtlypFw4HcDvMjy/Kzs2VGZWxDEII/FoA
QrBzC9EUjg4rL7kXQRFRIX8zW6ySrnE+Y78Zp4s9NSeDNKdk1r/1Fz+7D+DF+PJ3IEOjTuL6bJCT
BaolZ9JIc6kHkdBqw7RO30DP7UOBSQ1jtYB6fOzTvkWGp6x8JjpJFV2VOtQx8yQv2W3hZlepkieT
5kdO2anT72nOP3hG38hBO3C9ZzoDdpIbJmld10b5XYdiB79hlP6Ja1v+w/hFfu3ttvEYgv9CVma9
YxDReUu+lbX7EJdm/S1U+oRf7gr7QDBse/AxGvmQe0kS+GpEaA1NCG57OAmMpMIDyHJnlxec2/dp
zIMJZUrYFhitkAPWSYZ1VHvNRigRAHyjaHDROih9viUVsLlUiZFAFs8TsQl3Fa/qjXLlwwqzYkZ5
vyrZTQR8vuAyAq/9BCZzmzKDcPiF+/4mc9LHtwy66NgyyDTVU8aRVauaE8hR/QsKgHGitxIqYC1/
xL22P97pP02fVkhIs1JkFTDnBqURohi1YB89iY1Y4xl3mpSK8IY+DyFiZtD4yb4rfQ6GCLrVtF9c
CKkJUbG4+wnTfmXTX9ZCkYvHj8min7c6wHkIv+XDsDnzcJaI4TvtaKAa9g0PBVkr24ACTfXKpLRW
FnwBfPX02D3dd50Fiz0liOzEgFtQElLJdlalCbgUtoIGVqX6a4BzlWq8S4AE14h5NJbjhlr73xNN
qWaegQXprRJseTqlFiU2n8Tv57SX9Rrr/XKJY/RcpN/slebA6Dv50/eLSFaPWx/bj79885H10lLd
GZ3lQxR0YTKb6jWcmSexjm2vf2lFqmHR3hIFx8LVeIg/CtiYDw1oVdq4+4iS8jv1+uvJlbShFN/u
/0u1h0IrBCwYIaGI9RxMJxKF7BkZ+OwL2J3+0usPuChAzwW/1vPYz7PayHH+Ba26cT8uV3aUDBrg
KktB2p0JtmvmGjMqwvErCWBqnANddhCg1mkYrANqdFLBkf8VTBNlNdmx6DA+QCkAb/pYLAgFmoDY
kw7/u5hlXDo5+2O03qoYK6l6PwsK7PGI9HA7335P0c33zgilC8YbAB5VvNXWvGWoM+y4/YdsrW/A
YmszWO5v/4RpIc3+oLIHDvxSgWemAgYg00mLcS4jQDUaujyKfeU0Lh1Jtk0/5SErirekEOm9tBXi
jo3MReGzAiEl8DRrhGgocndk9jUIR4VntR3/TJWpZ1S95EXNwknh4225e+4sZTmftRoJ9jTsjkmq
ufan0TamtF/Hy68JGDUwkUkg/OqArOUHCdvGxyLlj+B2YKcGYqseburbPRwhJSWFn7YxaIP89R/W
mSDvnJERDItO5Vox8pFbmZvnEWYmfe0yjYRyjsGRy8nzTlCk8LElQBFf1oOiW+rGnZRR4VN88C0p
5KlNsdb8fWnlJne7UTar191pFceFwsly3Z7CtGiJqX7h+G7y98rsV/ChQsGqDKIU4/oO4vAAHqKl
gVJ93FjCNHKD/SUgstWzM3+aMURnynjKQkda82Lifv00w3bX5WopfVDDBFNB24MGRnOtjBRU+fqF
529uXRmR15L5WeOurKSKhuC9lFTJSshGTzBi0fQPvinzbXWyWguEx1fMI7vRVWhO+TcrPGPL/Dp+
1GqVH/0SunHGjbUdeH6dLaTIlfyvxEzWHYTHWBaSQ+VLwmlr9GyuoxQ8MRz8P8Edow30tt/IvuRy
0vP2EP3fKA40Js34MEkEioOaMFngZrTUUS/el/QfjKI6AsMIp3VjSGkFH6sOg0lCh7g4nt6vaiEj
e/vKH5GMXb93aeo8ZrVTyFAP2A4JvTyL/biRAQQuFWrx0J7idQmv32OYfvEz6Cf/2OesVGGrB1Pg
5STyaTQ6+8ymHC90kuJx5SqXwec5tKoQcqVxQBrvKPKcpWVEl4EFTtFfU9noAvpZqhp3PCQwFOlA
Ol5Gp0w2FbJpZ2LsP/MfvMzE/4BeCbmOMVHWMo6JRUCeuPxBJCyXeWmbjyvcn86rQaRtkm2AdgKL
D8jo+h3PLe5YrakOqkzqwlBXstBuUrkGSRCRJbsFyqa9ux8xyEkp7sQW2qzHdu8X8RdJmTA5ZD9c
TgUriDS9J+mEJCb++gQ13p593fmCb4r1gQFClGgX+6qZ8ZEcv1jumG6EM8dkeL8GPHVMXGI+lfao
RfVlxyCinp/k2jx41C28pfLJPGhlVOqRfpfiiRIdbO0ts7lYDF3QhGrHxTUzUgfLZZBYHof6HVnp
jMd4Ro9T0qXBLFNSQdWhpNRS1O5qfQ5pNkkYq48r8iuAx3kilenJPH8pqT2nlErJHAgl7tJdLWCA
CrM/3Im7gn0neB3YUFCi/NarK+wyGeDnZqG7uYrGUQg+QNX+dwVeBm6n1kYnIoIN3CiP3+9yCuzi
WI63TBnxg8yQco1ZqXg9+CPg9oSf1/AljKHrX2Ky4AVdQ4BLgUUyQdiryAWhLVUxJjRNUxHHxLB7
o5nhsM1CJrIboZf2B61yN+fjhtKR9I+Bi+uoi4XJk8poz/VsNyQJqJTWNd7u9Un9KekpyZ1etf72
jlE4KAKBIX5A+4Lr8mmka6UMNtY2GggQVd6bYSjNxn+pfehbzEpeTgCNKP35Ev74mNWoCvcmx6ZI
RUVAMFOlb8WRFN0N5KBl1MIoZiql3RtymlxL39GINHTZPsY21QtaesTtCGejlgTethKQyQJFjYgf
NORrdCS1HmloMT7QS4luQpT2rXT4N7MYXWkt/RoU8sciunmXziW3T67V5HfPqnj11uPPbmFIllMr
VWvsuyDkDPfelUigwPc+M79SkvHVtNxG79KaMqGpBYnug4aky/ml0KpHAo/KOSEo0OB1vEfxxGPI
WFJr7fvDJVv3v+neEt1AljfQeW8b0EeDz/zQLVy8nyuc07b/nkuJgUzGzog8SGYmVy50xkbdjAqS
DwCShGT6I27tGQAeu+8Tx0jFVci6L2ezH80ZTR6kFk3moe4MojOF+VBG3KFeDx1dF2NTBiRidmfg
OZUY6Gj7I0cyzd4YFckFURskrcmBqHQjQ69XrwTGBtv7TcMNqPrkFvNVq6ugvKgIZat8KCX0N8Wd
uIsGg+fDKo4GiixRY3JIpVsuw2Y8VgHo+MFE+OWBMxW9NhHNhMDC5ocdAM3JS31+USixjM152op6
w73YG33agUdV0K3JP2r5kweocQkpDb14ukyY2aOTINNGmA08QrX2MJ+K/CLMuMpBbf4D8hf6OAcs
Exfo3YmlIb4TcRGrayzGiBAmj9V9w50mrZbHEKAHYSgXrREtFk4MaNlcciZp2FyEsvgcdYZHL784
KGeCL+zh5Q4zpc/TFY9Kt+EmvbQ7QjiwecxFElEg5dC9uEu0KcC+MJEO/wnxAdhbUtENWwvnYzLI
2jK0yQuQriDfGp8Zixpq6LQGDv6NsrCvtJpufQYBxrF5SP1xET0wtSsVEfuA8+j2Pn/UvZ+8x9eL
ojs9k5C02H7DZIvxouervlzbaVgqb2P6HaOPLGiYHfQiTlPcKErrhqV/OPjRHJUOcxTxPsHnaXAq
2MnUmP+eaZ4eOhBtxjtC4IFJtdGfMPjJJifxmpiXyWSSILp8zPuPkZHoSyCRvZ60oNxBkZS3NN1g
4/vScfcBi+ah+NTHrHEkq/UvjJJ1EmaaiDJS/XjAfp+2PjjkVhHS6ESl431UlvWFddNkJWFKY+xT
XTPYpG5rWKXvNG2pCMdAJ4MZJRdrNs2xw7172OoT9Dn67pEe51laAr2Ug6BcsmpA4DfJa84N2436
a/8uXGijwR106huk+k1yMcnyzd8y2Ezi/ncSF5EiqKkRzkID2gBjtX61w6qjeuUKvkCnt6nB8rBR
DQr2Pb0byAfYzGT12fRS3XcyQLCdkoygSmoiK32VqhKjpq+dTGL40gN1hg+tTAnvljtBaa1tWWUt
Gxa0y5Nupca2kADXRIuLikAm1O8zIct6oDmQn8MW73GQUa5/YXT6xCBrllw5WRjVA8u86SnbJpbU
uXT27eYjwwOya3Dsbp7p38P/FcIDNgFJm7wAc6Dz7JQ7GXobcmfH64XxBr8Brzz74NBsU3HjaxPE
BekZlH9drJLMiw2C3yXg63Wpuz/TvYZFgB6Mbdy/ai4hup2hhoWa992NedOJ/lcdxXE3tHIEi+xB
LyMf76ps3FAyLbTke5PnLi4d0bRhJPS8uQqKwD4YNdO1nUXlVNZN3Fhn1GKDEs4HzGqpvet9uwEB
FpC/1Fcq1x+tnbFnffxvcbJuT4POLwgFytonKi3VAd4qe7BI3RcMMLB4j1uh3UC8Jkh8jGJslYEM
AFrkxmreulOkZQk9/ss0jEm5uddt9VViuiwi/m78/9v1BbNNu6WWx0zNc9UioiS60yLp/o+9uEKg
PvF9q1gQ1GbEj0UUS0FY9Pe6SSOdIgsbk0X7k+IvKe7Ft4bQftbVXEBl86P6sDVGC+Vz6oFIIE+l
2+nLnZhJMEIufKyVw5vLa8X82GUQUV8zZgYfT/kWVHAjVwTGcyV1sqTJPFQQt5EaoHO2YfJHSNXC
JaLd3mAnYBgLe3EPqv9kNYX33kQSxlKPET2TGNlFmFsV2iwG68Z7jvkpQIG+8UcJ1SxNa+2njyDA
kwbsg+UXurTFL6cOv+cgdAzmMB62B45XGyi+AeZyG29HGH5Jpev/uEEk/fmaRnq2X8Cz/0vJfL3w
IAUcLJXrdlt0MSMYx6dZaSgTy4+3yvFLPJ8117a4mf63mZKop3hjXRE8u0GUslzF6r5XO/PP27xC
wzwwpR2mmH45eZN77aeNCwu680dWEtHTtRk0mj6Qv80wR1J2rXDocfmW3DCBiTbOcR933wh1BLMq
cFaamMcYa271uggOSQ1iANy/tKeUCjNq/dHfi7MC9l6L1oBEq5Qgk9FHhbT9m28ShdTTDttGdrPY
NtEYBvgNuxd7YiJU1z8b7lgVrKlB/c7s7Swj2TDNLyaG2rxWWHcP4Ux5UhFbJlyk/FeXypsW8dWY
zkS1cpMKq59d7FjxAAvt5uLf04j8hOmD2atef2BEyNqieNUQDIO+ZBO3vO95agi10SDHn/m9lJju
ywjjPhSdJ8ZZvq4MAbrw/qsx//rwnhjZQ+bQwo9icV+RDUFdUZEe9uFg49dae7rmIVykxh++1vqc
7m6RPNO8X1iuY5/BNHhbkHE9FPEapDr1C22nb6XUc/91jugb297c4Zbg5zt2K7fMpOKyyImdZU+i
a7IZrpmiakscmFPJMmQuAav1SHEAPGWpPkF4qilW03kzA3agUv+NfT5NVMR2gYDe9EZ0//vOXTpK
ITCbUgENQtcVMfWorfUlpPbb+/34QLb/6gDpjGa27VDH9mVLivmXA6ruoL39OSVUoSEWU5elwbXP
vxYsoDpodfRQYipbeki1xipMg/q4zh4cxlXnnon8NBdfL6fQffc4JFRaMPNDRyNJTjbSuHGYAjlQ
t6vliGTE2OUdbQdKvyE3y+0aezUlOwcunutA+aFcD9oocPEiWD0lLITlV/3G9b7bEZYzYO08AZWg
+aEsPOHSe35DgMlN9aV3sCEu83eK6ZlzPyQfmK8Ku9crxJktjd58kklYQgZAn4KEOTQYYLuC2/WH
QGeUBu4O3pfZDEDctfaIjbPRKNs1Gj8OEL+oOs6LBqqrIQ4HYZRSDlVzSAOJzjwicK/pU1BD/noW
37Hl5Yly6asQPNvbqk7Km4WJ4BrzNOKsZ0gVkui5ctLAMspiE10aLUv8pYqZqDZCsRY2nQDawv5E
6R/LPLXg6LkLiI/Pkogt9SUUnxTqpnhmuJFbXm/qLndqsfnZkfcn4YdTNRyS820TqKcoE+T7U0yQ
mY2AoKhvbxcc4OzBDdyk2pOq52OlX4mjkGd2r3XspkDV3qKdM4V4oHdO3Ubq722ylAwVAkuOJN19
h8Kicpu6fjdrie9OlAI38UVtq3KpknaobHpf6FDC0COVjyomXZktM5ElCzAsDUuJYQ34ao2Tnow0
YUUG6YTTeadFOsGbO6+WEVi8Q+JSSIKlSC+UelOQtjiT6PKV+hUf4YKHZ4WGxtUlGJCglHqPr9Ky
ZLjlBioMnZQO+p/iCWJuxqEbKhUjFp50aVY5rPfoWVMlmBOn3n92BkNNGbtPAKBKhZPqSmTfjI5S
bFn+bQndLUuV6W0t85srZoz02QisNewXNoXZeiFuPVuRadfFLKgYD3Zx6c4d/ljUTxDkzAoW93cd
zJj7qQWrXdfi1lI8Rw+1kl6uoqPMYJ9KhnFLubHUa7ZLqauaFU/JRPm6fJzc9CaHJ0hRdlraIWPE
WgI6hc/bRmPk4xWP5W+TUmUbukXWyfAiq5NZGO71lLem5fcycW//4FvTMg4zurQaGOzQL0LTL504
RxUYU4NgbxpHEWgtEZFE5WQJ735PE8cuVGQDM8P/8P/1nBJmmEFNy+r8yb23myQwiGFiZV6mgP/c
kO5ako79yWISTImHlSEUb57DTBcCvMi7Pp5mHYtlU/MblsaO8xqAtTIjVyksg9oVLNdoLbtGdUtU
sKVjVrE5f+u0ppIcF8UNxMQ/JhFSe9bzukBmNxduOPEYb1e87vSOr/KemLQn91SsCZIUUIlUbwMm
gz6AQfolI94LRz5RfBLp/Rxp6bMDAT47o6Vva9RALbz+4H4lR7PTD2y0o0syRsiobvO9WyakxGRH
zIuDe4vCsgv1kRt6WaUutwsF1Kwqa1YzYt88Y8WF+9+t/wS2eZB2OSN3hpCdru2ZPpYI6VXxxHWr
d1rNwu8DN+fCWqK48h7/mz3THaWfUBDNRrbLoJPRlkWaW7+VgHStoRB3Li8xkI4tRqxRiYNPTo7e
xgiI/e266fhwtVHaMQN8f9t/3GTXuEad4sEGefpJnv3xRZTKo7tYr8OTVLU3WeRwUNP2Dz16C2dY
MUSd1wNO7SsMCNx9shKUWsanFCJgFSSlMo2SMnroZRlExr4Pd6ElklLDTuS91hrieKMfyzhANggx
BrcYJVWHqEzmZrMyRTIUQZSr29FmzyqAffq9fotjiQ93BgrPvB++gvTf0XH0j6on/LFWwFjDFuPg
XEScAsXxGjEyM+WdPmrX+LZn/78852jahpKm57Oo3Pw+RUQrH+v/Xm3ua4XgAFgkpNlWoA4wtvgC
0b2NMYVILTYqYf+8JiEdKxEWo0rUSKjFBQZp9/uXc7AiwNgEjua8XDNmlPr0WW6EwSX4NJrJHQmo
8JMNoB5cv8uW7x9zfRPj8hA1SoaJ0pB/Gb8zg0CGm7cQ40fg3PGQzBIyTyfdDc6/mh/941XsifGn
4UbtTI87qf72KrjpHLUJiaioOkphV1B6BGx5PhAHgczPp5c8Tdl3RugHPqte6MzHY3XI2lwTfBWq
XMklexLGK8OWj2mJg+yL6EaHGzWSutJ10x1Lub/mlI4Mj22/5IQxqexHEe1zMxevZsbnvj/oNefB
O4uA9qrkqbl713APf/XP4rg4mZWc2p72U+L4thW9DAsU+sVv28aQljh5yzH561zrP8Y5TCQIJryJ
byWcCIcaMBjLdw1NDeO+yyIabsmPzjHp14O+LQx+/XuAHoIdqgfQ2oDZRqVFftYIBvDyxtkCIb2k
YIEPI4VOyzp3Ullbe0H0KFTPtin9oeSRj/u8gQBOIQaP9fEa2tYvpsZIAm0NStmECYl72lFAevyN
DrMKVr6icaKDXU5dVqsHGcY3JXu629oTn+8cNo92fTyvlOop1VfQ55IX7m6xrsKyqkZzwIGXMWwk
lSsPBQeeyT4FoYW9jGWlFj5l9dJXviUzQg8aMTJPU1MfNMk/Hyh+HmcbbUrpW4rVlZ6lkaZPFifs
2IvuuhrtW+lTB4M2nLNvE5fyN5Gh+3ftb6blc1l12kPQFOCQ/uMs7B6bnCggKxZkhpJx8GXHUuZe
qH0qjWNCQzbcLP/la4fPFM9ZFCUjsTCnFLVGFrxw1bH3+BoJMenlIwJRNm6gnxNIbkvn/7oNGu9F
4LRaYv8mq0uZXrZRDPHQR7HdSplsewrmLMSJzVsxiWpRy5u0sFknOoqNww+vJOesb5T70ENejdtA
Dq6FLjs3XgK/s4r8rKJD1+b3QXsmdVz5nNKnvpq4GCymqr3S7RntPnpcFx9q9K6pyhU0S3d4CeVe
1g/c3+/9s88QfMd/pwdPtUdSutbLTdDRQEIGVQt5GHIy33lu5lS+yCR00+7YqBs6e6gTk3O1RHOD
BCuUO1cruoAZXJBGSoWEHsMeVDN9J2UmNryaj2A0AVBStYv0obMfaLk95a6EtCj/bOQ6gTAyn2ty
pisTXIUWEP85CWNoCm0vqjer2ltrjj6H5zAq5/KWB1wWLGScNH33Pcn0Fe1JQoJfAtgZaIyUPR9Y
kZtW8G5NSzemZAzZVMfkPT3KRj/yIL4sgZRmBnTVQTWybL59a4daY9l8VIGYo2LIJBebNGsgxyXa
jy6f3+5lpa5yZq3JBAxUKKf+9AW6oQ095+VEavTsSj+xlXQa6Fd6CGk5qI7N+dc1AFNQG9LQJkTo
mmVUqzJ5M3ixoEjNWEBt/yiLiz6BoGaTVoIQQfuL0CQwdncKFRD2GisWt2JJMQ2EIZxihH55V5hG
070oGzboayAP9XOdBbV0XS344HzHwSCFH4TkJJcLE/PSbaZwu8b33HIy62WT1AMcX76JyauCJSEc
g+bsHzGRr31zWR6OEs+z6gmncJORtWsdUdag6Mh+3TpYohIY6YT4ob+tR6WsjZGSuPlWlu9dIV+g
Fzh2J1dsUGxu5D5zA9DhiIgR4J0dXfjHvdbCUvxGp/BL8IGYA0Ik6WBW0x5/DHeEjhpqrvZnyJhj
Up/gb6OojNCHjyOyS8R0LO5azpVtRvUujEq1nD/kY05sko3j+UOS9zjQVvcRDDh5rWWpM3m4pGLn
GHp+O25XWEXYt4eI4X+TMrwyRqdc2jdiC+2j61H5n9/+G/1xy5dtYR40GtIFGXbVVSPgly09r6Eo
mlvnMe0WuK0L1++mlya8sKXB6CUSZJrkiSccqZ/xfnmDLQHRv5I5AfDGcFYW9pr6piWLETD2Uuxj
hmIMkv6q2c+SOWExod7SPn8MLaM2yF8McGUNMR1oF6PgbXg1ndPUOvULhxOQC7V5Ngz4yoEFhNDs
4kAgRZ8sBe9REE47frHVv5Xs8nXm401uQPQJ7w3cetDKLCITM7Tb8USjkNu3SRtxbM6Qrsu5sj6U
nG98VssKA+VQS2nxEDRY3vQWPDD1hiuOl12sJ1Memhe0zy4e/LNaBTQkFwjdVPuGkzR6gyK2C0qY
tjZ9oKIm3ErzOB4GvCNGD/3Mj7xh5sE8QNu+P/v6rUisdBD5lhK67hbPL8oQBmo45TOMwlCgO6DA
9aZlEB8d7sA97VY7C+NZfut+qRkScjYkop+PVq/sl3FeLZI9B/4kT5k8ei/rliMqlR4tt2LHqI9v
YanTshGJlsUouLw6tcOpzkkmmgXRTBAEODyiwidLYsXKNZBLSGwBlFTTshNZ/rXXhhTb3vJVLIbj
bIWhebdMPmZgpSyk/4C2TUp9I1HAHu5nGlPdGSBgC4vqmrW7kzYhSIYgBshxVORGNW1jrLCeeu+B
CQKv5LpT3VxyuXJP1Rw4i0lFujqmlMcyC09k01/Q+nF8vsLXmn2sqKzktKhbbsQv1A7mXNN/Y9fm
sTXEMW22lxt/b1s8xYnXotUokHkZB9N2EQh1iIBokmyczB1jepWtIM1qjG38A9BOgMUwtfs2cybW
dcZ2tx+e4luumJz0WToA6K9BDf41wEEIr3Ba3D69z9vp+AFNbRXK5D0TJhxh1GmKlJU11Gra2Z/j
rz+Rs3lAR48KM+HBOhdBDN8p6yTViCY7JgOPfPW69x9UoaQNEW1goGt0JrxSUvosEwwJVYInx66n
rwly0J5jFIvlKsukVDxQ4vt2KNz0qsQq/MtbIkwg9Zj3n0QouhJGB3oq0/FpoNrUtgJMRyBhCSD/
oq6KCYqKkIbIRYmGPwovEJQz9gfMmulGqXyyfhHZdfK6AStmQbo0AN/owqDdbcbWAgFNM0JqUaoI
VrDhczsMdR3KR6gQPAIn3gR5L1GZroJYWUYKsGNpOStXTKhAwBMzg62uV2t62C1TK5ftXzkv86mg
ozJ9l6iOXK7TKR3toEQojcK+hih1rg/jQkZp7Ao9rmNA3EUuXdYMT5mgAX941231hjvTqiwuyHC6
iR7GXcBMZhP66IRtA2Cd41x8pniFdyH33RdAIR49GHhhtUfsGE5+lrYPtVP9lZcEgpieVSZyW2qk
rMywkhkZac3cPgzQ2WtKtG3p9OxhmCGiF0X3neaLufdElLmM2vXUMsyn+x2ajWsKm0KQIY7x1qBf
hKT6t+eBiWd4AKqeIvnYengXtiEacxLskgkuHEucmlwiAh4DT0iVPJP0MFfCQPL8D6aYykO2KEjh
7QAmbUExUXvRPZd6GLW5Q0zIm5YGEWZnMaw/2exIRfqwdiUSqdJjxcJp39V9B5ECiS0T1KnlJfjh
/VEz2g8LoJ4v9MPGwilNZWRQWMJT7Mr5oxl/955gOUeZv60y8rQB+1xrf5DSR6CXVEl98YYHJeDV
mGawcu/TZwoQGoU7Cfi6RzDB9UnOe+uj4e6XNLr+shcpB4nkzpWeP6EWPZRF0Yt2ymrDMfw3D0/g
nVj7NOyXLSCXRH3L1gBkxNPNNtQzZD2RLdJOM5bqaacGOpAGJN6AJequAB1NHv6fGuN9T9++FaBC
8Itwl/ixplLfCMnNndOx0Xb1Y4qIze5SOFnBsc5IiwaYVBjviZbHLxArzrU7bVkjeRBG9unLmOBW
5FQnXOCA/AyEVAqk8zNUzB70k6SsMX383NpFinE/Sz2YZIqgWrNhpDus88IwhG5bsrc6OVmJyC1W
loc+EjOubGGQ6lZ+KhtHWMZSuegcvGNcTozASS0vIFzO/AkfV7sTxHroDEDYW9ghRcyPYg4tK1vJ
p8fYbcD+JRaGLMCld67w/KPKiYwCgA4puJdHdMxthGjFeFEmL32cNbGnOiU3Tv8V3yyHvIGbgPDj
vPRe7eOQsImssPtS4m32x0jVFC30Bj0+FDDpfiDAmEkgb+qtU2R80sO/NUY47J7oPJOZZkLcMlJL
02d+a2LYuPdlaCf1Csvo3Dxt0t3QKwJivtOA5grF+cvp1j4467ggv4YmmVX12V3IYMhGO/wKENfM
EKC8riVObxvRx2tun9jDTHalpRzHj+qeLDWlce+KgP5kRVLPyO1eVb648gwyXlXuRaeE0CxHB4g1
Sc2QasjNyKqbkYa2I0agLJrpFKHz9uc3RAlLr6G4wFLyu8NBAQzPGGx2ThitWnmwDGyedJ3DKs0F
92C8pXfA3dXnMuU88K+/ED0HIkyDIfqwPxUjrPRwBg+0ZskeFbnhsI6mh87SyoDuCYLXQeOg45wj
unqOBhzzkHD/UFTavZuM1ATdtNdd/7isMwdSv5kCslVXOKFSK2D+CUz7V6Qs1SHeeEpAt/gmfKMr
vn5LpqMI4y5eoSfMQzLzhpxtkxa7NDpyKXANd2JBD5UXILX9V1JM3Z7wdd5zB6cicIxhBSZ5BeBS
3C2qvgNikb5BA6I2GEEjXzLLq9YtSxuWfCFPOD0kB3+VhyawD7ZQDMGxfV73hgQfVjirGwpstUCX
FQ1jZCYmXRAlw7tmICj7rJSpX3Da2pfuSbcBOv16Nvtz2ou4LenpFRGTSgoCpnronhqS/xJRKLzp
bbmItHqCwDlD85OPXB7zAUcJJ0bKbLKqicmizhrpL5ndcv4AATgO/E8kAaVEI3/FCRgyPngGmMJ6
80eoRaYkLk0ulv673Hjdw2BpMtVvl7ljslFa4LyJZ2Cgsq2kN6AKhvMcmuhMnAkJUO9a6U41LnnD
hE8LXcWcgqc3bzCb4Jd+dFYCxikydnywDvTvh88AuMD5YaizRG30RcNcW3u16awNeioi0arGEFoO
OHiul0LBYL3+JGy7+31HeZ9YMK0l2mfcefy8Z86IgmXn5Oyee3IT2YcGrBbG2+c/HdVcdNJjHLfT
CFHP9iijDBjmFv4F/qwVq8uEYYzuawaUoiuLmeD97Wc/GaPhMB1Q7xqYoMrzBDEFAD+e+kwnkzeg
ZGfLAv4lZ80PaWiG3kbS3/OHSHBCLs6RpabkWF7wapkf7uCILX1fThWpwWDl4yYcmFaVZzDI5cBg
gZyK8CMfZciH1hjmLG5qBKQLGDbqR9x/SQp4hQL1yi+E5+eXLjhGhrr0kJG7gIJatdxtBF2MBc6o
WA9pL6mgGNltBLIl3cee5KUS3ZJip4LknroxPzr4+ITKTEncIegMTnAjYnk6HCoHnCygojmDgqCG
YRolvWX6AB8sE0pWF8SKDf7NPKgwPq+Yz7oyvGIYw37S7PZMcRMb86OmVI32irE1KpHuJVd6nwF6
osconAzEb/ItjBTCK9o4nbtDp5nLJFRUjE4ZV+xLCVdrW7aqKbMCDg6Z70+IgUyepPao4b3Ple7p
yBPSb5odBwajS12NqhHHcaksVCsXk7JcfioWFuyUX4X79j4lJmxJ/i8Tw22K5cQ8Ri/x6MW6U472
a/5b1B8Ng6Fr0Q6myre3YYGB8OunfS4EuJKc9aOAkZc91u9J4mfFDN2eAHSMWtIGGm0cHhE1DUoj
Kf4nXtFDcIMWb4MLNWqFOccEyrycqL3xLpbeWSUGcE16cIS8mWbz1ebrA5sW2YbD6DQ2dHljONOF
bzrNRqaqlUoN+MZue8EATrPJHsedKbwsOI4DIwvOVXiLgcgPJXWmoyTI+0XU7CaoARbYdMeKr1/9
WlAkLp+XEyv5NsHzPOu9mzzJjFINnyl50vWOBD4q9qK+mz/7cqdLT69aNA/Z/s/GNG5P4LFfgXz4
fkrPSh2tGYNuU7cAJDP01R684iRMMCkIbeEW7xkMVHXhs8C7KCyi/IwMeHiZlyJXmuVTc3NpqALN
c0lDcqlIFhS/1JBKlM8Z5t85eedjjqoJNDqANcqm3h5RQKgRt8yt+dW/ZeaP+LzTsyJAScCvGLNk
MxywEJl/tAaJiTrIzQVo91jsETASw3mPzJ1yWozifwN8al3AVZt3T4WI7RTUJmBjPbg0oZ6rza4I
ypX6gut4VFMToQH7Hivn82EuAv7KyWhwQshZpswXSaG41TqYc82TgXZVJIEU/EN/StgXDM+G94EW
e2INvdON9Kk/AFZMIhbLR5KYd0y8qtYEQoqeRuR1K/Si1xIr2i7sh+KJj6rZto0HIGUFW3en/bPP
nnexzvY3a0k4egrTUd+D0J0nhgl52uHID4CXOPx1/oh91HCuXwCq5jIMJr1QH6h+xUXRVP5PXVbF
KWcRP3l0MDiGtljdCsJ5SAstEdCkjEtgxq3vsPPvg8O2lpDKepF1qIPciXXuLcXXQTTaoVwqhapK
iHUYu5ZiX2sO/QzKq+w3VQGhfP6ejfPs3QG7MnqkEaGkK5PdKy0huA9vspv/QIJg4e+ysNgfdeEV
oDfmeIfybjkga5JUaDF7MA0YEvCurIAQyk8Xrrr/oeXPOuAJ2WxAkoH2qFuk2vDb2ti+Pi9GmH9l
KZJq8wPyT+wWlRqDkDRh5KsD5I4pwTBHm/FhXUPtW4sR13j+4cxBdqlHr3WVWCMxew51hrvS4DSg
Upd3vCs0I9GJUOLZS/kan8gj/g3FmpFf9RCijw+dIJru5PbfaiRgUVQinOiGV3hEBcPUjj7WIOkW
xV+IUbVwJMIi6gHjS3LmT6/G2g8Cg6N2wMZnJD9sOdo47FqK/FUF04jSj89na6Ctm/plmu0VkfH4
SPA9vYn7grDEzuiR2KAWImkgpU2EeC11nri6VcpqCQACvx1o+KTH5IFINJmycLD6tquTmy+jZVoo
XA8G1kniLfMshFsyji2MnJs88tKo8gfen82YeTQk1JkaMygY8CRUs4YK+/fBmoOwxv7tTnnSrj0z
7dtOblw4utksnb014uOHUZppLPq8wvo6jLhL+1VzYExgoWPhqjeYc+manooIIvSY+XZceiiokz5p
Rv6/PMvFvLJZgOhHx/T+NGZFQCzm8AxHQZZXFV9bRLybJfuUg6o2qOFqm8XMVQz4MdRx1AODLdkC
Rg0w5aRmxkGqp1vYRPcVfrfIe/HhwP9mz/+s/NWjoCBVBRkU5hT1UWdzrPbUmC8M9DSqVhFmANF2
a2CAvyPtH2rIsQTmpk5uvpGNB2HsnGNKZ8FPnh+fSZIo/LxTbAM+lC3UOUAJ+CicMFYbaLCPRsxd
QPOzeLSrg7WHdtbp06M2bzbikqMt4UWdIuvYthfxMishSaNaX+X9tu1SqYpoQJFlb3JwU/Cq2Li5
DT0Drr1UC1mduYaQ5T+uTitjME0VF8xtIFjqyXYpNub6GmFd15cM8/PyfFdfD+oSfULUCOlfAEz+
CDZeDG2BWstt2HSP+mgo0ThhljidPnZ5vwqx7cygGTiRH2Qw55cUhx4joaoYh1B5Q6fiZe35ikdd
emGBBcY0RkA0/1U5S9JtTwWqw/hoL0TbSqnuDuCKY/ZDvsvGY/v39PVJvgrsc7U6jNEF1AaP5CZM
Wna4P9ysywMxXy2pdZb+9pkeDsUlqm/vkisLUWljfbn41loQDbJJaN+R/KjVSyzOtsCEh5SmMy2+
ju8op7giy7/iC/EUgmeWVYkrUJt4/Rg+D80tp9kxuirEkhOQYqRouK3aQsOPBeKBdrk3fJcVTBwG
wEmmsaeTBe0CD0zmiOO9j5cnTh70xEZTeBP9Iz+U9LZNxGj6ewBIWv6afoSAaIaPLJ0cbe68t1C1
lPH4fhJN5aUB3QXZlfIJvyEyyC4yylhBDUkywSly2kOeiWaRFtZz4eIIOVIJmMuTrwadh+EMfuqs
bXqDeM0MeKgo53X/crq9NFMdI09Q+CkdvN8cNhFLz+9otK0nwdCBNeJNc5BjoUqurwpdYvQmTI2T
pWgnSkWksxHO4ZlW8bM6nDEbgEvTSfGFKWUhSVjS6WlTgBMp4Xi9O/r9RD4PbFiv1ehXqpNUE4Pb
Mh/mhLlBn0d6cQyNmxX+XcXi+ZOePf2TXgNMkU6OKWADbcqCkDAox6pk15Mbfhg3c3UPfJleYkLz
dUJAl2T3crJ0utUh18+xnI7WK/eaXmre9vMzFmDohz2106AB/2zFRWy2pXQLuBHqQQ9qTEtEwJkf
YJ/szDRvbsoH0FlrEIR7wwt+cFha/w9Ya2Vdt0UDyfvbWhnIE3WkwycLB+xCOsCBey/DMN3CozD1
/WjZNil731nHoNgrMmjrh5pCBAa9J3ouPKSP9hxqV8w74E4soH3IFK6ZxJCeKUBJoUoUIt7mq+Kp
lXU+bXBXanaAljoVArwTb9KgU9JKRN4NrB5fHo0D0eAlgUsFUowiy0hiSt257OwP2hevMWsW/OZ1
NvfHnHbPftH00Re9XZKxmwDvf4Lw4ZgD8TOq9CNQjn3JbKijpwk+w3pNDeVGb3d5nk4X4v4W5yuO
0cGCNKkhcI8L6DCargPT2WnTvknMaU+OC43hyqEeQ88kLyEcZoYcRA5RmS/8xygufppeDj0FiB05
z0eLNLmWultgg8f+VDww5BiiYxagSP9hOmmyz/5XsI7Enf5yVMUZ+fE28bP6F6L7Wrt8kUv9+hOO
ZorWrpGcynSMTmcHJsll+1wuggzzibynuaUJKfxBzYAr8+4yly1cI916FShXTMVS7okFVeCJ8TWo
LpU+xS7tezSJyxDCVTiWv/48laiJwZ3utyyh2vkeVLxKPJjd43vj65+F2km9hxlnrUk9fq9I3jBR
l/ofnDZHaAfiojK0UKOeeZscy3HMZxnbLBrBjF0ObaemeL1MC2T9n1d637DFzFQb1zTrNHUqdC/u
ki1vjg3Jqlnnvfb8D58qI6ZFdERWTmS6NTw+zhStu/OCRAVACF3QpPpUWhAWu3abQ+TJ7iwEMtQU
2DijgGWto2SkOgswpTjWoy0pANtkKEz2jzEjqBc2Xz8f1OEcMLi7ZP52YJuTDhOzna8Y6lup1A9m
LVzPHbPZ3H4UTZb6EQYk7+lGt1C1Ps7bGbkDGLC6YUj+3ZFZ5eGYgYF+qhSrvWKP/XkuePthpLXs
yj/7oEGK4fwiMljeWKhSDK5I+6IWMTcTCVm9sjFdJN37JY9wIPB5E+4NPZ8JorvZdc5R5HLfSVlN
RWwXz3hhNSXjubcE6q84iCN8krW6T7QQzITlhOCQPuBzEFHamhH8Y2EzJOIccWZ38v/VfhrmPvok
E6bv/7+GaXjExedbdTByu9nS6ZRuJqWq1nnQth8RuwR3taT9+W6CPHQBhcYfR2pLNXvjt6UJg2Ik
wQf/66USqK6JXSOS6LQLglRGDzlGNS3G92XxIbTaX+c1h79n2EKORQw1nLzSgz7XavkwmCTYhtj7
hs36D0HTkf7zMcmvWTTynlXwyuoqzgqtg3/sUKoqdZEcqByVDwMrrvxPpK/OsRDR+3YoNRdpucZ6
gi8lyHAlcIa+4KzP09aIHRQ+yVu1W8m+6Xm1rtJ+xgARSuLAM6e/70DyegydKCj9nnlo4rxaJsZd
1Fqx1YYubXTs4w7/+QFfRQm3p9nujBwn4dEJyU+6W2l0SjIvBo+jPcSuPj/aGSvhjTCuuDMyC49f
RpwdpDtyYx5Vzx1qoJXB5e9B7AIzyqKsVblSZP77bpyc0mL9coK2Ab3iJ+278sui3xbLuHNUKe5M
EurcGY5yp1bXuY1B4sFKzRYVtCGH1GZ4YYFusREoFpJgH6Sa96RPESMvX6Z82RreW2YeGY1Rx2kN
T8e4z4QX22bPBXfMduCp1191TwDdOxslZiFCbuWLfPcLcGcaz4qyDzOHoyK6JQVXyQcZAcrHcfEs
XJxADAhV4ZeUrroTkPdquPSTouIfd/n61FlQGHbZi1iNKucIZ3hykcrV/f6D4+jgMoaUUid/Xe79
E91Qn3Wpu+axCQvLyEJH4n8IECFruK6tKbIuv9podlTcjIe7ds8fuEua1QJ3162K2HcPmdDVQP2X
4EjOGAuVcX6N2XGngPUbDc491hIhNDpNjabMw/994jJatUymbO8wBYu6E8hYSQ0GiXgJI1e0wYZ8
2B1AzQ/KvvMIjdR/Y4tpLEPEII4gkC5kPgsgd+xPOySo4VXo+RRsk85HiQmTGciK3MSd4vLx50tK
QSi4ZEBAoqEqKGCEkTQvHwVt4E5ey/elZUVzgVFWurGjVytaPVNmctW2LUHaTFuMCgLAf7f31AUE
KxdBKLLP9qlQLFnV7RPFu49vxCdSUQlkkMm414FcxEoi/cZB3HQq2dZ+VgUfF3qdwlSZU2hYokdS
t0D52F6Sc4Ezzuh0I27xT92PpIWkthqP/4t1a85ek84MnEXIRTDPPl3G5BqXO9Qd7utdIXDHSeTq
SxXp4OcuFywb7qOh/7KIoGlnwTpsBYyO/JZOqpdBWaAGwcDxCLxZoT5VjFR0doN4uIyoQOwfB/B+
iD5cwZ9g2FdCJV/IIYgfimtZmJ94ZmEsXXvAB4/mFNZXbAYec3D938taV6smNG4TasgF0qS2tpSH
HuKBNRNbdnXkZ4IZEdwfgZk2ozKG9pIH1VJFhsEESr+bxGdTB5e4Wwf59jCtSDx2ckxbIFO1ysRE
8XIsD8jHmO6d1a3RmQMBf14TmTdma05XLPEMuPIHfMFJAONdbivbJA3fhRlUBNmTcGR/8JZ25oLz
CtMzYgLXhJJZWZi/n1Ex6CNITHgmRm+rHrFO7d1ubGmGRbzW8YjhrY6qk3CT6Fff8SGl5c0ERBzj
p8b0vU6/BdZadOKnXD0EWNirx/xLDRg2tor8/FiCYQ0d+PgwQU29XkNxL7AyNTTlAwKIY4lPasbx
/4U0a8lDfvtGaTzZfcHP7lKVpmNeZLX1Tj1lWEH0e7NaD1OS3N6ZofGwwGfFEB9omhL/qooddgEK
AEiMBBVbExaJTKSuxZb7TPpdTWQu0tSYdQLzdY2Goci+/sKUwgTXIy9/F1aJ4l/HQEShL3n5Ksxc
SkTenqcZiHVfAMCHPVi1qoMHCbFfvWrSUP0O/tllAcqciZxAuTavWmQlZUpGCoEdfIJlxVxq13gL
Krjr0IZp5Otmfxei7kpV/wXYWs++EQWts/qSlWcGcL00RoLx2anw+ZVgyoK31E1n7eJoF1GbiMgG
CBaPwAGXQNb/zBrpsDuOUr1Xm3FJF8/UMcKG1VKdyMpJdKxdjcgniMhFkk+eUJKr9geGzfKkO/Ap
6KJKQ3Q6RNHbc4cq3QyQ3Go6fjNCiPyE0SG9apSLv0KVNBBjp7+9XolNN+PjaSG1c3iUjowoxwFW
oktQQ+ylGYEoLoJQdaPaH2g0KTLjDy3L8IyDBgqOJYUSjFc4pzChpVTDx5w7zzOhG5ugV+6ibnru
lg0b4GZ5AssU6VnqaHZUqS90MbTsQkCZfabL0CisO654zOiUwSuSFnzj0mNRK2EACMqihjf4xA5w
9uElrIDQLLZyriPrwF/Lfv7f4NDUqpsKfNG0kXRUWq9HLZQVo8Vfhq04bRHDRrHETWcQjh2g40Pt
RmOIkMTLaa+nRZki1afNwQRzs7otCWNtZ05eWmDhBuLacGDbpwX3mW16GMnChi1lzXqpX/c3vQga
bB7YRXIvlLDjO5mFuCZLj0bkOvYZFR8T0oRc5xjFvXJp6uidsKIrH9nVkTvxd5v3uB9oBvposLm6
rztwLQygZ6UKP831FXmzvgWQAuWK7PALFdQ9UFC1czrUD1sl4jBgoD2WpTZ6veQ+UnIaGqX5AU+F
rox0Ug00nPJgAsSDl7NgCBfDWxDafUctMmhRY6kU4pGsvy18T/yDC0wfiqeI1N2PbaVWIaBtcgS+
nuu7hJJPUKtGXS3AGW8WUi8L1sahy3dzWuL9iZ4ASzCB+gF475/UWxoXegE7Ml/IKNX0O7HK19ZE
+RCb+ezIgu8nuH3SeO+GFQCXEIcyx4Rx4M+c51h1mUUTjhLdtNacNKrvg1+k3K9RFIXfTvriFULH
xKcoyuV/Fpy2R1WcRFs9SxMIbC7MCrXRe5T2+cev0ykniCBqYJtPxqtBl1yi+gRR64LAYQFTLzi6
RNKa8Bz2e10nhH67NI1y5SpxgTe7XJofpl1rfVdJPiWi4VRRLNHrsA9hAOXBWx30n5CtpD2r8oTD
0K2pM41wYuiWVCI5g+2exRK09gQ/klb9r46TDGvnVOcDl1A7qnobUn1WEDTl+nwLk95GFV4RRl/u
/aPul5ztVbOWHlzp2wklPQ268upe0e7VEX8pasvZICMzakM5TVuocakCXcG+ihXMTHYPAnOPsxu2
Ba7BZJfs4H5sf2PHqquaeEOeY71Olzus09Id74FgSlROY7x+YauKMsQHc1hIwjn1Xt0Q1oqhhBD5
YGGzAimqlP5MqDU3KIN5aprwtiehZSJwxqqe5rjPpfTx23QXewvPnviVMID+H/CRvhdOANgqFQer
+Iwzd3gv/aHZylIT2d1xPY2B/KbdDggQJsykFbZ6vxUW4qDqSFU5perLbUqoaFIiuXpwR/jwDuF2
8ZwLxKS0VHzw6p/voQZtPM6RsBNEiODOZ3SLuP9Wlp9rF3VrGZ+tPGHBn95xlmsL7U/SS/cFdDsZ
vfPDnhAZdiDpL8mWiadxO4FrQqamVkXYp6pXmCmjRlEJ0rCYkM13PVTqPjPX4MPfkz6mCUOLIdtN
klYjDlGe582nHGnWWYK2+Rx1mMAJ6NUwKsnKGUgnFOJP09/ttaPH9Re9D0f9mxdPsAhdeE2Rk4xy
W6k5kwGRRfIeQ3U0fI3L0KYoQLwE6WVfdsnEaCxKG1mPoldgOajNaV7TllxEvLOLQphUW5RFd0AD
h015MgRsHQDs5FXYv5BKTPV7A92urQOmFgV3zg+dOagzYLOwGfA63J33OJ3K5jUADxAkJRc4iCkG
VrGMSkSh0tfCo4IZC+pdHy/PyPOTOVUi8WSLd51C6GoW253YE5FcODsr7QzrYFtvgrbfpGVDgtQS
nWPQzzBpWGs1V68+xDNMOnlRi+VDkmicIVRwKNzvAmKvw8PsTudVEm/f6YTNhHgxRvw404leoWqu
7wpQDNUuY1iejipcvMb+vf65DWBaz41zTLelo29eIA6Afivsri5unHmq/xrKVfKS4fhOT0lAezcC
LxUZoIMRQIYIhBYjRFcWtc0qTNoUGT9elYMbl7tthuyZTnMwAq9ijpkp9qLAlY2eap6lXJZLSIkz
H0EU23aDvFtUkZeaONaVEFEMR4UdE3vJrlmfXn7fEjOhc18Sdq4dX5KsN7ZPC/UK5U568hlx/z6W
Ea1ORrvq0rpG2yN9SCkxPBkBm0GGtude5g+cwY038bf3pTMeeVjAQ2HoW9VjQgF0j3eCLoPEBunN
+bdGaWwirVlN2i0lsFtH9XPfS9kQyFnvlCMr3WSUv9TCqL9Pt792wB181vBBhuu9ZoCGWdeGpLYt
w208jHgeyKyFvrlLmOXhxDiUcwN/OMU+oKcl08FeUYnEYXUM4iiykUyUyn5f3pHdBHj8lZYL2Aaz
n6ASDL2J+6cHhpNiP54Upn1sPeMKrx9Hvpq6XmjokRjCcyVQzMcwZloOi103PynxF6O36iqSB9bJ
E/BOkWWoNt4LnU9l1llpbR+GlLdZC6Ck2JP0rFDKQB1U7PHcI1i6QViNjLu41AN2j7tYcYyYI76W
5RZFvH4KTBaHgycf3LLGNBPGJLRwYaKIv6gu+zCObKD0A7dn0Jc+Jr0qDsJBLEaEqVU7aUDW/5Ff
fiThynfvrrYDcgIHJyu0L9yaPnoO21YjpV1pb9/efmxevzFkmG0cvGr23v+mBvUYGJZIOCJcEcTJ
crwWC6s/Z2pcnkmnq+8x7FQcWic36Bz32bkZyO8qFTBgX+XoyrCuqP0kl7bo0XoYguOKEQUwMGxy
QhxIrKHHUVkRaBnB6LCrM6Qc6FVJnZQ/jdCAUJqMmrrxwIJWyhSp3o4EYhbSWzFNGZ1OkGMQ75jM
0eYYObBD9jGwxIuIE3o1HAXDbLVrP58BG2U4SXgRZptIBt08WdEH3g7HU9fmKp+p1MAkaSKYUwTf
jlvWp7DhTSpl0cpnq1YWRxzxqMLHVLsZETgDHBYkZpTJMG75Jg9VuEl20R+UgUXlb8NIC/zWET1D
HSxxzbE3bAW/ZGemKOFV2MxBoDk12pRcjY1a6hgtXRgURR43LaL39Y7o0Ir2EshxKmOjrApf1l9H
WZ3+mgjm4Zt6Jw0jlY7VZ8Ep1+mnvwRf3FkkP1I36vpTD0F+arx9MMWkylv3+zXUc1B2MlZcEBeG
JpreoYIbT0/DgrDlnRl8lpB4sqDwp1GVz9pbN7+cBwfhxRB5axA1io6dUzBYiCRYqOSeYBlyeVDG
XdoUjP4EewxQyOKljrCejPvfad7fzn4QrTrg/+0ZX9XeKgU1AhxZGSaubd3HRviicAqDteGGWN97
l94j1nJn26Rb/wxqmAe8ZipilJDWq12bdjmRhwPIu8SMpE6v0qILrmEMRhRgIHjxQ8acGyfzj2/N
G4ZQks44XxnMqL6YJU6Z73gXdmv74nacqQjZnqyWnBIu2CtYpd42qPVBgybzxdkYHAeTdg5BN83O
M5yQeHjA+zTnV0Pyqd4ko5BoW82Vcm2t3rkxEhnz/z5kx+eTYvfjzw4h03hWZINcPfgq0Dj+3cOU
MvDF3pAF/CdJ4F1j4sem4ERa5x93EuhsSuoc1YLSd2HlMWJfKUF3H1+ftaAJT5ZjD3QJKZLNuyQq
NWvNZV2f5BJ+Ex0KNiCyhFddbYWAatm+BnssE5RSJ+gl6wJVql44EDBENObY0vvhIHGlIdJx1a1+
JKrFHvFnrKXkMg2c63J5NuNVb9wZ86+QnzKnw9L285wd8GguGbeLykw2YvRnr3nVkzzlR1XGSwTv
4Wum5EusWH3S+0LL5wcJHdap1AwQWYRWUqwv8aqSxDEReIn6C+k7IbN4PY1wdSsWe/ObNykXv5Ak
zDRSy8OYk7zyvT/c24EH6lJSL+gUfmJopYo1NrOTUVV3eeDIG0Wix/vfB481gdPlBEX6eofK9+IG
gHyCZHrejrrYaKcG441jHce67IL38EuR/XT5uWBn2RvtkV9Cn6Ri3bp+lOifdWsluKlOK5GCKE1a
czR66E4TdmNG4e4HhrmnqqL264i9A8b+mqi299gimClw5RGr44PPixAug7fxBO22YYIpICVC4vHi
E6wm1KSJP3t1TW2KfhIJQLQzg0T3yyulsqd7EQqfVI61s7VlZZ+NaM4Tv8G4L/xGEiqmeFR+ZIq6
9ljkjFBXzLqBFZ0DLIYWj7bA95attJ4B9uofpzRvrdSCE0rbGnYl6z3q+yZIXJodd7pgtVrAFvst
kjgrGPbRoBFb/Oeu8nlBOy9nIPjeZXuqlgwIlc3Y3kKAV/+0nls9PjDGfzGKeBdu5dh2FdbD7brQ
vC4dn76puHVQyQc096SJnh4rRpRbp96mDIxxhK5RP2Oz4k6cZf/HbRcDOTGczwiyV2n9nOgo2RCp
pHsj1F6m9UH4/K1aDR2yygfoh3+PKKH7bZsU9Tc1eT2mi4mdad+kKNi5wrAqWPQKZarD0yn4wR7l
7tAdxiYr0TDDEpo4dZn1jeBhB+4imQVAikZNmBu6knYtFekKtqFv3Owf14pIqvoOTua/qj6sItz+
DYpyXcSu0eRYvhm6YpDgTUqQn6SDR6EdujQAGXCd5ovpGHvdjd0pfs0mpjHc2/NakJEzBVAsrFJy
doY0/P8IpqjAhxEi5uaof9HuNGpPqM0PpE1D10yYvJkQxKuR83XEfaRG0OJrIOmnLvtQV5/ENbzr
S8QmT5LXSCKEFFKSC+DfF5UBJDFcszA/9mzh5zgAhS8RNtIqEBN/QoU2KhhIUvnQhhs6PzLjq/nx
6FIYBI0+w/MFYRAUy6shYYkiT8LSJl0tcDL6JBmZB6nOuNRcl4adBSJJLCU4Hpp7AE3SxclEi4Et
oSC0D13XV9zl1TO/2TIeBDmWmj5Up/XaRKfiSQhilL2oMjQzyi/1DzBsgOH0uEWlCjZV3ruerwDK
+ShLUnUnig2SzNxA8k1gy/a2xfhkJs9tvxDEYl0ZbJh9x1Fmi2l9eDYQ1oTWAfNQE0S1k+DbEekV
/jehKyD1aoJ9lQyHeg1AXeR2vyxftlcr0G/QoJ5P2nsUWvWR0Civ/wW8VbtGlywdX2U8Ak6KP5v4
AwBvU4jZVEQplW5AXIIp7XKy5z93fqduijT0JvXco/IPP4ywRVjDiEWxaP1ofSJW/LEurPMmg7tg
Y9laVUI8pEml96mlsYK+ai9xz6TtzMYetR57f6I8QRMphZFLPk7OPFyPI99gbtCzH9v4snzicOUj
o65MAe5rbJKKp+dZlCxHaIzD61bMYkB1sHitp+eodvrZRBjwbmg6gchT20EYhn67POuhGTZRfkKn
EUD7hf+J4HkWVOqsvobY6aBhouODDXngXxNPy+YASzA0YlTK7fd0MPp148QQ4DQn3tHPsMBARdo8
2OuvG1eiU1pxHA1+ataxft/9kINjRE75o01Vm1ltYOuwb++gbfiH5sMgphFC0NetPC6q8ya+zMEH
kqyUJ+Ik7rQcvrRGvFbQTt9vwo1q+E6Ncpiv51zVBwEjZ0y1olIPbsaYejVvn+Q6oJDxzsLGuroe
q2MX/FzLpZBHwdNLmc4j1MX50VGHUAUWVvsCqoQnu4MlY4Ak2V3TiwRgfTY31Lr9RSmwfUYi2+bC
UbrStS8FLkO1MO69M5PT5rGZCFNq6ouq6uWxcDxgoIXW4Gy7bCSuuEMAmgOLEkxs3S70zGvF1cXJ
0jb0y67JO1P2bLUed8tXq5qS6ewyl9gSulf3t3F53PwpHT1BYLNtyXytHi3NpmleVZOoYoq2L8Tm
eUfmTwMKuq8zVI7rMacWedAZGMLfLGtXcell3zbUAY8IyNJGIHpHareARus90IkicaXAlNtggOIz
mLKxoyvPgfSY3MysaSg4sNr1hnguDPcho65C0394IXvzIvA9KvchxKfsh4tlSqcZJKWjMeJoIpGT
dypjp5lRI9O0LITSLQ0a/BILJ5ym5bkQ/SAL3gfnzUAoB/rKdCIpOiufJkVhVatKT4kAHV9AE2/9
bZN7+pwhaeW8zH+Qnusa2/JYTQ+gVtKxuAo4diaMs2lyxF7opTYrPuMFH6YUSYYMzv72MQ7QhXfw
61+buAY7shcdDRzOB+dx/j8jxUiOnCph+P1sQWUqOJB19IXbQdStOqFtpXtzLuPnOC+ROoA2jisq
RQR5aYHHfS27MiqEeAlwBTSI8xP52ZHQ1MP/KL9x2TLYOQrfKsjfCMhC4BNe/8x1RpLUwoQb+1+x
aB8d21pWjWCP4ItT/uMG3xJ2N/wmt7BIw/HIDPhMwdI+3BI9Y7ap8KIhc2T6F3/gzMKNFl5M68sn
2SEUNVt0idPeiPJ+b6fHIebjxe0fau5XF90wdnQOYgyqIzjDohS17w9AH4oWrjMJG3t4UNMMTUu/
YbQjaSPGnERAIvwX4XVpbFR6iFYTeHd0Y/JxGTcfm89IHHww0w47x4Q2aw7jwYwNVfSyXm5BVIKH
mlP1x79o7Ch723dzwIVcrE2FD5khZopWryOBvbBtwuFe2d+AmyBygA46vYJrVjJj2dFBW19VJHiL
9NiRdGOpSVtR4dV2kHAtnT84nfeMkw9mYtoVUJXgDWb/NlDOuwcFXuhjvnustDHBUx3qw+PQBRZX
pUTMYsF6awNZlCJk2lZKET5tl+SVaAwDHU6vZUyrxB0or6eZBoV/n+E3Pj0aO68MfzD9OwQQWK98
7OXF6IfnmnaGLDz96bcIvoXFCbLXli882cv0XekJ7636BUoBfUaibw4d8NPM6FIxBiinxMyIZkNX
WZurERY7dwK9sKSW3NqgAxLBBsMd19vt9ESSOxNFkEjkSSyxMOCSZmnlPKLSH4jiPC3f9Pfj+kuR
vLjmgjzXjyZwk77GtO6bzmRMAotrYVSa1rS+voGHcYgq1r+xWzZSd46B79XQMqCbmxxp5WIetN+D
prcgjmJCteqNkhkSGB3dCzqzb3iWccQHL/1nWIuFGvMSOzTnRWlHUTXLg7TTQBUQ09xtGRJnnqUP
sR74csd4LC+aXK3doT35CJvNFXHlcmVXL6O7aSjsJ0HS6G8Rp5OKj0ZQVim1YnCFTwH0pr+on5Ba
Vt+F5U4fOhT+0FmoelKwIFxcEdSINFSdoWJIpQSOsDayTPiG4DL055aDmGZtBIzo/06Eqb8oSSpT
hQmBFtYZZQesN3MQddZYtfd038KmuR3wgsIS+gN2or0OOKpdCwHTgG6Oi/mRIAOdcXSPk4jeQzwP
SjqUbs5OEreg2TAGP0dPnw/TCIN29QB8hFAa65VcjIwhV6yVubV8LyOcKwK8soVnNEBRO++3zsLO
pHfpaEstExrYdf36tvs14VpLO2y8HdtmyuXFVUCUbqkvW0Q4bJFckDL45KhioICnX3ZGPQYE7Mt0
QTKMfys+fUuQz/DdOQrulMIo1icEs/G3zfN5COYzUt1Qy0po67w3ybfQnwDrPXVB9WijGzVCVXYy
u09Bc9QzRVYiMYSwb8UkB3UgIFnI13jfSZo4U6PfZguVWb7LdxG6UiKyxI9SpATde62sLHuMJhpr
kj0AOHEzP1/xxpJpfBlRm+z0H+B7fv+YVFmsZ3qk4u/M1Dn8ymSshwYK/e7mIfhxoUw0W9QVq2sb
8n+1sDXElYEimxCUc5MGVkBe2stThH+t47vxC6HtBXsPAp2GRmOSFBSVQk8qzUgDvLjL795VFcY4
V2qqu9VZJTpkCe+OvWcaZOF6uBjMGAKQN+l4DDaIDUD1tvzggSUn/icJuo9eSibiusnAhG2j+ZKz
QOEXodARFl1fldJ9uKmKuyDRc+f08med1P0If2ZqOplMmwd6KzO4jBHqRBR+2CDBxy7F8QvaLQXN
xE7OQ602VkRSY3M9lqpi971RmUx81hHWoP1t74p6nsPiqgBN7N4m5JbCXPM9s4hXsit2DUdI4brX
w1ERkh4ebuZaVnz2FSi/ytoiUaOVsX/z70e8SVuEoIQzMzvErZGXNO/jLCUslKDgAxuEnd4goGaH
s2Azg5+6Uyvvqt0duf5dYN5qrE4//3WtnATFJg0n7lcgTYbwPqBhKL66D3um7G/O35uYbAGurXhS
/JhtyfhN0eUacPs72o+1IEzVXY9ET1wDuYxhGT6YPNHhbNkVLBsyFv5EhlDBb/+oJ3GDKL0gZHwA
q0fyKrCO0WwLsaSW0rCTbCrxvc2ZcOGdOdcJmVntq1Qw7tX6SX7xIni/zsuDemogGnjMAq5zkGNG
tSLwh52EdeH0OjkaWKuqO13jyUsCXTl6njw32XjMPmPVBLtSH8fafw5D2t0FYxb+Js893L24CayA
2HQ6DO3Y6Q36P81yltD7F1H6i7yZzrs5UW7/zUGgLraS/Soy3b4D1ooWgKPCqkT1qhgJfUyVvxTA
kSeG1J7ACNAtqw2od3CvUyFFyK1MM+DDU9zSZ9GlXDAecY3tg9PeU0Wnnf8J+97H4Wg8wakse1nx
Nvimm732eLAr2Du3mSpy7cL3EapoyoqHZhzuqaCtvhIdYyzs7dCP4htN1t/6mhgnkM4767kRPadp
8Am439O5arO6bAN3lEpCF87EFjX4p3PpD2QjCwkvoyfCylzExiGrS3bjkxhoJhRo+QkAdBvOjZRv
IfsGCaEGg1YM7tQU8JpSzWXt2ODFUjTAcII0HncSzbtwnYJOTNHMUYvgygxk4NTAZOntOZ7/LkUH
kqfh7QCKP8tsrgHtq+C552s6YQj0Qkm3kLHn4fXpym6xSl2drprQpTc+MY8bkpfUHVrfQWWUVXDk
WjNTpio91rZrqFeCq2A0xnK/QLAAdhysoFgoJMFIZzgBGu93jgvF1bn5GRoirb1aKt57vtndaVTI
/0lFWd4nZIp4q7npIKtFlT3R+Gt8mmFKCqVIVMLgLNgaHSUSC13C9fBRpadS2cmd3UT8yWsbuy4o
6R/CK4j6dZplyc7Ae8yCaD6sbsafREw/oavuyELh7fpWeGBnoc6YJozPQeC8l7leWivCZmJBHHss
NRAkrQyX9OaWT7fE4o4A2Djtq67pTh2gaM8TIcrPpPWDu9Gs4Uua/jkzdj7GOP/dsUIOWDOdayYF
En8a4n990QQX9Oj78DYp7g/qEz1ahnU6nqGliWE5guO6dzfy7GqzWW4o7jCBsICD6OB3hDdw6KB6
BC4HUkX1aFXa/Gk1oQWp2PXZyA5HUUctOnKS6XyzckQVDn0+Whg2b4rzw7r8GxjTC0fev94wN1Ey
EL68e8/jcejRqywIL055j2eGvLVmKcZcnRtokGi+TA21lZzjGV+ISG4QCBF1VnsbzI22UxoNRqcA
bWN6NSMbMITNYK0ua/COoLQ6Vi6RgwKXUjyTeFVetQjT/u58S5nvGw4+6LHi0q7e+n3FGdqh7hON
/oWUK2WzobZE6xBLZUXopuIszcq2bKvN62qqfvuT/xU1DGQV4Ird1RiqSJl6JFlnzok/5luQuzpl
PFa+1w6fUAVzvlmHhRDYCK6U9JVjn0CfzJweDyVTzmjm5y5njqQZtfkqjjpevMfWazrdNtJxXDeW
EjHIYfuF5nfOFUJGSoIHidpoLorjpbXCPR8VVfLzWy+b0xPsy2wrePvQKjRFitXKbOOV1lDJWrQJ
WpSIrcIbCUGePp4rWRnjZYMXVdrlSYbx5x2C56+Sc4Lo6UELCaCdUE5UtexfRin8miTTM18yYlXF
Bg0tND0DopPmX302elpFRsp6cRsREGBfs61BaMkAAZfemoShg5WsUIPOvfASTkdsBMTxNYR/1Jwt
DieuU/pzGwgeXknxoo9Q44cIH4bh2tJLUDx3QuWCliDYMHJ2jxu7yJorIbI9uL7qfxUiRNd6hirw
20UvX/X55GJCg4eXPr5XuptuP88SaO8nE10tQ98A6N+q2NLjKljnoEn5KLkFcWrcaLGq3t2x2/aP
AbKwIYkLnXrNB5eKb6jFyqAY7rlep7AhlwqkzIqo14ya2Ruqqb3A9ZXMlyd/o/KKc61JIJ9waxQS
x5dKx6pcthMOxvHHvJR65LwzJQsNDYOpCXKkSVvWxKOYl8THSAmoF0QWrDdCqloLSSjAEcoFwUIy
bV03GoWU6HcNbMhrhvSzS4dpV5XSC17fCUwY45y1qDlv8wyTr4dkPjDYBMT0zbO+8qdhcjZCY7zD
Niq6l6yi7Y/kEGvOGr61nM7d7uwaUHdY7a1P6ktQBI9c4NbUXGNUY/9P7/MlYfkMf4vskmavDPm/
qYWTmq0TGRuHxaaKZ7k0Pkgb2zjii3LOXh/O4IL3cRdQEg8S65FAWN4BzCVGYtJioWbIuCloENPV
iHFaZiZwHqmt1bIiU8HkbQ64UTNcrADykP8gSPFwjecHGPdDET0TLZf7gQNblgxIyRLL+r6jBDvw
9DcULBmZM00u0DPeNk71pJD6uKvkcxWlJhNybumwKgGbX+UJ21Vn0R+hVvIpWWZ+rBEjfhj8ZFy/
eMSyXQ4+EP3MjI/kFbJ75BxLH774TD6uLzyPt0P5tLioo2QCiIjp6iu5q9WRb85HlqJhVbMU6+0h
Tawm4mnBd7tLTPZOUVZwJcLtCvTubr7zxyHYoj4xnP0vbGs+kJyKvAPL578dwV6Wo912Gg7rcaKf
LIuuxVvlMCd2+6jCylj2f6d0uSa1OB4S9F14xicyUCRdkq92oTnPgqRUNTpqtF4XZR+89sFHbTwz
SQ0r1Yw8LS5Qp2xOmMkb0PD5d+OxQJPg/QVaQ8JdvljRaw80oXOJiLqnSCooaFgb0upFmgC2vpAo
nICQa4YDyaYfz754cYO+7uv+YHkaEwD19dXXCBs2VMH9Mj2fwYjVGiD/K+V9Bu/XpFcoyCD/B6PX
7UybcpGi3vKEFOEYuJCPXFf3RHWs051rsyrxgWT5rAKDDM03z/ROZCPBzq7cv+tMN6JABpFp0slt
LdqMz4FVwDNopSLvZteyqVofQuLJksjMIX5YqrpfKgiavKW52KxRBQaOQ49VDRtbUo9hGzwE8jGc
ST702ABFCVVfN14of0rgjHXm1HntZry7xZLfG5q7wVzB/hi/5WNcdodOfLccLd5yOF9eTKvkZGIp
5fKUnyYlRgYDL9//JUukGjOCSU76HyOaZPTBXJCEvOkwf1/8rXvxslTGzI3QQgXO1P0le1n0+tHG
vD/fB457KjWcvj2T7gF9RMiyExC1RuSzu96p7vTI8hWRnp4aKJxajxZ8C6SwFbUpfvSh+RQwDxfq
ueiFMc2orRsMZhMZqsKWnw41osQ7sayZXPJMUW6gfRk87hhxv/ZeT8XjEUexS0KmqU/HMZwO7Bi3
pE5jUonrVmeC28FRIl9XBDf6tAYK2Y9HHpjJNzPYzsB/I2PlzGdyWHEVR9gZn5ZJyxh6+NshaiF7
DMYPGZ6vQsNTKJNSvxSG11FD7gweqGiZqeLy3WZSM/TrdA+1HZIAl6tHV7tNy6tBqyHnFN8zOwmh
dearWx015+ifby/Iy8b9Ri8SBcfgK5jP+YBYJr5lKgiAolUbgXCeYsE7YF/+ouXdx8NFraSpKKl9
KfenInOPR0+EPySaxaYQMRssdw77y7fCgCCjABMN5J30LbaeUAf4xCawwrTE6d5EaOW6r9jBTkyl
5JKt4I2lzHbvI4lBpwVqKXMzrGtq2VYRtKsuW+gaxv5AgEMN4FYI9n4/g1yiu+wOYhy72WEhwZ0o
bBaibVW7WUQPcbXfSC1qm+wHNH0v1c8l3aU7ERL4DefPn++Eo5PfkvUKzxjfwHeNySfipkfaHlrJ
P4Qwbpmg0dmQb4g1WTBj1gBVr2DyiFV3us4jikjsQyuVpKfKPv77YdXhH52fkbY8fvVmTgw2Big0
gmIkyHvYhzA+OIInp1ronxqjuWLDRqTBam1KxitgGZPlZjKXmWq/QjtzYk1dUMMPGhiMegqC1tMt
hP0FDIpOop/hOESsYO9hfuXkTCoQPYA3OI+Nhu3IAPFDqrGC0MuFCROgitZ36RlBj/0TkJzT4FJj
dKjIdgu+JyE1Td7dNym+HvuQPxpQhGO5ENY3JbNKd/yjIUS71933OBWEDRQbx2peiXYCQP3WunN9
SqzRf6ScLn0ag1vkh2z+/x5PSPu6wFogk0bIF8NnAji2Z34m/8ATY3UvIk+K2DNPfU3+aGD65KX6
twzS1pyHTXevZKFsJ0WdyNOKqF21YesiYWBzG5CP7cgHa0tiD0nDrKRg+6M2AJNWieNcYMnDS0gn
IK+DgVf6CLOsZPLdWGJRDsBMII9A27ubgOZpXbp1A9meVLjPzC1DhOsjnnd0vOduQeUpPo2Cnyzo
9leVAGq/rvk6kairD9tvbTilc9PsiNRbGd/r/306xnIoXg3ETwYrSklcRN1CQOMLPMwzFHkEbj1d
M0QgQdGzdBWh1lsQuO14sJWLrWCUbYTWnPgDfmvylZGfjOI6np5fiPty+Lj94o1HGHuYGMoANtyO
q1L52zwikhym5aR6OK2BvTTRLyHMGjRqQfqsAKWFOKVjvxkyThfAR/tSDaiyGnMPO3j4hROByMET
guHJTpVETmBeprJEoRlW84MIkiHVhtrySdL9ze+HhUvIJ+ZXDyqyRoNqDh9fbpOtL4WH24Ep7wC2
x/JAogg6g1jjzHOl0LRwLk47VyGBXXtsG5bWRI1khORDQg/1q2ReBNjr5GhZ71Hxsdi84ypQfDJj
GMe81u14Y4kAm3MC4S+owqAlaqJizKQTN91iZvYabKy55+eja0sMhkcz71BrHQ84y0NP0R8dZlVi
MHozThtQQwwmBvFRU7vbwaMYkWHbWfjNb+ydek182ROj0ujncuisPgBClgZGWG95ebS7X+SYoz9p
KBkNI2sVzFhzm/unM7V2jWXSwPVCxbuv+Cnm0iQlLo7GZxfnc7WxASKhg+cgB87AvgIhAzasNVsH
9ZkbO0MOYerEtBeGW9Yu/YMwZK0uBl3m/oJ7OAiY6YUzhSboJ5tNkweAjatzvHcvV5GOu4VGfLj5
QhD7I30ZmUClZzn5wfhxXUQmGZN5Rv8hopiY4mRMfpktCoJatLhMkL3NTWlAIAVrLm5nfw99J52t
pFmsaewbVyEWZ36lyjSah44k69eD3SroOjz5+5fx6edjxs97TaWWxxJvHIOFhnZ+KTiD43AGpvPz
g519n1E0BU0BouxtfHG90kDNLlMq3GRb+DZA7n5txarjltU3RiUzPnpOA2/43K/wyYMDam423OUw
lLXCTbt0pOWziGa8R4ILZTqunOnQFe+QJp7ZIFMWg9fZl7IzLu2a0R1cs5DXiyDLey621pjeXCuv
1vgfVgba0rlTVUZAEs2lWsQXc5mH7SE7Or3sjpQhn0ORiJUbg9J9BONuevNjDYrN2bU5rXs/HPNu
YPZbFwv0e4o3MQ7PO9FKD/18qCw+ErKjKcNNYTm/nvS+MFeSKkMD+RQ7o0IOSU5mtObYl++agpHO
n6Nzs446Q2+xs9nL75GTkOZljOKH4rjWCePl/YI5l7EeRJW1PyjIVy0/3oke6e2O6bG71hAnjyeQ
IBKoIrxyfkXc+eTwf1perNBEFMq6CBVMbYWkrLaUHOpXWGypBKWf0XGs4AHP5BsQZ3unPeN4bCKR
7rydLfpmAkMd5FkpOmRe3HXsoRchcgVgea0MZRlaFfE6LtlgE6efr+WUMACKuJ7UuV0RxTLlg4H3
N+qpQ0ECxjgl6JZQ971NGYZ/AGfoGnlD3lBiru9ptcTwzHwE5nRJ25IUm6HiFBokXNxoPQNh61o7
ru7lIoHereNHkKRqYh171uc23Lf2WmmpkBlxuwEiS1j4or6JGIwveKJiBfaXKQYRoGXa9+YRmoCI
kbxfyyq3zC9xHLyQRIS+pMh8jZeoCmjQexBaDjoI5NWB4BYGkDcn3/FLYsq8OPk5cXpqy3vNp5iv
iOalsNgHIV3D6mWzl/1gz6kwLmHBpOBuHv8oG4wlicSmy0FKsU/3xfN6+u3PeLb5VoqLkYOb+kBC
IIaUNOcIyy2nREzY0AAMtoN25LvMi90xEflbPlDpE7WIszFfF9gRdSMwjUMnK2vom5eZO80gKTka
WPLOWFm389tW2EpG6w8TazJ0e2/feUB+hm/+RlpgpiAx64qy7b9py27GO+qM2j3ZAZME3mf1btUw
2qdKt7bNL8pODz/UwTLVhLhgUn20k1SWMAF+xF4xs+DcwlwevuhhR7S9E3t/lu+K0dbQD4r2RGLH
VHSIHIzmSWl9chV5XSPLC+9Is86xsK7M7WUQ9W1MawCo8SzAo5ZIPWG0JZkZV3GiuR1/otzSv/hh
weUTqNTuz5++SHHhTFxuWb7FKqH2h7A5ofVifPJjPJGTE5/6TwDyk+vUrnaeV3VKKfV1qK+vtdP9
pg6U5T5oZuzMQbrxnWGCpvMtsyIEw1+QDxCmvOwOR3f2g3+IDzaafLcEfaCHMrgXS2A3j/2t4wHV
ezVGIirGvM0KLgNtKaTq+eH8sOlHlj2tJOX5KBvJ/iFDmwEkcorjbKvi5vBdE5jeZHdEW9J8Muba
t4YXl4wUSkzmleY1wbHKFxTblWsCSfzAsUqxdQSpISVRLA7/GtJPoUUvqG/lbuo3p2xazKydx0pO
Kvyuu3pShKNEhM3OjUdljzuebzP+PbLV4yEg1bd8sxmnffVAjXvUcT7Sy54aQXZdqUz3N05CdibV
ForS5sIskNf08Orf1LIvyXPEjqugJOfzTVz8Ihv6QNcoVozpO9fcDcnMBtKo/oBloxsSO9Jx0oA2
FX2OS/gpNt1KkAa56D+HIIltKhZ0qb4ht0S3zQmbd2lm6w44UMwx4urFyN/93IclWz5dKG3JFmyC
J7aXvXaCvFU+8dFJQBJSKX9x1q+3J/QebZJOSmYWDByBWoz0dYQy2YwJEJKH0vOzjIa7gKiirvkZ
1VFNEW0yXSwprkouWYmIsk8Cc/9NsuEE+zjfc23fc5bnDqzbBmsyjQ8cm/cdkBkE+M3Hzwv4Sw1Q
6PV/k3LHK4Wj3mo4pRpsUhD4wI9h1QQl3D751Vzb+7M6DX/lUozim3GkfvqdQJdoxfFWZk3zI8g9
zL4BsG2cMOB38NQGIpmrWtpW3Wq41IjiKKjoLLZi21KGzyroiPBE2zRhkeonIKYrq5mB8HnZLJo9
1CyeyDzTTHCFo40ZgUfJt5pu+N1ul5Eab08mzFqMXEmgOL0q2/sb+M4c2dW+K5eYq4yF4cp8mdYr
3EGeMvizvoUBHhDFa9KOR9/dOy1WFRQav7XdTSx3RPJlq8uF6T0gsGHH6Tg6bfx7/+VAseK7Fmkf
qqa3GgwAo2LulCRNifadQWY20b5fO8f19ntfkTxVnK/+fffUJ1Imq3d0U1cBDwJ/MzTLrcxVMrPO
aU2jhop8nJc36Dwoggo9GHF6YbKVxoE96y21D+oTWq6ZiJgbMoV/+udt37bbg/7IWIgnPqF3E51f
TwhwBl5hHS1fjm0XNuBLZVLomQsnIyt14h2aKyg6JRx/tsA43CuChxz1htWEo5bzmbsKhF0nRyHr
HOTrZQjKzgMB9g/bnTR1E52vkCnRZaDcpEtzYy7k1g7Smk+rUxuhWYJzWG4n2ikfkM4u6tINoBkD
Uj9bkhD9OmFYtpo6l9Ys8Mun8nHA4iGmroM1Zy72mUH89ARCLW0vVU1GfyQOUCyEm8ItTJQ5pt72
uDFD8KBBecoDMz43hlNV/BbThifEp2zykNyMWmT1WyjksQ1rF4QzhJqxjjv7urqiPmx/2P0Z6VLN
FPc3veSmv66Aj4e+ljiZ4W31V31kQ2r9KbHbBVZKZ/JHKTmoYggjiAzSTismIN5KXT0mpvh1Qcz7
C7mB0gQdS8uhrKtF8e+jyVj49tCiZEOajdDRwTgtLZubcgm/REuExkuBBd8hI2EOYzuSzkTIvtj+
XiU0M07dUpF6EZbQFPM6LDT8EG/IOWu2l4NZqOGwNm/jCf/Ci7eK9kvXcHIDtOOINeXh420JdbzL
T4qgdWLsMoowVOndm+PluXRASG2zko0SYVXDirEVjD4tcJA6MNxBltXpqvZAKuG/7ra2kYTr1vbl
FmmfELxTy5163Wn/hL9pnrqNhidoG0XacHkELYo7WgXkcz5cixh8DPSiAWcp/pDwFaRYyylK1oDI
aXjFrpP/jVyW5TVYd6P0CbVR+C5phfXsdJVtIU7ERDsVyYN9bMEvSJ1HxLoyEcVJ2Gne5G11/1Ir
I0XWB4eNyiV7nLMjX4rZnbQo+6YTI6FStjwkvb2mipb52uAAKrvi5iH1GMBSET17LG/dVpursYXL
V5zWG15bfeHvh23B05TuYeTA5USJCtAHL+FbqMh9S0NCYEImcwNMRAZwZZ4O8iQ/OJd8FlnvUe18
vw1onEelCsLBxhrHarF8ZfzGwlKYgP3ah1t2Zi/G9JL3H3uPGxdK79mT1i2Fg558LLdToXrYgtUY
6kexAJrZuGTmpvbzmxNgqSOfg6L0PQwW1/sR/gAxAvfoqlGxw42HI8oVxqVO1TG6HbG4Xa9srZLs
Zf2IVq9PRBXPujI2O8E+juD4yX5N7FrRRYtNxtjo4sEuhMuU/Dh7laS+ihTV2rC9ZrPBstMH5wz9
K1ugKKg64Dx3h5SboyfFJPPN5OO96FM3XR6NHmISBKYkPN8s0nSH/hwT6d4hlsoE4VpJWzYH5kXW
26PU5/vtmWOYpPE4W2qdXYRnHo37Bu9Xhsj33KpqZpgcaRvJvmXKyz+iIGr6BQxPPWAfyO7Wqvrn
OHDgXttZQj0TjJ9pKXJegfa/CmQVgNWt7+GqRb8D+ARwPDTztjC4UA5IWLQEQfbhH4cBfYdzf8Mm
+QeVOvDs034WJxe01Jgiyh1g7Zko6C+IEIpwg8qb7fOfObAVFhFfwUh/j2IvvnjBVoZFDvLIIWRu
ASq9zXRcwj5/xS2LvQdDW+RaaAosVCu38/B52cplSuiivmwo/RryvtcdCsXu9AEgG1+XQ1Hd20jU
WfGEiNqyM890HUUtHmN1apWNHgLu8uN5ON3wf+AsnUEMKGfrzkM4HtJk5IRgZ/etuJTYm87RI8lj
qT5eSq9Gv/kLsG42uZcKG7qcZOh1SmmdLjiQKDDpD/U8bfDYMgsg3d+JbaXDbCcPzmaqfzihkg20
EqhQ7er/TuhmndK+Kx1ADg30WLewsVz6j8/bwulsuPoXY9tGplhp1ZNasWB+1NU5HK/eLZIgEPva
Jc4U5bPjKGat/DLuLFB6QcZcTYJo+rohD+2QQQqL6lBC4IXLXZkU5khdDQr7r8jrpN77NKVJMWVP
RiqpFuK3U91QN/ljr1aGXkbD526SM6dpWt3srB5aaXEP/6Qdfy4zq93vrLum6j7MzOT/uuJe0YJi
3GO0gwvmHPWavACf++1eR5gjipE9JLxE5/ALvuH8k3N7cUjYqhmunLTOsYzPPJ5qSdvgyTBS9WYN
9ufauitWqYV4WsFqbF4/HB+tpds2NdWb+7HmEGtvC1L84uGh/SIdF4tF8/iy5bN+j3IvypSphQnQ
v/1EuNRWBsJnfGuN7Hz2Pm8BXtCHZkmFvXQUEgfkbJKgfgihDjUKVeXLvHagxzBqghcdz17ah2hq
z3Mu0OQL0CL/5HAWskTtSsktgFxiKMzwlRmpmhx/CwRkuhNopGd3LqSNbMW9CBBz7npvUaEsAV/c
V/FJpHazlRS18Ni+pGAfGpqaWujwEU1Z+7s1wohiDY0bHTj1GVoD1810e1Td2EPwITuEfUXeJ4ko
OdHe24vbEkpx1Jz2EeMOiyxapYGA6mY3a5dtgP/myz4/4a8nV4qI8ivNrfHoeFQtdInt2N3Ybd/D
SOpeY3SKYPSPq5fEf3YCAGlu1Eg0CivqM1zxH2yK7ySSLsFHPSDxRXcGNjXWLVkPrc4vfirfVY/5
m5n0ccm/f8SQ4atJZvwhA3b1HgNLWbnisomiNeo5LnYOuDdcyrEELSLsodULTJmS1n10v8Q5qH7z
MSt2gOb5ordCLXTs7ZlCYw5xlV+tfPQ1g0nUL471GmU6+Jv4l8DX88qsNmTeTbhOeAFEed6UZvZS
u8CbhF0+oPNUU8yDEVlembR1eXY3qKV+RgWqOwTbLuNgwc4I/uFOQDkBPVR9yoJMVPn7zfNFuUbF
IVkj7vdq9MKN07CVSdE5kqU3AZBlCCU88ybO8K5fXDeG3MlMsW8s7/4eSBiAc8nuP8cVIcGb+t7w
mS8EIOsDZBbUEyPuukR4wd/lJU/xWN711DO7DaMxU/MYyLFSE1FR6eEw273kn3CUloTLEH/U7iSv
lh7UrOQkQK229P7OwnIILTLVx9N/6Xr2Ar5/+dWD7g1w5g622tCgqsQv90xHr9aggWS4KBnf1hvb
NLjwwY/P4e7XwawXVjmhwR+M+sJoTprUkhtI7caWmmtdaJV7J2if6qatWMf7F0FFcl2c89X8TWhb
++3OlYZ5M0XKucigpY9uLa6I8F9SKxH6Eb/KFFaO4EcmHqGZZMWwr757fmfAjLy8zL6DTycCHQ8N
3ImD1K6u3ZuhnZpVjD20K3FOWsZpjs4FJv4c+whDiwV1iYc4aYfuRAHAWMZyc6yodreRYEBzChfr
zEXWqEz7zp37F0qpsv5LULaJ1BnOc+DVayCWlH0lDW8JZgFSb9JOQhECXNtBNf0qyIZne2GmZP5B
9XyPcm7JndcjHkVh312jO3MQfvFx5pk9ABV3Tka5mSTKYEZtvzHQgZP9VTEXASH+2miouG8EkPdN
0X2jR+ZoGmjdOrsGbAUnI6rhGf/HclaQglWl37Eo+ab3Cbve78bLSVwFTqTAo2ECOX1U1KeuJGOF
n6VabpJLrPODCwjB7jm18UoLDig/AY6wGQD7wrfWScS/5jUyPbWGW/5HooyzhoYKFUo7jbaYHFZO
HEEFiP6G3hNEOQwYqmcyMYOF/P74q/cW9B5bvtWJOOM9q3tv1AZYWR7jdMJW/rJ2R6R0Dh3q3bUU
anqfDMfRD1376/BsMUlFgvE+C05g7p68Y00W3JQSBblKddv7eDKD8PiM0nzoeEnQp6Rqb6o3+Ob6
FE/iQpTQWW5xccosWVB2SaJXpUrkqWd0oMZOTONikC5FNwBORGta5j+qip7DKGIzjkGCNh4IvWqD
2Mafz7nZYQFD/ebxp+a4yUnqJoOodPOCA3cMddTNon70AIAU2xw9mfmWHoXcxf8TC9rJxWtyXXkX
jPISpJcoRN0dTU2T1VgSL0T7EobJzSX5MvmXn2w8eAPkJeI9y/3Prasv59ud68L9+KMBJ7H9iwM9
+aVD8lalVkJy+5RecCC4Moznrvy+9HU8v/nzhVC7VP6JsKGdfBO4NUMz/oXUzLp/CJ57pUYcjHrl
hG3fPHglMIyI8xd0UcXzmq/JONr4pO3OmmtA8zEdD8cuKpzPTrsQUNYOJ4+PRKXP/2O0G82XpDSj
Bt2T2jhPuINbUiqD0+rNdDNN1PczsJW8D/9p8R7m80W+R8CCdC0rnjJnvl8to8VWXjwnTo/tMRaI
jyesbhco9FMrJsT6LOdO5/6WUBPx58CLJ9UVfQn1Xj6j1+ZRv5jNQNL8vz7FIkE2BCl2gmxnO+82
H0BPpXrF8el2/BsA5iWpWJFV/PmynkixHBa9CnhMu0BBA/ETvCv+S3lAHwpOPLwq2IPWXrH5VC9D
L5Nxj1Ycc90/9rjj8BnMznqhY+UG+8tKoHfmnkDhtLc+ZR1ojLuJBHlgVKSeG11wS7CtGrNhqSOI
prHBMfcrkAoivF/byay8VD+L0X7g1WGoR33wj1pxzZjATbcBz6Ljm4XJdfvrum8Wn1OB/4PIByvs
jC5KHe2+NMSJHEQ5aI6qMQFUni6nhJLKL43V8SPiEoUS15jhvUAvkYTaszw1UkIUvc/Aq/MQy/VO
abVN9YAtOA6vLMxYwJBgMxUGZ2YSyszXU46q7LNbwebz8E1su+E0wLNcwymfYIySI5Nfo/VeZUo4
sZXL/rleHhKcCmjw89GiHeLibij6CCMN8hWjYgdVo+nmDKKlKaxxpVnrjisxnzFM4vfDaoGpiRAQ
AuIE20G3Je9I1Z6FV2zAhi1uHCW/VMv2DgJipg7eFYnowTzlgYXhfwVliYu+VMJzk3VWNHpae2LP
5o9LLqTc97BqB2vnOS4+C1TqETAo4Wmbld2Rq4X9oJp+C8/P1X3oZZ3SMXJTYtsUjlWyDBzsL0Aq
7ACPteorM27J3N2S7LpmhneHxN+NTE0ciXTew3JeYZmkby6f8LyPoV5J/ue+V1Wqqv349lxaHLUo
HnwGkr0a7+WdiO9QxMIwxKAxr7Q62HIuLZdQf+N1qZ8dCWAE6BXvn/o6gI0qh2ljswmxjdg5JXdE
RUiaBDqxjVt3Lr4Gq7JZ//OVdV8NDENXkH8ShxKcb8U1RBT3QT2iuMgPuvqGa4vhj56oBprmRE0t
pWe2aBIs0yfLgntvw5piR7mrsmEBVRti4LN6sdtlgN77vvbnazi82dFPYRDQGThJdoKbTL6Ac5L2
IzUwTeR93bzMtvdYEosGe2WHL4ORCU9tC5fp8teQg63UHSVhnR0hLYgkkyTbkWwWNXjCdQI0+s6/
glbGmMoHhg1YWTI8L71Y0R/8AUq8sC9Pa+yefi01myDai04O43LVdNgM+j2f4YJzCW8w6mkWyKpE
KVD1xJCzmLEqad3S2+nCo/gUEnmAThLoichjwyA/f/hbciPVsiBOa88qWF3pr2G6BXOF86n2gKwt
9D+a2jj5jMMrVDErvvwbx2QJZfizZatL2o8x78qcUNTFz3CwFWwDqyvo5ZeCYzKzpEnvfyv9RV1R
VtghxDuCzppHoWI8nt1/OyPyosVMbD+vXiOOUbxt7EOzs4u9awMjUARn+RBrb8abc8kL+0iFP5w2
D/6M4CenCbl6wJTRdeNvYcDuuCXAL0zoMv8JSW1BZ6CCa0nCvDYr6uaSLKYzd2qMgadC9pzcpY93
mLX2tKrYwEaCneuyeEtPE8NVKp9wzdff+4vxvUDA53gi2tXWzOTozI3CKwkkRtLmVXvxs7H/Pz1y
1QNwG2cJWqmYC8uH4Tt99uyL8F9m6D5a3L6ODrYuGTxGBZyKRmzRAuUSdHIlIEMTOUSai8NztSzo
V6XEX7qNKQ9Z3WwU0I8DNny3zRZgoVN/okGGVjtVbJ7CFlxidsitQHaFa6kg7AX1988Wj2cQIpjo
MZca/oWYBFnKjUoQren0z5HdyICJhwGdoz1c1WT/VjdUYnP03PiIAoc8DjRpF7t6tCwfg3ZB0eJy
e5zzEtNTXRZ4ZSA2P/dThqG0s2hm0JUAkQ1d9gi/JryA86hyg/a2nhevfVvvZjcAFo01zHkGroo6
qC6V/v3GDS9XcSKQKATorPRT3nW1s91hQaIhtwcEO7UgYwiseOHFVmQDLJDV2hYYgHQYijvmyK6R
Tw2zGOAB0++Tq1Pk1BFGgLM7L3xjYC4cMLERh+tCWYnRjSgNU+us4x8w46BjYRjI1oSHdANKH6c2
BZO+9xve4GxASxOQ4U/mvFYO2qvrrooBoxJwjlh8YEq0Ulz37HFpvxgkdX8dJaWOf7CLLegWhh/5
DNDTkMy9pgGss0+6i+gr4G6SXYku+zcmSBsUI1LO/KTeqYRTYLJ8YCwq6tRjaR0SU++l95tiPrQW
J1KZpgzAk4EDSjtInWFPROfnCuAe2F3EQc3/8n+6/EijXF4HPwR9p5YPApocQuaaoEkQVCNUHtRN
cN3vzOecvLa3s9uTW1xp6cMA/tMlEFva1j+xU7WEwsv7BcdG6sr2cuk8M18uWCAWjbOMsZpXPsh0
JYXtg8L4l1NMni+AoczXHwy1JZlTKuLLg85aFLCOmHmZPoi+OQ7xaaY/NKjHjKRQDHclR5YTUW+r
OlqDXnnhQy6guCsuxzj3h46r8gyREXBUaWDSB8SHVRHF8TQoWFNA90nNj0Rvz5P5TJMNdhGv6aFb
hLnxncgbhuxQXJJZPY/15HXpSS4JEUMqlUA6MDpSxWcMqVAXtuLF9MzRBGAp6NNjFi0V1ojqpwnp
WiEY9cxjYBmau6vtnTdcfSD3hPjK3bjLm78hfNR7T3+Hd5+KdVV4kJ04PjVHnRUSjWE4+gJx7oXT
092kOGQRS/ZXw5lgKyvEz9K4tO0cclxe+VVAgL2TRVl2c79UnQMtKFHZBl0x209WA8piotpPYJ8c
saLk1hSLg37Za6AjenhlpJWcl8T1INgvRE839xt2SZ9LTID/hvRdcHiB+AHrLApn8P4kVYuFTxr0
UlRNACepceoLRExmdOgntuBt+Dv64xxsjWXHJp0bSi37iZOLXqiVMvHRUaOmyVtqyLhG4qsJMyNE
4T8L4TkPUQrAPj+ayu56KnzNivD7OiffqG5pySqQbPdNeH1xNBoIPmucU43nYTbLyYr/qbXhAuBG
ij9bYFfeyykFgced9JpBkKIpm0LzwRbZfkFJDGSaxui+5Wg7TYTcl06gFdO7FRbhS8s3KJ9J+R0X
ZUflK8fpYLMdom5oCp3SY0lKUQsXGljZpvIavJWWLecI/bhNxVu744Tnx+2NKX3+MKXS7ng8nTMB
QN3Hta4okjKmwCwHgVTIuEzIovvi/sHo8quNj1uJc0FgZQqO80Y+5c+REQBwOiEUM6ZY/udw33fa
ZxzFF64VOie9bS/x2wwqUjonQV1kRsxzfugRw8zpMcI74/K5qgjt8lM8QLInybGvZd/NhIEK7dwF
JFvx5VrQL7WXBx0DHD2jgcINRHgjhX3/S/rB5Pus6dclaF1M6Lc8tEEnMLiDH5gqkdy42LQ0MtDp
8tAlUHS3PdYK4mT2RHCvVfT0YQdiYaVQ4JDnZGLhpQmcNapBuCRGJ7W6FajrFMw6TyJ+0J2gGQyP
cJhoY/F4UoX2lMF8JLmKuO6EmVVdWSum/SaD21NC6vq7FcV5gJfUJtnq9LnEyoiJeR88RbeCHNKL
jylQzPWKHMeKMMaFXOvjRaTXL7GdP6PFtabhauVLrbMzNHTMjSLIUUJTQhbtBTcIbYAuUx0ghOm4
yKwMpEB54h6ejEmr/zzN8b2Z7KBr1zw6xoYTWQgRhXn9PgtbDIJzYKamcNbGcbfwwiTnhpjw/fjE
C7TadANg/ehRQ96+vm/JW2AFutLPoz/f5E8BsmMSB9X06Ubl540z2Fkrig7tmzWg/eHtJgaS7Cu8
ojo8Pkz+1LNRC/E6gsYhVbfZatoprtk9/1mq7PAUvzycu4fG+XQ6FK+NKEpAJoJOXTJxHKHL6igY
Uah8xgwo+kkAIGQOgJOJj8nn3ONYM3AuI2l0E2eTEOsVddjFcdxY+X/z5DP53Onm/nq3MNxZXs9r
nVag6KlVCk6SGEKwyZ2ippSBkYsS2wqj+6Dg5ixmToktMLC1hPX9gVtHJST8ytbF6LFkMCSoHUZS
6fVSsqZ33jwm780ushrONguPKTIkgkcBHfQ0Om4Xm20E+bWkRprzgMB3WZsfRej2okCsx234j7Sh
LYVG7Kje4eVk/whAmoPOim2+UyhwX42SNEvp89NWOzJOAfRtY81/zP44yix4+8EKRzX0VmOwDbmw
Nj7J3kryhc2rC/pS250+4y9W0LVtomZZ56Kkx0plGzmn9iABj5nOo56Wzu89X8vewnApVDNg0YEs
HL2g1DuDUi3zP0W2OSlqIT6z9HAEqIABIgFA8NeREI6EjJIywq4UTyflC3ZISqqLzQCBZdydgWmS
Xc+V9aCa2dcdnAt1/Le8x0VU2AaE/7mgZCaonL/vOznugVddFr9laJix3en4jyQ7b1uS9p8GcjTw
oBdMyLHv/eWGjHLcX1ELVzQbFvyeAwbviHIqPSb4+LZuwKviPyHRlxypihHyQKgv3Gyjh1QDQQ8C
uoFmZhIiOxrhiTjX4eQMA6lH1FXibAUhqtfL5ER+SwXZ4FOHj4RlXA2xSD1LaeT5Dtbqm8tH7QFh
rO+mwqHQMn7Ni8jyNETA14mgcRY9M/XGMb+lO+IV/5jNC1kVO6w5NCsZLIZ+PbuuJWoEzEUzNiE5
VDQSN/mbaQMkP9B9FMJMKZln6FoahJbHy/t/7IJPL6g8zApxyP83evmvd2yTtcMRdSGtC7/tkY0F
CLG59eLBvhD9EcGY4V5Qcc2uCgjHUO+0YlJ0aiDGm3l0savwSsGPMrg9v+rkTKqjGnu++xVT0MuK
LogE9QincDKf1NGd9nW/+0YiBOPXIgrV+DkEzy0mnKM6p3nD2Chveyk4QuZemtgY1ejuLcUclhqK
/U8hjpqBDCsNbkaGgXFSWZwjfxtcEIQYNFTHV3jaeOLKAtbdSXMcMMB5sA49eeE0AYyRS4fnAuCu
PzjZYIwe8+E7lDesmkzzggQFihYs+stJHOXCow+wlN3ZJFi65g+kMH2w0APUFb/wij6RmXCIGkPc
Dbd/QZfh7oThu8W+3H4YrEhb02ByMjQNfh5KPxtTDtnVVEa3JrDr43cVSPyTIl+kzWLIc0tH9HQq
eHWOuw87rENYcUykiKcsiSCZ9vIvT8b7aY14hcNC6wZEJAeXBv7n6tq7Q6g60f5MM3kMdCwqmvmY
bC2z70UHp0NJC8uV0vqmt+8jBK+pIloNFRj+U0Dgv1w2Gkf66V6QU+7UZmIv2wpBBhEX6o8evFJ1
ttjWHgEjwm6EwLt6s/hZ4g3T+POrKzzQHe4A5NiK57r9amWqBRVReZT4WWDYA7Fo5FwrGKJ3UnhS
LAaONRVr6LX//z7R9A3sk0OMl4fFGgHeL5G1Q1ivEV8DdAvpwxAhS+OUrmv2LIZ1HIkypxWvWZXy
DPM6tETUIs4XZ0OTsGiNb+Mo0/BHs95o0m1tBCwSA051QNWbkLihUI9dAu7qiJAcKGHnTbs6Dkas
UFoOCyKOMnJZr89aj3UlfmmueOQ1JCxUr/knlLgvsAhDvgjU4tzTso9KYvmHeQs+KRswomui2+la
TSS7gJAT/wKqzt4+Po7YkI5OVnBJdCmRiQDxTutLf3S3kA0qdUWhHCwiEJFRHrxQEPLO0gjtwDU0
CtMI21a4w1zfcEq2a18poty82k09uythsScaRbjaBy8TNhe2HXKAz+c8KJGgkMNUqQj6mP5Q26CJ
qUI+qa6X7TS6zEPiTjKFnFc/+GyRWbe1k/wc/5URDIp+hPaunHD9dMoZek6QcU/mvfAJCBHMC7Kg
j54cKzQKGV0Az9Hhkd1P1Xu7pl6M0deABYmkc9UJ2E9e9DY8jxlrKeXM77wgQRMZSCYy93bde14X
7I+1GRbD7dspwPmZ1Nx1spoUSSWL7HTMBd3GZ0IqgDiOKRl12HTNMtwM4MnX7S1ngmUNq4q6wTyO
o0ijrtF2PluNgdESNBrHV0GP8NJgM1V9LfldgAn6tVxG7j8BKPh1k/u+eZ4ke1Uj2qlrG3DsZxas
JzGgeU45N8vopoT6nEAr8RkijY3EZ16MMRwHRRtTWayK6EJZfT7061YtxizuRZ3nNLADtl3NiQMw
90O0u1cZK74p36Vi+nEFgKF96UFXh8o35os2BD14IJwtW6gmVirXfzJtEHWh6ZiBC4dfNh3Sp92Y
ZcYHRFwZjt50t9Wa4YHVrDITGeImzSdowyePro7t7u3gejUH/UozpueZLBmMwQWnV4XIb60ty9PM
8ZUCF8cetrsCrD/jcbwdtcGkl19mnjY06CrR4Cm+xkbuanG5fai4b8jd/z2Yr6F6McmZxuDZ2mFP
3Qzt0e5PZ/tVA+UoyLBc4fG2YJb8U0cnJHOIgM9aF2FdBIO5X+mMQExufKqZ7n7Ub67+CaQN7N0u
CC0JSA4Nl3BKeLL1KX+2wA15YfRXFUrdKOwyP1GlqiAZ8nqa95EaQMWsrTQhHu5jByqIxtvdmsBi
N0X08ePXPVbjgBH822SuqnUkueu6DHzKN8bP5LHTrXOAWShgld4WmypJ9MG7K6/aglZn5oRXIJiC
oaS+zipggttX9mV/BsfWqaVPsNYrgkNnM4wBqOTp4JDYF1kXnAilKrbChCSsT4Wo1BojrLg+//Lv
rhVu0EBZz+7EcrN3o1FayBA+GIZ+o6AvFv0vpZaJ9d2yRk+XlYmoChzuv1WjX4rfYBh7syh0Mb1A
l13IT96Ewc6fat2x0lG6ubKZ1gk0v7v2uWvqsF/V0zEsjLZjwHDA/SyrRBztkQl3VFBsPn9ec/VE
seveHMqsR96VeAK1hh0K/vPt2FkPlOmFinSvnBwq5N+tnC4mM/JFZKS+SbdU7Tijp1OGAU5tDXrp
y0ra00PYJw8TbEE5qqwoVvIfJpb/nXTw7t9MjjbiA8LG7xkGjpoi1xCGSSSqiiWFNRYYrbO246B6
ipluruzOrfE95hCzHLSaRIdRVvfPP1SADdOgxeauq2+9oR3ksY1dd1wvOIw4wFjQk+Mdq26hvWMP
cpAMcIC40WAedWi4WLW7Kbdl0xMBZfsEkM4C/jARbs7DLsD7W8HKz2blOLATg611kNPGtjxuHyZh
3k1xde6ogtWJqdNroCpaODwVsm0iIfAtcDW/dg8Lazjcgkh9Uz/eHZMJ9Jen5zwvfXF0RZGDW/Yv
oMLl7yxho49qwIsWxEOSiVkkvoNfafS/qYq1pdC6sINlnKInFzEaD2LHJG4foAZPYQZ0AfgfmSo2
zHIANz+Y4p8eiX4Fzaz660Tu3UOpNp65s51uZIajNkMRIh2d3WwSF7S45sR5WI8pOnS6h95mq8NL
li8vuBs6QSX6c3+bTL/KFPw9J4fQ9q2nYHU0KyxvHR4qejWtiQZzdsxUMyDkLUd+za7bJqgTp3s2
DPBilXmtlCmTXkSqYtmJj9IxNrPScyZ3e40VTfw7P+nlGQ91j54YF6wlX/lj6/t/AynZzlo85Tmt
kvqzrrsmv7DOVa3eKNB1Ugd5mRUkEN+E0iLcg/qh+nnCVOOi7CmmWpO9dWRv+kqmafWLUmBPuer3
pJ76rU9SOsWml+dDfegHa5LvIUvwIKL5xnut068bowTHWQ03YyVRZWkmyMg0ZnncNAjXSow7j+oQ
/0bVdWS6UwhbaLPPYlKj6w+JrcIYi8wb7LMot2wUEduSJmAOe44ViBPBQgDs+QW2S+bionygHUf7
oxZGjvhilf6pcz5HPezt4v9MXZqQf2SYffH7KrkBIFECVySy+Lku5n6Y6zmmE+WXX8gxHbcj943T
2FTXvm0YceSOFsdR7rGC91U9Y0ni43/JC06jZXlU4dNhjKAnXLPza7tGEFwNewrtP6remgzho1Tb
el3Yb91hlLXEzKeloEHwET85qBiGS5bwAF1eWNLjJrVBwqxYWq/JSe0Tj33zYJrZLRKLPz/3Rqnt
yjrEi0RxM3tlsg5sYzj7QWQ5jXPkKHxkE2lupPkMusqKJ6mYP2fNvZjCXmXLYo3Ss9ldesyZysEU
bHB8ayP637YX4Yfbt2gpx/0Y82x/eaFGDKrii4ZQDJ5ycifU6saTf0u1x24gjKv8HWUR/AVG3vHR
o7y7Id6V+IBa8O9Ze6mEBCX9cF1MnWrjwqq575K4BaAoDVp0aEzqahkc+gXFb3zUFUuzZvfmVqH8
P+kpqEZ+rzSWtACFwJHNlauWWDpSXknjdYFudp0eszBbAZRwUAgqAb/cM7t7Mv38a6hoP3ASuIlg
bdw2qmCNV7EASVZBM1Y9W+YB38hXZGlpubFYlS95R50qXGZkdkuyHwWx48bE8Nr7JikgSjlNZzl1
tcAdKjQ8MON9QH+WpcUUD9+oeEga1uLeftB53frbgxiovwRrq42fWR2u5Tyvv7gycHEkqBcdM8hk
IjFJ8Eq2/ugcxosRxLr9tiri6Jo3UZt/OIo/eUGoq2xrw+qEIaqlZFrVR/2mddYb8UR7ZPvGfvM7
FG05H+0Dk5Eyu+yOwTrGZd3nfXRuL0O8Grkb9sWIWFl5LEcS2eaQs8R9rk/2x0IDTmQoh92H/NBz
8vRsnaky0t+waaMhQxAtntLPS8iwu48t5YH1+WDkSqhSlK+T2BoidZuSYwv7pywZaAgWeRmpZGzg
TkZEdZEXgTKDE/2ps1iIBfO/SVcbwX27bkMbF4Bl5s2nwFsitR8bBS1BsRy1nn/2T+rRSj4oKvlf
jwkDR6F+Sj9EgXAjwKA1dDJTMZ3Cjtga1q5za5nnrs9JjTCo/L6MRHgJOrN9gjp8fbP8MB7tVulc
6hGJF8GBmhBy2C9Mfm00gBVWuMbhbQ73gmyLiN1Yz8memEZ9HTDloA9+Z7kwslbyN7UVNzHDu9ES
5p/VSAeQuxtTeFFCKdhTgzg8DL7Y506gaumqMXqV2OY+18Rz5WQk/XI7+m4ngwEkGc6tVBGnx+LU
Av29RrJTLCQWbiIW8KQjer/ViKzDOzKEamKX6nyOcIzOTe8S/OqMsZQ3mV3RiI88Ni9nCxHmpq6r
a5jn7ohU5i5WwayjHXoTDvkxtMs7oKS3mrvjRseS14MUjWW4TjbBfHlt+c3lAQTvLklrYxwZCsDD
doB3GzfY51mpnBNrQq1w/+2JsCKgXxLfzIn/6lsqdrVD9rdVo/UfIAAs6SOngvy6iKIC3pSSB5wJ
Z/woVTlJHHMrVn/5KY97c9KrDTGYqw0kkc0AatU6pBbJeUMnrmf3OFy6kbqY4/z3OHBS8iCXoKT1
mKSF5r7fF5hgzzRuUQ8OiNIOxt6oNsD2pjlVfHxZrI9NdJwrXEJ+ohwG5mKPncX5o2t8q9sMunnR
++DPC7M16tZoWKLVvarQxQwJ8B+AYJIl4lEwPelvjBHKGH0+dgmAfjEPzqlirBMcBtZQdlqMjKoq
FFXEI7igc0BGNa7BeSNV8k07+gOu9WLLtgDRn085EvB/kf0a3yrut142fp6qNTe5Vc56WlYKyTp0
F1i9P0+ybrBIgVjanmFnkuGJ13CPK4BdiezmHnCvV7rA2X2bTOoehYBFNowGiUixRMdwIU4pf+2z
3JZxlHL9tEFRLRjE+j90/IIVmOORMMSits4UuCs/86r+6pxLGV71fnPhykqdMDGtgorEcp35ac+o
vu79sNJlmNTPF4TO1rRdnr/TuDflOQCvDAu4UN+r7LU98U9aIIVCYxp1GGxNwcP1F/e8rDGKrQIR
Op1t0ApAwWf4GgbQKE8G5L3aOgEkP2iVLQPvFWOPZ7j/IJ76kIlyH8f/n2MzXMkW2ftLX/863Eyd
egNqXcDspiHmfgPnWbYHAr+Ri7FGJPEihIJj0z6Klui8ng8HwR+ZxeXyZ2Ibq+HDKKbd6BLToj0E
xMixSjdc2NfHJZofoI7Ekm+1njP4J+u4HQdU1qwlofJrDR31uZksgXMwRQHqgtGuDEsW4lmLU6FB
5C1mo4GkpKCT8qVm1NwJ5ZcPeExPZICG8o8ujnmuqkhLekP0W7Zs70IsUMgR18pUVBzO/zpz/DM9
3fGv8PK9t7TF3F5wwhJbJNiQGhO14FqTr61u7QXf0yvxsNm/dfnB2HdjtKqHQMxGxzq5JPkza94f
x8zKDq+cFYJU5o00nUVsEUpqfdSS0o4tU8CkA75mA+U2dInrQ9LhOvHs8CRwjaEMJogdK7Cpyulx
47yXxQ2lheKNdYNki2re1ZkKWsBDs0OUgi0lsjMz0v7cG+FFYqzpti1BGitGyMa9YqAXgExiamrU
DxIsXKOY9UZppRNVSOH4ThfYkbWaYgcmRyx8td/jcadE3wt+5sGtf2vfuZgqDBMClzdW8ygU1kMe
HRfPU9bk6ugb1UEPFefOP5Jlfr+nywUuy4I8wqTqrOWvPi0SH/J5LGT+D5PTgXdalKuGXXYBAvL7
BfUpVHBabjsEE+rNKjOfopkrDGolIQv5hd7LGZ1HjhInGUhcmojDvPz8AMfGDAyECePEPLl3mjsr
OGP34tPlPLGViyS5TMXj5VKFtUzyfJMw+nk3UkZ3vu7Ah2CsFMNh7qd0Sm0ceuRDAS9Wf2roDQik
wlHbDE8wKXys92KuIkivLDhG8khI6PiK1sPqalK1CKSVrq5wmb2XmvEFSr/PCZ7nowAaAuz2ZDjw
lMRvFtnOfeNgKZKc78QtLi0VwTJnFpdQoFLPIq6NUn+UzDk0DmJsmtUbNWisK7VPQAKOwDfcvJ7J
bjSkxOuKqJUDRacmFtQ3jnMhHyTmH5M/1W39Mu8TJ4e3bIpl66PDJzThSuqIeO2Ja9zLfzeaZb8K
HHx02ZubxzjWFepU4MaLFBGtz7i55OXPN5VQdxUMEvhmLjfLr6JM4+4z6+tc8A9snwt4twLJg0uw
aSPWz/Cz0lX0PDJL4iNipbG1Pt3msA6cJ3rNA0wHs6oN3KLh8oA7IO3WqAiTRWxOhroIRe0RIWSw
F6kCzTxIl+MZ0v90TICRotP47rCP6FF3tSur2R3xEuhnOkm2dyRB1H/2SADYbC9mLkoBgRpqLuoc
sEs2X+b5At2PJnpNqxcJpS2sCTRyVZ1H7oVxpd74TOxzVIQ1ThX/I8bpQ7bxOcKxO/7aSpcrbz3w
DFhypsr0sf0zEKTxz0MoeIwoDp+rNJ0EruAplrGbp418W3q/+LfZ3cj1oYrpZcV4Y3W+pnyrWbp5
5nTEBBCGzxDkC+ck8MhTP4hH9vAuPtpIH57pREzQwMBKlRGTNvJNA0Q7VXQIOByDulZ6suUydgUg
kZ5qGL4ESzJ+iTkw/afjfE3kRUfmq1hkhtBFREZuxE3qpwlnxpBuqUxsbkRAadBATIeqgUbrgPS3
XVQ10+Hc/rvU+3w82JUncqVnvrRTaqk873ljSyt/EQXnsiCjsW6HDkBs1VQyJ349Kmkk+UNBRya6
52bFmVIoKIuysG2N3bIOXU2qHIWEZO8c04nYXWy9TSCsSpWYtn7eGKV/0NdyQ8FUwYcu/Girv2tH
1zxc1TeMATuIMsvjLRj68xZTqleX1fljNOHrBxWNOcEg58eb6ljep4CQ0aWGIrLFGmPqmf3jz8lF
zhI+ZC0Pk76QdhRf40HhcXgLofB+cOv+8kZQ6IICR0vdLr8FrAih3igUvw03gmZtvfmj7AuEbI2V
1bJjKV1+/v86itxNBKDFlaLifZkWPwZrOIS3F7vwDo7d3Bo+bCqVwBrttVtgMa7zmpb1jU9/ezDE
ogzD5riT668BlPCKeYvdAHhWeb2ajHr+GPZ+BriTc76SiiqjmbvD0pJz65LW27IKmsp0o9srZw+W
PPwy7bDfflvhXwDUvkYkkrcsfM/mTkv+GE3ZhZB3zHrAjIwK3IopIhZlCDyUjN3/meEmjHm0Qzbq
jKjo/Fw6xzg3VJJAKLv9JrxHhm77cgtRMQKORn4orTksmfj0r8qLL/Wr2S+aKpiIToD2+rUaiXrH
F1xWlO3sOA9s78miGGTPiHR4D6sVdqdSIONZvBw8sq+q9DDb5msKkU0XBwmMxY+d8Eeai8mrmkcH
8LMwez5DJVst7SMhsg2T8jy9Ksny1suXHB3+lPi1toYHa6m7uh5tZ7zDlMyMDsxDVGAE6uNdyBgz
Q89EpX1cmb7L2Uq7Nb8kF+J2zAqoYEdfyUZSGcnVdXXPzsqblwZTn7Ss+bkPIKksZlFzMAiKhyX+
6dd8IpIeqg7FLCKdMYhiwTwiupqfQaa0d+T6ZasvT11RaYsp9xR1g6tt/7EgpY19uZYIJj3ayKH2
PytqHMsHIPOGvZC8r60x9OnlNhaXkXe2sRGeEb4ZqMz3ezr2rryMrKAYU62809lRrWMrbbxwkb5c
83HLbhg3AMStz+WZ9KCcpwzlXcavzGQG8Mq/yj6cGDBrVFC7W/ik/J73H6IRBfkH5n0XjarTDFnS
qOHrnjSlv9iB1O6PHvSjM/yi2ZjXt5mBa8gEV8/0kQutcY+M6VOrVeCntc/OZQzUxDuRsx8zNdIu
SjKohSMo0E1NPb1wRvqfxT5Z5A52uCUDYImZ/Iy9RtDtCJBy42Q1OXPBAmXp+H6oPX4kwrZ28KL9
eqm8X+N9siGklwueVe+Ww0fgBjIQ1q4ACShdObu3UqNZXzHX5BA8mMPfd0UTlHRxoTk9k5FL3IX2
6poukcLSdpw7KS7WfPxvR0AwASZ5rpWuRuQydmevExQqSQC3XS7JFECNnRIKFkmyDpDj9375cXuD
eoYPkTTZz9wdmYrpI+WUqjek1/Yc6lmQs4hu7mTdjBwpU48I7uurYsYFzQ0fIjKkfBGssMT5reCi
SLBH25PUH7r8DCGv0m/tiw//xh7gMblWzU90a+0I86ZDruAkawdXGab0CaajNJZnbcve0OaPEUeM
+ZIwPS+YEjorL6+PLyFM21yic5vmszHfx0ZGhj7jNVZGolpXW617rxr0+eoSK0LmdXW2aTeRWyzg
1ABA4CG+cdEO077j07tpqVw1S4s7Cv4+dWoYS55rshdhIbYX2Yum8Jye87qQRtGg01dKNk+7n3jw
UKwBODx8nj3/9k/4uQCIKNtsQeoorHJIkg0psg8NlbsigIXQjd/1mAjd48uJdkkHZusUg49a9KBv
Q4mJtIuuIKLtx924BrZpkIZ/O0vk0UbI6ASvyrfsJpffiRDsHqkMO5X2uHQwAVAj79cLfgbA+4KB
9zRHs58bSYFRAQsgy+EjRldldsGrAKqFydpgeWtyF6Dz5r5XEG2RZjv+199uJF56MqBWfZbL7Gww
Y4iQr+dVbR7YVtS76n0mxZo1H6KGAK8S1cioghNfD7M4dRhbnblaFK4E87vH7RH4aq4eg5xmJbr9
nGOGx3cTSP/czWGVt7g2jfl2oAQX61kCd/4sC73T9NAGqRHGTPz2Nr8VtX1qC4GnfuNrAVScrstx
+s+UQRE6ygul7wKe9YtOsep5EKg9nf2sVcZPWE7QHJe99BcHWDrMVj7rqxic0cU+eay23rHMPBhb
i2hns/cVhR+hS/Uxbgxj87xJTfkRFD1ta+/nowWUATVRbpffVTR48OoPZHMlnAVhYYMLAt1v4SIW
EZWq0gWPWmJhrbogGqTDAYvvwnEzYyBgeC2ELNRi/8JieG8mu7Ix7BH5U5Deg/Ia9XP79bfXAVJb
rS5X/O8kceEUyTUgi6+m8ruB8LbR8q4brSEnYG5KjzDZBGVgxiUZT2vF2CMg8arldgM4I6ETRQSe
ZYQMj6sWAKDuJnocf3DL54NOC7LTuLkRk8D/mNAejDM07mhwEn74h8V2BOxOwVcvjFVrunEzNt6g
K9imhPI/37UpuevobCanqGsfISwU0NxRmcFTfay2fPeNSW6M2DWYWaMlzG5uiLqJk7W6M5YhhuI9
OR4guR4dec+LuahZGhd+KKXBzWMcAw+pvXEtd8f6HOi50V5UGUvWUh9ozVlUXEBgSTDO190DLJId
H8Pkxhyet4vFgJiP9+mGODQz5V8FYkarfDNGxgp4hY+OKyYpiLTGi/tycgYmIQEdxRbTsj+G9lga
a+nMCrrSs5/4NjteP1E1pxzeQffJ1ZJmx30POQ1A7tADvEUJZU5VTAMHN6/hMrC4a5p6BWFS0xYB
lB3P1dr62p9dHnpVBYWoi381Uf5G1rfPiP2mtXPjxirPdGBqhTE1MurayH+kp+LWQzM9AOor+NuE
Nkn1l7I1KQBb5dP5YOOazlbJ94bxD7uDHUavQtfsxjtAvn7BmzS3+eS21fjpRBhcAkdXltt26PF2
ASUtV0Ku3pJjNvUqLJ6f5zDxwneu8kVTi+J5ZvOzq9BMVqcSN22wlenirtxsKFkD43wpUcpOzAWZ
f/y3hy/SGXQyLngUXiLqLncXEnTe88EOEA3A3uK/MZvg1pcxyAfLSfg4/XZx6HqHPEA/bo6IxI2B
LRTBsY/KlUpB+s2h5I4MYX4XYwEUpKctnZBqFtbmNrNQD3toy7dIBOmd9zo21/KGo5vzpNMx2Mjq
Hq1nrmXZYqwVOiAUCH0JnQa5qLhSjPAlDZJuKCyM/cDhjHd05ZjzyjWYcVewrWWmKMcK5Mt4dsNa
xzV+2DWV2p3ixZ6Thy0fm9ucBWJkTsqeUalvGOvtA2e9DmNsn7+ZTBCnjdaNmKjpsHfFfw1K+IoT
qlqXeZPtlWNMtgK6X7cuXZ2+T/CJKgvxkZ8gX8V9f1g5nm6CGWxwMIGmer1noFmKie1weAoXHoSC
MimJC7RfButtfaqqkcRp91LbvSb2wWnQtzN4xC/Q2Uw/I0yIrxR5QSWjOSuMKoO/jxrv7niXZekL
5ATORs6SWsJ7lsG28c0MPvLMGCSJfMHQKni58BS4O2s5NNnOaW24VyzJJC2gTHuQn4xJ2gyaI1v8
l+2svFDqSHjYmOZIwPYtQA4tg0Iy75JI9EpaHsYITWP9+eSb+EAlXjPa770yBp/QWJ2PCAg9xE5a
D8v9hS4b9ZVGi+cEpq/gxV+/bcotyovrIyE7EeAld6QllgMhx+QWASaIBTwZkwDErdQ/8zA02C7O
hv/9ktU/pKlvhoZ9Kb0FgoctRTh5pkTOKMs2WhG6zg6pXSqZUxMZY3HdK/B484l77Uo5lrVJ6Tb/
5stwsbjd0GLU2uuBzalkCYJBq/JqT8+R5hkmDLvtI/syVGA+aOgVjyRvWD1G8o0Qcp8PXdLqcPe5
ZMPYBECejhb+UOBUdZJgBiAqN3S/YIAzKEyu76dTD6cVTQCpWuIlL0cFOonB5MqEEQyQYurVzo2q
XS1myXweBta79LyG+AngWeQ1WbquXkKVqVf+Jqq/MFsepsC0rm85WcRkI7uSLdFF+iGYvOiRXZZt
vMe8Sw1DOA36eEcTLxiJKCumdOrwlWzEH7NUvYMkRsmb/0lBUeutv/61ghwlegilWwkoASB+/dnh
AVEEZpeMfuBTw5l7seVZUQq/4GNyzx5IF8wFSq+pVu0YLjYXgTBiveIViQpeo/oZbhduhsiUKFgR
6fyFPMFuY6LzOymXvPefJLgyH6DpF7L+5CxkyRaE68NS/2GHDWkBZmp/iryU7zRwKSsBZ/hfwYxd
9mvBT5NGjHsnpqk1XxyVbxUF1+zJQ68XhFwkk1qs6oqK90cZOX7dk35IbTBnN8KqDzypZCjBFkjn
lYQGujuSunFyGlOV93OqV1KB17aBoqL5AMSqGRKRLqxSYAQ+CNvOHjQLzJhtMJiJ1+mYuCTnsb0q
eUWK4hl/bUFqS+MHLFBUDYO9hRwB3vy6s/gcDWav5cTgDRyAMxUnW+6QfxXtyNuQOlAJoFYEKY1U
fT7LSt1oneiv6kn12LkNPzvs69PTNTUFa+E7wGGH3qamTiTJ5vmOxr5k35HxYuFKNDJsGV2G8NFu
2DyLtudPwd8yiA/pjmWa+Gqy8xRjZBQLAW5rk6wj7vpqo0bQumOpBdJgAuHIO6luQEIhsQ3In6LE
4+DOcLVXKXQ8sMx1PQVWvfptYfH+VlfG/7RIAIfHXxjBSj5iSfmnJxRoMjRmmVo1z8E1s9g0GCiH
9ty83Q/2q0vrWmOm/No0gGfSZnyz/sbNumO2bgnVQ0iKJzQNAqyOC1+RsYbZISzB4Kdj0q8+7Hqy
hZueO+hlBbgHcVSNVrJCwAyW3qLzXisWFL6853ccoCZgxh7NmN7MMZqqypgXNC4dxztTtJ3I5/rJ
DuzmE1eD5nqjNgrH7aDxC48zLnPQVDst4Mw553xJZl8+aFrlga6ohGtewuklbBXTxDNomMzqNYID
mb5TvsYrlVu6fIaZ6THrzYrrcPjRwl5FTlrHKuBUJfvuQueJXq2TunVl2skYstJQ5nBAqJxej6hV
/LPMcgh1QAMMixNWfV07igXAvL12HXRYxYXb5FxbwS98Dp9dGhxybkFbMETz9kt4UhCbse5arIjE
Hh46blWBiMeUuZBJJqwzRBexAEwqMBHmOqVIrKWzmB4htausbZnH0c6+ukLyeqH287urIak/mW87
Z9IJvoyFOuiyLPsaCLstPxuIHpFwnU71DtyE+ZJ6f7tSOy+mpOmlp1H9NPV7GPTYAzlJXwfRGL4+
nlLh3sE/aSHsY2ZpZTb3jiUtv91tbiVrPvfeBEhhPVvcoyjjiprl2kFMzXf9z5rpwx7yZzgP2JdD
Dk7wAwTcTGJICH5wJTmWKFxXgxCUliwl+5XcOjjTRm1Iq6JsIbF4SbB4UqscZ4khv+eLLHKu3Jo9
ktCVLWB3OYlLq8Ax6Su3XMnWrO6m2Mec7IOlo7nhdWpOg4+XVKq0D78rLjXhC3lZFeOfRaqGVSRm
3EQPOzOxwzTWb/Db+mp0pKCbtEM+YRWtFwJrax30UG0SfwFi4CPwNLlNlGJoUmxF4uXvTmCgYdUF
E9259XVfKBpaujK/aZmO1KVCksF7HbsZcfpzs6+YTiAPvF3GOvhIRs8cptzTFU7jfLrUNCYZvC1u
nfY28PJE+Zp5LjDqWQFTL3+4yAspn66NGgY9J0+45HBbHX7Ia0Y1pviTDllN0KGa9ATgRUGIfCp5
N4MMVoBY4DbUYmerXW4nrOTnYzPyZseA78fXyG0QTYf4UcYPDOzLm/NQk/R+SD1DbrbLtsFmLhnr
Aq4wmJ0aRZ+sx3eQmkTa0GtdQs93mD2qKcptLkf6EJnEwMdltzDhxZxAxbzlu/FXFdccxwTe1kMR
NYxDdZzFKeFVJBMU+41DVE75SlZCv+tjUzl907qeptpiRdxjyPchHL/tSc6YzfdkoD26v3w0DGPt
jTiA4sssUDTziELXgpGtsmmFmPdALQottP2ZWDoGkETa8EpiSqxSlS1UQt5B8A88V7kj+c35yuui
LxTVlyshv7sKzMVwv800fwuy/sCDub8DIGiVNyyxyABoQYrqi/byc/9XtYStXrmGopXgeZsEgYwo
LSYVc7qvjwxylBQkCISMjiG6G//aqmsjLIAhu3f9kpbNt7+XIWOvR/kWgQl6+NKCxwo5Lk0y3vfY
0SUzVkSVy03SHat2ZmgBOroRHps5HuqRuofGGMg5vmtq7LGnpKVjmRD64+CkQCRrQmlhUHQzmuj0
HGqYBm4RFETOXx3YX3v5BwWuJ5lSEoYL1VIWqU3ITQGZ5hdM/6SEQTZ7E+Xy4JwPOQnedMK9fMdB
MOI3w8CR/V6beXQYyc5s9MJ+GEgD4AZws4GSteIEB6QFOUTP0L0c4XpnMVyVykATzUzwj/E15dN5
6iCl+puv25C8S9SRTLqFPD8U7xEUKp1ByS7FYRxH3H6T5pPmWnJJHV3zyem3/A6CeXdlvsT+LXbO
GD6yWG0t66fJTBtgVmKmpvaMWgCW0/O6rka1amf23d4CmJQSTvu3JJ+znqvPD4XyjQ4LglCUqsq8
2Gt0kDRgaSyW984psyyuGymn/WPyb92dQ8SfRlZ6LkFKb06MpXIIAcEUyNGA+7eGsxxb2+jk08Z5
HUYGN2KibjpQZHtCV6b+mwifmqxfftxr0zNEgFgJns+azCChBTVnr7MHg6MODKw2bBimdkePWUf+
fORBftXAw9gwXyyKcD52ZWJqOlTFVQMa5xoCd6WTG//MDFIhTQoezeEP505iGtlzaIDq3MGg1vp6
M4PoM1aSOXIm48eCwT9420IoezAbUsvjxfLb00TImoEPlajCKeP2sF1yy629RMy+ivvUxlH3z15G
OiCzEvEQZaSPCUfzY7huY9/2NJWDMDBbyoHDpSR/ojN25S/COgBiAFxhzvwS7hK3YuiJOnF0vay1
ZnVWL8hoIKmzRo1GVBmOwsYiC/KXytSwOsxE8z0IRaJbXrjWj47gwlFFLDVTNYRfRJ+4at4vKyhu
zWwKlEalLoRoTPWO/MHKxWjoIQlfrjR/nUJeIE5bPWSaqC9oOZD8gm6yJSrGojqvs4xDntW8i+/5
dZUhZ6ubxWMiX0CI4n0sNmPWQV9XqxnAvY7WwY9Q/fcct+9q/XDi7mr+gdqP/FqzZWStJseERwwa
IgcSlPLpAhiyz1gXgZyaJTfrWHzMNV1e9wDQcxR4QPSLAdtRvhcEFZtqSY/aSwpIAY4swPyp53bV
5MOGJDWoZbPt5zGTNScPktVVbwzWlP2QZgovQAl7XlNOBzR0EixYzZ+E2FobtueN0gpCon/R3iR8
YQZOYV4lZzjIyY7JU5/aBJGy7v49kxeMa8loZhI+6NS+zfhdLjqoQN4mPYMQyRSV0A3xYORqRwx6
jmr0LAigcKX47AkXandDTCXZWP+H68FUbW2PvToVR57moyFB9hMZG7rV2cfseBOkLHg1JTgQ9OVH
pbSe+bmtSfC4H9rvqJ+SLtHS2rp3hnPu/sXcZ87ngoNrjPG8jX+Qdn9Bwrh9SxnY7frkRaezC6hH
R/fdHVUKiJgIqq1bJJzDF+u8dPCV4vuYQU0AemafWBBsXEuqNECMvFJC4Bwnxl5ipJl5cZK5eKDM
mf85Trm/x+bnrumD7YSmtHLQWw4Vqa8sRToAE/f29Wyt7dhYXR9P335r3XFZmSXXLDHgIjdFgNEQ
trecl16HTOl66/AZRuH6tJOGCqdnwjj//59dMkOIsFQayx4rOUFrfD7HWA4OViJcgxsdx2UVfJsc
dRQeIkTtZxDqe8oHJ4OoDMiNjQWlCEsJ/awH47eofusFllM6bC9L6yYlszzMFBvQc1JsHf4qXnzr
dsx3SxszlskVpYZIHGlDJTBJPFJJBEQjAbZyBIzXzWfZ6A3dnYrnBga80TlIiYqcS51mHyJL5ZsK
cxcKNHf0FE9k6vAd1d4vmdM50MRAt8i0lQOYnNd7sabXQVCEr1AV6DSk6qXYcudAbBZ5jCUSVUng
sndwe6cBJznMYGPzZMlHsGbXtD2PxQniqhzLWeiSh2Zj7VSjJ00XNfW4sgkrs2s+s5rVWVBtwWCk
FCO63P6zMgvGbZjx7YgKUfrwa9rRANvJu6LfXnQ8pqNmOQpdzcfZauPntl6Sc59m/jOVBXSQoKHv
A9hApiBZ12AXWY2wQvbIXPCs7533DeAoIQAjURN8LLioIgYyhgypDs9x5OBiUeT/q+LsJptAjxWW
yG1mDNmub1xBsG7/Sz/7Q+fU1v/B96C/Ozeva7sBFjzRVehtGjE2UYmhLMLtQhLmHTDFQypZeR6w
R0eHHDG1YfemJkvo45/zP+Iiet+MqUgO9jfVgXOwql1rY4Q+6O5SV9iLMqH6kA4DCzhCEt19qtq2
KELkHN37HOpxqYZvK4avbSprKExlwut3txfxstqvRrhOZ9jBAkESCJtkNy9Hho2xD/v+Y+fY7kfy
7XebqH058ooN6+uC6EgUBT9S0vS390W0XYAp7jJzUB7rBYYXYLXruCkMk1gNzK4F9pq6l2gSTQx+
BiW4AUZ5ZYuVA1E2d45dRwrwfA+LwbOzv551/9v4wvCEE7+qrxWFRELcxT7OasNTgnP3pBSAc2KK
E6G/ELUBVte/f+ewVapfV+KP47G8gIlP2yCMBTrtH/qnJtUKS/3KzLyV30A6MZRNv8bQZ8F940x2
nKuDgSt50buOMhfF15/HkvhrLbuqI24n9Lxct+LmaLlR6J3n7fioyutVPOag/JvXhy7Zfn9dGy4S
Nm2gZTINzJNJ+tWnLdaCMAX0bYpAEkWH5xgAwKpz65YtpWIS4pFnTepxl9kabiypDpxVJBKpbYLa
QuedBXvZvrLsUsPdzuADtoAwZoVy+CetrCsNiaEaJX6eY+zPYUeDOtEIhc9u4fj4w+6twpM+3Oqf
T02igTzwPDc+RxZVNJJfO3S+4b4pzcB8QOzLxmfSMrISLSLPsJ4F4S6zLwoxjLyf78IgyHqjwvNL
OGfSCoOmDRq5IM8AQNLNldkZ0+Q1fH3ll4Mug0fz3IU3t/+zSbA+1ctIlaNt3Hg/3OTVNEEpm2G8
47MmrQUYvXcYRCl5aoQUhOTyiiCHkDZLxkmAVDsI3NzrXGxdFTCsfUVGHArCVIA65/k9SSFLVnvJ
04u+pzrDvvfRuDv30wGaFUMP7asG9uzFWcOXF0gYm53hR2nEHXqpnC6x+C3FNlhXcrb8bOZ8J5+q
E69JzY1fu2HzibDQ3mgMU03Rd7eXAwEKqVA03OXea45RVxb292e63HWKjFkZI2/SqiwrEC99IjTE
eT1O/nMIBFqyrKHogFx2bvKfokKeazxWztns6Wa/1x4fQpdgznUPBgxWB9m0Yah6NLvgkVp187e9
U12AXQ/S0yikc8xfidJqboqS4Nj5hJB61tuEgJJcv69L6SqhFs7dVCzEgeQ5NGfrMdcIwz4QTfMl
2pr+U3TRVRkhgVBqM2ONcHw6GIkEcgOJekMslqJqLtJsM4wAilncQenjma68L6HQY9WWF98HE6PZ
0V3IBeeVS8xOXOv6YIpQpPKpYsefIAih1DZd4OXRnB0HdGMGFVkZ2bsQSukOyKCimvCpagogHqdy
peL52jOSwN+AMU23tYB+ZTnixRgElrh7+lgFGmQ2labu58zJDYhYJ2y88xjP1MR5ycnAD6DJX8LK
ZTmSUlWDu3jnbQRbMC6hjjwjwxBOPUS8XrXGXETCb1xlWQdLPAOnvOc5LHrIaJfDeX4d1x4affZ9
hNKTUKbSstJ+GJLE4F4m2YMR/muNifYaL3CEz1M2M021/py+a/DSHJQh2I1mBSlZFm7BbFrQAiIq
L11L0/UtQEaZuwbGEq1wySJnAYQHozndo68d20cRVoE9NeIzY9+UI3sD0JLFdK140dA4uCUUcKus
z+5dKyR+8KqUMgcnYPTo59yt9Z50RlbpO1NX/tPrpwxlg4lZWlzlZiKd3N0vScME8MR5kKcuG+D2
5qhvJFQaoWYwHyxN8+3ils4Pu4cBFmLYPHHr+lubZIu3UZJGtMbNIkNnn8yuxtBjCJkY97hLcxqR
2JyVsdqRTB80tpeHPTaGKj7L7MN4+kraJHcJ8LxrywTqaq65/o0VNVqua37hRHiY2OybM9Gz2FlF
35QTh2i3L/GgIFIQftexr4dHAjb5aGjW0YDgsxr+Oc4hpjZdq0ZBsgbY/EBnWtfc/iIUoBeqvzoA
mpJWnjpBxkaiBGd909kobK7itI9rL1DEp2x8o8DIm0quT2FZ/GYveF0N85BkwpCxnpYhqNxMonP6
SKRXsVasPnDP3/q96zRt+ekmQCunqyCPlwDVg3+FKcxSwM7zkJnQuisIez43UCMeeR8evPKvWZWC
XNc0O425Z6yiI0IbWrG5Mg/woc5QCNWXbuyFlkvv/QlGX+AC6snvpxCIUcrFmyPxXyWZGZrF0TWf
7UDF0QDyhrDe20vEqB9vzCdYqFoU7x09i4GZzqmOhhjS4Nu0l469aCLtNq/IUp3CJBW6HJSPrFWk
1fPGhSwIOW0EQWBxkfJxCYdCVrEoMUoucXygO5DTKOn4yEwc+S9lxHiXS5St0GMF6/lq8m799JHa
VoMnZevlGgs8DjzW/MhAhEYqZZjHyxUAmZdBEJgFCZji4uSrFLTs2xOZL9JCTnIwifbAKqp9MsuQ
TeLDeyVFdsPTCXFPJhkdPsg7mPMqtrjZIz4jExPetaR0VhKBkD/FPAB4cjX3dfda61utM5aV+PEh
SQI62gNiuu5G8xwd8lqA/xWKFiM52HN4tXvyiKXs5aje47+60lHCzApI10sPB+OnbA7+laI8nn+E
bmt2VwhgGusjGO24ymZYxDGSBQa4c8apNFGBNjMTBVeHxE9Dor8ksmXbLOugePkYhS7ulrbduIge
k4Oe+dE03k+w43+VSTpng/nT+Wft2ZuIHskrlGncbdoTw44PF1aVkHSZF6JNIFkRFZMMwQlGmtyL
US72vE7kOpVTtLjQLUk3zB5DVrA0nKsn+Xrm/m+EII/cIFBdPTF3VlpFArZ3vNKYEMltkvlCSqul
HKfDsBFBzDA6LamtC+IQcv+Cp0QJ7hE1GkCfzReiJ3bHeqZL/Sh68djm6rT2Xl7ilUqCZ1n2v7EJ
KhuigvZ6JffkNRwP/+qWlsgb7LVTI51pVSbZV5eFCXt7KJO0O7w2+HEmZeHE4FtPHBI775bOz3K+
wfuOMEBcHCm+q+lEoVoXmYJQLKKvT68scy1nz9Hlcml0HAcAGih9Hqdsn/Tmsc1qR9xT43CNb0BG
FYz8pVFLAUaRHb6oDok9MIS6RFODxWIg0Oly9XRNCZ8yas/VaFDZvW9R3EX5Pm9dsh6sATCStUfd
8IeWHSIunRY5000b5jFRDA91bLfsmGYiqSW2GxfZrxRq77lcXyItgBEXoLPCGMv5ZlEXBeBih1nk
ELEz16Sjqs9aLtypxSpbUt/krfLERdTUSBHY6ZbiunQisK7woYi4QYbB9oZf3ueAwcYF/EEgcvPr
cAFGWFlRepy/s7REXqkUlhaP5hoKSn7tPPCqh/p3lCPu//lUXIfotGV6R7UkDGd8AGvizHJXvp35
/c2VkNMGXZCS6yyglxtHLEoHIxRKJ4JApV4djZleUMHPurhSlsS+skogAGZYGQhP8NXguPm7Iv1b
jLGrGsfkDULu8Fz8x9Tqt4G/eCYcEGzG4R1Dt3QxNACkHYH/oi7BUBi5+8eajJnCSR2xGBeu5ZJA
+XzyI3etNLTUi/JhYTLaOYOl8m+wDBUhL4lYSyNHZTx57ChuegxlYya4A11lOuKuWEOfzFTDMvzG
VZTQTQ9cxeFluTDWWc5J9csaiZO6VZIPEHY3h7I+LxBM5REUYJfpKCaZnTXK3hFMOQmnn3anjF3j
S+YOGCztYYw3dUsoAOJapGjAIrYWzADd7S/7jMKUWJzHSOBUIBsPB2+txA/kLUGRQBUjP/hpUKZ3
V+om4u1gx+pvLFxUyYCURETCcj2z48i0de+9tCz5dM8qEX9Mc9LAb0JTwakMU26ui+n3NEo2TGCA
UnPX6B5z/oOOQqlbn7tIg41xVSPGG4NcAwIeminI/fGbRBNGsFFNyWtzvt1+EtbrOYyps87OQiqD
qjS1rGcSi4xUzVyVqZVC6lPG8djsSv7cLfLl8BC/GqwNq5xi2kTBNEA3uvDzkmet3m689/fLurwc
E1dQeW3TipL3PnCyuonkBnO+OQoYniSUXsCh/qbkIqPlil5jW0bzKfQHaY0+Dp/VKgEX62BVHpy5
9PJBf5H54tHSDffvIgIqaH4u3CzP/HLV+DvVLUNIiTJxbJOTkW4PPjwuhIwNZv8eo9oaTAfUGlng
bWWQBhOs0pRVgFjVf3Iy+Ppj4zgMyKX8kTrtSLaHo9gI1ltjYgEfnCbf/YjmFCiNIBq31ZfcAb8O
4rHiUzNMS5geQIbap1KRXhHIUwrLc6Mj2YjpEZFKZHc+l4UicfMYT5DAUm1lNjO8jirica5jE/LS
TdLwad9qD/OZv4huD3Ol1AJPMoMJ4MyBOynd0SaI92MSLR3jMzF39mLVvdkWmQyQ8A7zdmnYHbzC
yw+lnUnxHjCpLl7HwKF6mUXbuahuUvG3in5gbW0YERcHkdhszZLXEH7nPsJPTO+xR/I2vjLJs0g6
WIqBLBwrFFtwMMd0ZDjA2AcBtxyIkFYshkjBwXoZXDcvsUxmKgkTM6xy4fVZbjH3L1a6eSKmQAma
MaiRUGInVyHUr7GK6m3KyWh52f2dtAbJqUS9lrHd0N8BS89AlvSA+ydIo8dVuDdnCrKmRiH4ugey
Wx+JwcJHde/2cjtbYYXiaG+bwKGb718s3MtdCaGzcrBdFdejt8VG1FvDzK7axZRjv5PLQIbzrakM
sMJj7exNFL61QWM85bXY4i3XiGEy/UGW6k/tckwi90/BH8nYe1QaUD5zqJryXqPse2Ud82UNFHE7
J6XZd870YgCiRz9VyUpQnm0Y/9NhoqioFP7safBVpO+03qDO7tNx0QPBDgPMh0IdJ5Jel8ruE0N2
H+lEewREDOuoN83Wc3qYpjTEljaOjDzZ2Ge+akTKbBi9EvKr7FMuklaUpjZ7wZTjNuKwEYL9N1Dg
irOsa4JpMZl9VCFChk0G5yULvLJTXuUTxv/bLJxicSX2mbDBbPQeCKbmVlszf/XWHDNcFR2reyU/
nC6WFp3Z/Lazb7Z48/IYHNqwVd5qEZNjVmQ+lcBn12QT3WOZNO4Y5LO6lB2+T/8RwE/q4k3ZcBiq
l3Tj5CHKyui0lSnicq3oxkxt/zAFpJTXi1xCzwgqh+zpq42oVz30/pqRGs4qXVD+FAa6iF1E9cbR
GZdQI/uYa8Nb3vTW9VxM4f+Mi2MxyG+5qq8v9sJ/KcdXnaKhecBKt+Kh6d6DyJFqD8jemHP+l8RZ
Vhgm9Ec3+gxA4Am1Cjh5WIIK9C+dX6o/tYdplzR+lAB9cHj5qhXy5HB8Eq9lEHev5jfZCFjrdGH4
T5lv6FNNo/QnRcjMEcnUCMtcuytDcMLm3NKK3n88zR6WRd/zC5JYxNrjT6ogxCz+N6a3+L1lYOt4
MmkSq3IoQEm2HZn8m0eXeLrxytn/pS7bBfyByN+9fJmyF8xY/uV63cPT+evrY9bcPjfVY6XAJ5t2
vnAAsKGaHq3wtOySczo4R6q23PB8jh6+Dj7LcwIUn2Nqr6blNk0xGUlvmNt/8EQXqKyHytidEDHi
TLOdISvBwNxByvOx84cnP8hBKXDuXiVqsTVlRPJhauCOUFINnwaPQkMD7NjgNHOGSl/LLBt58xzc
lqs4xIOYh5YIsQtFqhp2EeN/XQ4Mx7hEOxmBEHh4O5GdXjLVKDOUharVBW9gT8S+IpEDP8QBAwMz
JqoaFqobbF5qdu6UQ6/wGgC8moqWSJh5qjRcKPPIwZY91kiKUBWFpxOhJpLimDUWYWO45leeqXHe
c6qKmBabV1yHePhgNZfJwkJk1nYvJ18Vek+O3wrJDACmX4Zqy4Tx9CeDEKEZNyXqJ01u7yYeFOPh
R+m5KBV0LTZkEyDyjMqvvFKQn0bzlZ0Ld6HB2nuR36+v6XetQs/sSrEgNmbRUxgWQSGTpFsZ6Oxx
Ep9FSvLDj5RD6BOnqS6GxDCVqp3G5U6wAVfrYikkf2SXORt45lNOhxHIdwNoThqN8+tXN2GG0vcm
MuHul7Dag5D6KrZIJqihpzIiju7c7rQdCiJVQnQ175nQiep6SHmlQcTNFuCjf4acby1W+WS6c0cp
wPg7WK1QL40dlngTxOrU/PlXjmGxAkbQgSG9sMy5544S8uxR/HjUSQ+PMbBaxaW56aiUh1jIqao0
zYhhgKqgYeTxqWv6itOwQFEVFQYI7ofTvBASd+ShchtlfTZjGknQpP3FdhyKhe8lD2MWkfkbY2bI
agYWBKkGdszrKfyk+dsRqDO1ft39Fxm8lhODGkys7S4krJF954fmPgEeCqi3DznJfFUzi0FgTxOK
q5BOOrNN9QLZooF/UkuE+RJrj0+qSUnk+xK51SsRUdCjsipIyHl0imIUQ7aJwrjSVEdKa2FIVdQ9
M31z1qAMjJaOQieKLC6Yqg0YOtlEEPw/pTSNFV2UV5hro+NyEoTQNKdl/yOEYAjpS9wMKj7D2KY4
Z8yUTpe2XMLv0gRKSocrqIV9yOT5tIE9UBz3JJ23UWWeBb3W24KZXeVvLgaTe3MKgYdnQXmhiS/u
n/SW4hD5Uw7Ti7oVD+y+dOpfBJRfo64c+YwLSVEBeSJCSy01HCBnYlgy1ObfNBJz8big5NVVir5f
pa6f2VGW9bA9fS3ulKjS7ajy6CTG72krWLVrHHeL98uI0/Jaocm/uNFqJp5lyhFH2+x/N1rtGcK9
21HyZzF5YmcLcK8XS2SIuLB/b7vyFr5V2qpxWXh/IfrMXxpLISe/pAYroRrPu9OU/kRmr//RaNGu
r4U0EauVtq9xMVc3URSJxbqT0l4k7NobQMenndBdhx1C1v7Rnb/8Pr8BYbcT3o/uYY9GKl2KuY2S
2e/hmEHTFmCeRNbjXaOXuzVwYZuBgEsfRGRCy0We8kWMOvyz3C7+Y53Ws2Wbt1gdNmq+S7eKV1QQ
mj4WDqyD+LL5Q44ywcApWK+yzZ+8GzcHjCjgOcI7RvR7VS0wuGmo4VLFqAvHHINI5hRqZ45vvvAe
Hwzh8slTiGXtYc+GWvKxbDSXN+4qcaSuukFwCc5AZRocHQ1rLySzoVTS+OxeKCcf/Nbzq1vbuimb
g5UwNJlqpP+A/Bb1QUxOSbrUG2ZBkHDzSKdxKMqpKOHX9KFyZVsvJxk6/ddBgGstwQKrGZ6dVxoh
j6paRQctPrx1ffAI6j/jZ+TO1KuywUSKPuJ4w1MYE794TBrIzym+ydOCtOZhaAzr7JUfU6t0OB9+
HIRzFd4iztZPVC6vSDKjediMBPdLr8vrOajgfZng7PayVuBEYJXGQq9qvn9rFzn3go+BYIU5sfz8
b6+yQlJbF83tj/BGMX/F/MmFnzqb8TjvaB2KSVtFTgcbUyeVD2h5RwzuuCOQWyic4Kih8B90jlYg
61wGbG534DcjmrvnVvPxiP8IM/NwaBGz8PxOWrbn6jjTt1M4LIeORiyXPPJ7tCj3d/Ng8LHuSSHh
G1KK5WUxywac0GIyh89C2sRrY5LmBczCxD0WlUR8hdVUreRWxjKr8+qtExPUIEngwPxfhDROrMX8
UNuP58lQIoXgAQZ926pxpJ0CpbUF/T7+t1kG8XxnjXH+IxQH76Ol1LpMwCgjen/XyfNI+TP1y5DH
rlL3ca95XU7Gh6RmSGlb2k6Zv3ncV7VekcU9jAUGiivuQFx9yWQZD+oMYnab+DxyV+I8oXXVAMcX
+Q8UEkKl25Kg7sD99PFvsKRqjlVzDRx4tQ4p164AVfReurK+/t65KGhPb4081DX7B9JTdoCM0QsT
qytxDC/T8rP91tNZCtLGzFqPPATUDfcAUAQJa9zq2tGNTfK5G1yBQsklNSDsouLgr9R/FVL/s1YT
3AqPq4CIJbKKcJzHCdMESd0lrypmT8h+MxQVg7ciIuH+Gj++do4u8X8yW5rc26NlCeYvCYD8QYwC
DXUx9yv6AJnIpp0NjayUT6FBt50POR9f+EE9vrki4oqaObd351EoBtcshsdFAmIKKr60VCR0QAwQ
8yzUJJ/xS+gVSWWisp/pYYaE85sj+74U6c8lWW4yt520wIEh/TpHXW5rOumv10b2UGcXZ0bkcbve
hGSIyFA5gHCRdjKpBJg7VZvgbQgcRyb2b2jmq6geVfZe1nFsc7HyQcUUNYz4DfkLdNloioelHEoe
vBuBfP3+buzyi5I2GoAWjJ4mQDRfg/F+VJJjcdbwNOKHzvHbZEJKIu2V4gjKlIYwrMn6XPmnvWJd
zqe+t2NoNfmSvaqJHmBq5yt6+KepzRBKaZS/9jrIBI2PfjMlTCSYmUNXUJ38J36Jw//xzECFJrRE
pdAXX9uiXtRYx01o8Yo9kT2ZVo641JCZ5NKO3Z8nXLuZI4Od4EE/KYH4wDqtpx/ZhvtpqQSKm2pl
QCIWYaIa/viTXIhcAUbn7x2g0dWMuIGv+F3h7AP+PLCN11/VpbAL/mq8oDjejvPANFTZ998OSVE3
XxxNR6OqyIZf74Z2KL4tbGdl89i+/iLjlnbVuQd485OCfzrXdhiXi51DwnE0MYk90qM7EBkyjL28
w1EzM7rmM3ZfAoPASxkcmT1UfqqQ6+FGhNnV2Mv4I/qprK+5ZRpXG4r1mWuQvRq28WPVzO/vJ6+C
hWy7UB4PFFYcF1bcG3orGBZa5hhAMvSburuSPCC1EdgiYhxeG+j2e8gDFNEoomqNhQgp98yAjoes
vVXyNq3Cigt2oO8jmIzUNtNFNvcAGcsTItYGkEKmbTXPMBAx8dWEm1plJrOnv6aKEAoo1qgYH3Mn
wwTAvs3mQh/O4WL7txD4BcN4ydhAfmugncssUT+o9kujXihaScuRiTkgznQIesMLId+OAtFZ9yUQ
PnUf9gvrJgWlcj6+7YpnpnqF7U/BHoFyB0bOZhKCDt7GfQdm8JRxLoPICMzfkljoVyzejifYfu59
GMxyr42+KtNvB0vOqM2z+OkBbGk+0GK8PD4IpfJ0QTeW11UfN78qqWiu1L4CH6ooRvKY9uJ6phW2
kYx4ZHNDb7DMzI+JGyuWDNkxJIh42Y5vScAysKnrsIUblLezn1pHPmchGz2qjSUXTsjF7W7WAkou
l0tdpAKSm9/K80h1jXc86g7FijvG4JJXofV/G/PdaqarVyXaZ2FeUHWJREHmHrfNy0FCXj3Mxc9l
g8tEAwlfFIqzmook7jDtpQMKczXZ0Z7oGYKLnQ63eMSfLuzgvb/JpRJ9bTbEbvUuNmTNB12/mlee
+t5gzZeJYJ+NYfi3lmGCwWv3HP7Pe8rhbHE6IfGoDBPrMqOoavSsuvvuj4ZvW0bsVJd4Ia0OBPTF
Y3RvAGuTbR47KVrFJUUyIh6oY3Mvf2rnI+JenX9hvkgyo8IC4Q/+fqV5p7XvNtYnsp/8Gc+RBEKo
vF2Zj/Cdlv+D5F4YWW4g2cyhIjEu+hFK5tyH6nMMKuxM6+Pk2X/+QYCZiyGumjV/lTxnc17vbKv7
4bi07j4LU2BP6yoNxXLLR1RnE/ZHDhBhDYvHVp/xNgL89rXKuBzKi0vsCsgpW7EkobcYAU30+18r
TrpqXlUIgJ6eTKWSVp6vNFZ11YnTJeMabTd7mSra167gDtrMLGz5F905TZwDojEuDYyWRyj1xTPQ
lMafv+z6pi6RyT0NfKsIdDJCX1EqlLf+FVrTDcD5wrzSr7JOhT9x6jXr5GPw1bPAdagBaIQx8j/B
gLT1X0XgRpUFnroLeNJbKPj3eXv9YkqrGT1ohwVvC/ehadXNvRnllrFNneYW2medbRf027+X3407
bugqGClcXCCjOpYso3G699py/fHGEj2Rah3ywivbGOHs16IL8QvvYLygp/wrWpWeYadaYfzQTjG5
csfQX2UwGUBRJV9nkJNMUv+DLH+20Twzyck4TWOV9UUSGqjae1H3q9vfPLTYY6/MbA2lF0/OOJQU
dYVViOeDRgYei0mlGoi2uAzLBvDS7Jos971bwtIrDd5P0Hdcozszn/mb33i5HagQXC3t3woUiZHd
ljK6huA7ajVb/OI6RD2Prf7TZ2WYOiVoDQFKvSCtWBH292IPUtLeHDPu1S+DV9hu3kWVhp6/8E9n
1Aft3WLfvxHc1CMgSiZQuE1kMfi7fpR2DImP8n6oJtjVWGnpGRBpYp05MGpkVVBmnp7i3NkYbHIw
iWIdQK5sQKZzcJqfuNEYXDvggQ+zyIVUgxkI5b7hexPro+uYXKWhejEC/25FBjelZKSgC97LqG9k
zDV19kyVh+ptkwRSii04phQs6KgL8r7jPpYcQ3MSOurMVNaR2GyvnNKaTN1k+PkLimlJ94v0gK0i
fhxxqT2zTxT9CEezL3uiw2Y0n5JObJb1JVStQIFSHKxaZ9avX6G4ruATLkFabq1zZ4/E3yO+f1EI
PFCo7I9pFuTe/WY6Xp1m9G909rPgKwxIFAsU2Pl3IaoBhLuGh0h6UsPaHbSk1lC5Xh7sMFkuUs6M
VrKKmB3LtyaYntgFT5gIRNP1sPSK1+mvfbiAvLttCbWhbOoJlpr8gKH6IGL2l2cfTAYwRyjralm2
DRrxvnFHoxMFY1GcQUAuoEPlrUuvREgAHYHonZH0zD1dXd1gUHzJGxp7CJfZkcUDVL4LTaZAiFLQ
kAz25N2nZzyl8/v8uUl5kWnUcaTl4wbnI7D6Ep/8JTTnE8WwNkt9HLMAjbHZrgUasajG73oqba4M
A+AEyJRfF/AFrxQd0uYvzzFWT26J3/w0QqEH3U/StVeW74MFUybYiS3mhPeJ1yBdoUzdIiobSuR8
p4V5x3jmwqJ7zEzOvFib/cIJn45SMnMpWeoMd25ZqGqJ6lZYpza14Y7d9ESP+tHdwPce2A+vgpeo
fGRWX9NLxgVkSKiQEl2MfFU9lwsg5LoLabpdk76wWyEG/es8lg19UNnMVvMDpZt4EeNiu9p+M2X7
55jgofP5eQDFfntE4o5BQ6d8YzGDkL9c17UWriys4ZjdUpajjVnmc/eqEyCOKCvf48qV2Git3I58
La2Ml5bqdH6uccHUdDJAzb1S4arcWe0rGeLwarVmFXacAqIPjqd/+pIjsCzlrY0DdXlrDmLHNCOS
/4v5j/6UXGpmQnBsVfzRQRP60yjLThGaF5PR/Y/szAVeXkr+F/+0yD3fp7fgTYzRLCLPbjA+gt9K
2eOPKYOoCCvk7jNpcR2k376U6vEkXPyeRxAPfS9mEoztHKHLPcDZ4Zsa6qDxOOQJjGaKd8cvotSu
3AMCbgcUdKuy9k16kgus13NtAh1LG0nQIZ81MapZ/FTwvnE7mWhHscD5ptlhaOJSknlc3+UTs6V+
y7QYsoZsIPUGRyN+Pf6fH1ccrJhp2x9DcbEEU77Z6ohT/JKlmlq6I57wznRGwdqc7jnufA/bWpha
d5H4xcueMtlUP2rldor4od5t2XVfhSdy+qMlUuXPMAfnqZpLStVeGFSh+mo1JkGxh2q7w6yk+3ts
lBBVs072fawJ1UGDUSb95JiBUazbEZCwnyw3XmEBTOnjCHUvf3ZMppZEYCrbFwYaqvaNoKrcZv3b
8HySqkqgrYvfReaFn+ceLsS9C73GHd6NUpYc2hUodUHvhsskZ3HWsKx8Gz2RMF8z7F32tcZsEIoS
LnLp8gYiSoAgtXcIxtI0DyUwaJzxXE9I9BKVn8qr4rT62SzkzPQNT9o/oQqk2MHly97H5cCgSdvQ
LRIvbqF+38dWAhVdX/YzxltT3lFDgyrtRHIQSlUNeJt1EKVQryPgUK8SDYYkcD8tSxz5BFmEZyqQ
MEvkv9NbjJAZtRHTNebPp8gL/PBUP5kRc4bjyhOmUrxgBmgMyTsOTmiNZcs3EETQfdrarygxusTW
e2s55Tg6shNB4JDEjDJFLs9YiBHW+suojX4YI0t/EYzQ1wi5h7kdpp+K5BR0M95zKsthwhuyN4o9
txNh+3f/Go6CkOh4i6Kf+62ycJERhG4Nn0y+3jxgeyvuOnxUC+5Lf4jun7rRi4UXkg4o19vGIIpA
OmGKRak5c37hITmd0bdAL6IRBLxhgUBCqkugRVoV5MSr56gjw4AYZqSG57P9G/QuruJX7sf2+G7I
VbX6X6A2+hyLithitSLM1nOgxYQsN2K+ak3KjDlwYE+iIRFr/cjDnoLWtos/nSMxWLYvyVxLHscc
V9IFItrK84/kitnkQzRnhK5I6kUx3EAmtICqWBZggKSBMRbIPqiHamELU0RQp0JkQzIV3+1Bk31J
l6kdyc3ZadpmTb9B48CQWAqkMV/H3njN39dWDVqSM3t/NKx8P3iLGR5NJQ2fmLKdUXbkA7JxSow8
+9ZXO4CVE1WY4xtA1IilqKVI+5v/jX6+G3pP2ooXSI1wWrlpdfKymZ20Vrf1CapkEWdlFBI8dSpA
DrW0SvIvNHvZ5QtA6Bo95FWeu+uApveydzT9voDXlY7MOjsLTZMUdVAk+dTdV/5QP4GBtvwj+0/s
wHyzMyq2EmZt/Ky/L+SaIizQF1tDsUeSYZbKxBUPeBbCU1pprAK4U/5On1XvapycDTROBlIqww2D
i9llJANqJ17lwhCM2rNvKrZlC8XCO9O9y+zG0fy8wK21NkB30KV01cOLqfaCRRTPfGZbdvnzfzJk
Eui0cjUiYY0tXVFgT66ZXVnbzLizMNaZ8rqqUH6mJnpgcgs2BIn+b4VEJgNIQ0/IVBhWpzZN1bhR
GX8w8seyGEzwnAkZ+4+7OBnncF98oq2T/4uDWBpxbZDQgTXfrDMzHISbtbGiPGnD1qurHeu+dfin
GE+qUE9sG4EGmMYHo7AHaVMjgFGeSigSutfoyjjAyTBLs7LQU+hSBVmoSZgd9cYXgljOJirVI3P7
VHRRgnYWz+L6wXDURJtTmlbtoYY9mBKDmnve/lxOU5ryMm5KpSkbEnjfgVLNEa1TVuEJmQ+UEHjY
DsskhxpcDVycovqKNfP9Rtin9HIf+0WOsMpdUTImudiq8WYD0Hvbdxj5I1ab8RPGUHgjnMd0tUgC
250wjxMzUpRcJI+sGefulGA50RQiPFU+Tf6Bj4d0nZO0oedfgJgb7eUYfpVCHpA73e6gWcOAarQy
ZHADza/KQUy7zn5QSWi8xHaGarzPgBwoVUkj79hUFyW7F28rS13AjZ3CC4R+AtTBIU6L8Iq/1z5t
24C/5KdFnW/NeGZeNtAiOxZseZ1wXQ1nR4vfGAaqATZKvLHX7QjZVxpnVZgOGXAMyCGL4wIrCA6Y
NECeSEyn5sBAho2EljX7/eGESzAS0YSiTWEfbgmUc7GT8tlJh7q+h7TRfvcKEmpo1Djsnq612I+s
BeBccJZU+eMZaPEBdVJhDp2TxRMShh6MCpe8Rsm5B2ewCt9tpOv5IWimMQx9VxADGYUhTgmgosd8
HdZaZRvArHRzFRPV7ZMHsVCzmAhlD+312uNPlgSA9S7ymmaVnoBZ/wOiipKfVe1yfSMq9FC1Mgvq
KiQkHa7ARdgrgstL72NIarjtWrbBQprBUDqtRqZrbSSiZSrJs8J0yyBhL2E2q5srlZl2J4nDWYAZ
ienXaKUVnNfefCjkAVLaVnMZEdY6HN3HEmTQpWDtQRYYqbnjgh5EW4YQSBhLGK9GVabpQv8FPcyZ
lzyzDeb8ODMkb6LTMAI3ya0/dqpe4hoElCXBDOcoLK063YHEzLFOnuJ44h4WhuRoUZ1ZWLV0Vgtk
1dV1pDJgphFBEhaGioI176pk/bGjdcnfJ4uqclYf7dp+/f34LRl6ReHY72RBrH43WrDQMYRe0BJO
CRWv4iR8DezeOnEhac5twSDHqOu8c0BIZDsTRIKkV+liHNosUvcmlZuLjsmM0fnTsAmPSOrj9U/S
HGUx6ivGKTLUsFTgIkBnelRnGibp4NoXHp9bhMiBmA3WpvF/tRXuLsAb3y7nlb/w1zX8mghpoioc
PY1CmcmgHud6NFGdWZkK+WzENd/Bq69DpnffZnV5mJDjVxKnw7ry50XgyGmvcXjaLww82sgesdrf
REjG0KGLO0SjxcJPnlgGjYvm6HCQAaiNIY4FdeZA7thHmNa7+j7Y/aPdoBDkg8D+VfLIzx0vsAnS
m4RnzQLMkrFmjHImUHWaNM+EyOscopPQmovl7Qjo8kqOx+zZbuuG4FNQLcWnZ82r7x2T0OlnWfTz
Md+B9WixbhVxknJkLzWI0xOxF4mKbv0qWpUn2mUh5vwnx6lSJUryGIkXGGXI4lShA85nNhouKr//
039RpSPGbcH14/vdHgrs5V2Jy6IRUhjXSZM0DGwHcMrNiMVMUHHd/0QBKRu58EEzSVRMcAGG1xQh
37Uxl8lDrERuCEHs4wuHjiafofjU9WkBe452QZ9qspmZwNODMxE+7jPTk48ZjiZDBzDTOa20D9+7
u/6amvlrtUy3s34s9m2KRd00U0lcbzA52RlUmaFS5OcOrgx+hiyL08hGBrIvsbT80upLwk4OI/ls
894sqtx51sxOA6C8a2ODXXQhU7klBlvTbE2H00NYWl5h/RqTKzJzkyEq5rwRfqCNKKUWLA8QN/KT
zQGinuzgSSET9HvmdHpxb1XrlsFSqGWHzbwow2+crTG8ArQnlhb42dlIi6oq1aqHqZUf5B/aMwD2
mSLNuH+8ABKjEis2k/9XIQltBPxz014QqiqoGQtFGJJddwVb0o6XGAsypIv415CwQb/WP4prJXEG
6gzCRJZYmq3tlyEERgjTUxI1W7SkYW2BOKHhCBPoIGYWLNZnqQtMs4n7O9euCQ4dffSCpWivR5iB
WIUb4yWUYZYaHWoTC1fAr4Lvl6NgaJbL7n6/bSCRBPHsv/ziCzJzUxATBVIEITwXky2d7ez3fb3k
6HCG0qvXLDje8gUIc2avVo389YpeIFOsHx99f0KvY3P3eSy0GlTzts4BqhDY47SnUhFYt9Qwu+EL
nK6uT54GnLZHemgmnocBnKA0bauNPSWDNaexC5RV8NHhGV45rUCJZ7EN0CqwI4Ai5A+8lBP8OdSW
2PA61pVwpn7MT57u2OlqequDyDKkJmn4GMC0S8vshr1/U3atI9sYlU2lSFZx+YnJ3fpU7S3Zh8rz
6bZ+S774q1Jne95hhSBOtVuWw4lNYKoUVEaP6fZJAWXMvbew5LZUK0tU9VK8QVaI+tRNi7POLjeC
bWcNd5eO6Lt3++BF5r0UxLz4XZ/YmyRiN3k71RhdgFHk5rbEfncjrkxY8IB3kj1wWWC6mbJ8eUW6
2nMAJe0bugaouHW9+yey/9jDk2S+oBcKUHruQm3LhYMxDq8XX/b4rN1PZ1KtP7hLLelzJrvTHbKx
YnuT85kZvI9MFipJLuDvp+z9ENogLe2ynI9pXlKNBe6FEr1t9IKqs3172OcYNHMDnRCaiI/yGQ7+
QHoTRfBfq1Mfze8VFbI3vlS7v7aZnB8m8UJvuLf44hYOSa7GhJ3mAoGWVuINiZFfj83512Is1h/B
2eAzOYJkorrH9PbQpMrudd1Ckek1Sdk2c+rndc6deQfJyKe/LZ7x4S9xjeb/NnRI39mh6BPxKwVO
LAZs6Gfu1Rx7ublrbqPK44Vmh+C0k6JvDhBslpoBB3AkY50FSSay1m25hJeS5oF7262pUkq/2an3
MIq8QMUExhHN2H1nSgdgIA7+gGSy0Yn7QHy0gDvm0w1EDKVh+vVju/f+Re+tO2CZkeTNbF6UcjMn
YGsDeGEVkLf4dActPBlnIKUy379yqA7+BK8M7Va9F0l8rKl5yVhFrkgevB0zi5S9Iyq8CN/wrRiz
FWjc2KS64xlhROXal0/NFuRhEIyXubNsyjIrVM1hvJgWhhB90hSlh7nXWLJwnebKO0WO8UqxtSrh
waIXL7F1l/Im1QVMZRmj4b5d9wkUZzrAfgHpCoMk3Ca7KTnNSkcajScYa79j3Pfv5kQ6Sojyi9MQ
kpXsgkhdsV9AdYC3awTq+96K5y6HmQpa5jt1FfW9hd9vVY9RQsc9Ag0htzv6kOc1Rp7n6NPCvD+l
P7K/qK92rEmyn5gZ/mQhhAs/H9WxlAgN7tH8kasWH3OrOtvbwChBqkC2dT7zdz5l5CAjXtWYJ2zL
L1oShjzs0DRxe6WwiQydeTOqfTC065Yt5tFsjAV7ompZf/DowpaXkZuIqMwDD1PtrMPid8YRg6L4
nKQ4W+UALbyvtnOJxgn6hcUzBdUxG7Ur8loP4lpI+vgNMEGsz/ucXlBC7HAlfoxjdJLlFrJro/kB
uECm3t5G2uUx0pBfpkxlheRgXOkqUgAtJqAfzvdJ1zBYHqcVMCuuuVZbKAbG3rdl999OGyxfHQWs
jSdo63Z4iwnZbnudMh4Tht99vcyeYdaldVK0ewRMEkQgSmI3TiudgN8Xq6d3+gZCtPvUFpV5IEaK
6pOhBey5rfXJSsdtPjaaCMbiXvcZdOl6tMxHbjTNfQiGtrC6T+UX2zgV69nzwMBx+x0oxtwyBXuH
CVOjuCUyrlr/zKFsKqsfd6PZ4iXmp1tNCXvhenLnMAbhNckwJ11Y9GstEIuxuV65Y4Zpvz15wJEB
/J01xLdF9ua4/963LY5rXpb7Th4deWHEN4KO1LH6iB2rS5Fz8Wca53igoh2osLvo3DisyyFi/2iZ
aJ+HkiYRrKf3cjpC4qdNmNaW72+kMol2XYEoVk0PoKuNItog1IqwOP8fp8xOV4Gbi8rMqSEXiNZD
Y+12Tqefck0ujqYKvpV8l9iUXL3xeONFDyYzAgUI0MMrFGQavVsEG659ST4C0yTqVbLe7CXhAqqU
n2eAnUYrpQT6vyy/DZ3RpmC3DfIo+Jw9WJGHXk3CDhw2x6qLvfrhfSXFQPRja4E/LmPkWeuFDJW4
6fBltZmqNUhBOdCqP/aT1d9MI3x3U5jAmY7H/GXq071RHej+0NJdDNNH1SsyLtR60XK1yOugOWVU
yF9bDJRbHQuZr7OGDuzaCPxmsHjReCL3y13a2OahuPk/yTB3jmfvNZg0GYrud5DplKPEcwpJkwWl
FqN+Sk93aPmvY3uHoKvZ63QUDgQNxydLwnExqeG04n8Y9sXGnbXHx5rxu3KERADY/9zTg+wsA8SR
ihzOJlMmKK47QjzQJtOZDwn2mJiVU1mqce6BPqSFvxCLklfcjSAdb26xbR90DwouQiWqCgY8qyGC
TxYx1mdelwhmK9FcVadtq7tf3OmpUWdFuBe4qjj3e5U1c5B46Jj5632Q7ooZmIVBRndTQ+6+V5JP
oBHwdFzSlFDztNjVgeHNDDD8Mf/NOUc9CXpWCXVAIovaBG/WxNwQKBtp4p2F1YHELGfN1NZnF7Un
ErvtkwrYBXHgGl8OG62Fxjgp/aP9SBwyQpsBd4X7qauF0b8odPbcY2HtMkyrUg/0aYAmuylT3Nbv
t01q58rhN9MAMBnorgbKiYGUFY2s8GKIyQzsPXPiXSgT9s5NYa3DigaGUPzxfpX8jvITO2y+7xF3
+zo4KK2zjO/zwv6qWuif52Q/z0FIz/SI6OlVvisZZCv5Drk6YHDMCrZZqYGCHNtfIFsSyADuQTXJ
q1cph/jjYo3HYJnI5YXp77+MH6sKFqxN5mkYqtDSxSon3EYfowtHOGXwXpxCgOKTmdA2B8PV9uDP
vSIAJj0QPbRQQnuK4XKhu5upXrv+P/UFkdN/gGsiFry6U+zicvdBd3KmKjFgWPNBHfFLKwFJMR9M
Htmhj60XRonA/h4oL47sPD7dZOOX7TXuja3vU+UIIexg2ZKGzIR6HGafxcDkFLvXZZjOO3Bt0Leg
2YFd2NknfFBaCY2NDwu1PmWcahll8bmp+VCupDGibTngtZ0g6l5rWJW8ZuI8dBqBi46UzQRl5evs
2KvOQXWQgPIYlFalJa98F61JVM/LDOrbe0eokB4TPL8yeUlZu/hbJJAkcj1WcXbTTIgFtHEhrfGB
Rm1wl+Dhv6Y494iFA9NBV8zrhsX0b0NIGKdYvS4QDOCvehl7apdXTx9cX30+lXSrRabOs6oDjjf6
nKdDYSB4iUtMWmDrTqzRVEJt48lft0d8EukhF6m133EJYJowa1j6Mh0hOsO2N+tPmh92SL7nnRr8
82ebEv8hav/nu0ds/j2GFC5yqJZN0vl1Rl4r0YlXYorpJ3NbVB9Dpos3Qi/IEWrTnKNsaRllGhJG
Jwpr9CPYAjdQ7w6NewiQmP01gMXEO4WaXznn4gLt1/y2bgPcNylaY7n1bfESUsGoNk+YeNhApxgi
/1gAy0ewSGuH1YYJcahUGRzqPY9UU5a85VnEz6I1KGACA4klikFCgjCa0VFpxV2hq6ncu70818pv
FIctJGcIxvGFDW0p22fc8aMys1yXB/+GCf8cdz433onrNyp5ydp4cP2RsUyXQU90UovaX1SKvull
YHcvaE0SsJ2+uSge5z4/AX3a7a2lsyTg26jmIpHWVr9N9q4hFhPabhRh+dL0mE6xVPQ3XFk/Y9Td
XTUAKxvFVSmRmEyNqIqIiLndi2tNeJ9D9oNHGJuCCwl61pJDdf3s9/0adqX+DipJiXiEpBur1IFn
LNhSVKXi0KaV+ec8e5Q5TYKntsyiXmwRXN16clUGspCh53F8fm3ruld8i9psb/QGShvlRWP+9H0i
0mmII9904CUvogDG15cW224KXkqAWIVx7VaIrR1BEEOWOVYxuqjktv2lfvYiSpoHRmxgJspMC7tN
egx5N2tUaruAhmGTitAEITLzeYJk5ldppPLU5a3hwAN4U6dKHBrcdpPmYmbMSvwUa6mBsOHFuxrK
zdjK3owY0RLCKXoY/TJ/x2V2HGWYvhTqcuW/PlgykZUHgodsI7RuozHzuk2jK+3c6sr89K6AjYBq
orBZ4tcAUsnM3EPLsjFgkftbHyI02V+S/JB1LuPvmIj7KiaitgZ2F7VSpUl/IC+YKnemZNf7Q+3t
S0MWnwzIsFtdtBte4bPk03y4Io0PLj0bw73UvL8wuPRnQwNChgHNxEX3v8qY74o0hMev2I+EhYSk
++LYY6YRmM80a8IZwNvzQ8lVnY2qvvvwewst7tqMdOjYjEZ7GZzd1lJh6qe55+2eF3qcrrAX0EUh
2YZS+DneF6igerxNz+urA1PfH0k1YgVsxgWaFPmfkVeZoSfCK68SSYK4pv8IpREAyIpZ/mUMwu0L
wv0eDD/HsCw5fEIheYSU/IZT0vU7k8wjiQSzeUoi+uSOkUXxGVXh3gq5Q8igdi/HSqo3F7P8aljM
z6NtBpEGCovFlsN14fGXJwaxiFbmB73jCd8mlMvGgE3OQtcc6btKOvBaqI6ehg6bZBGRtZ+tlYKL
Lifa/LxqWtNyX/FeX386fDvg4SCpCs1TmTxV86mSXSs7+EMuiiSbIEReXR/FTNxvMc7aK7EdmARc
mySaHoAUpf+HS4yh1I97kaizs1GTVUgIg2EIrOEfOPTaTJ/+WXtKPb/kHmGzC1yzmZuZTU9sOloC
YXTpWGaxpioLpY53PHYRulAZnewSNQMvo4MtmX8PtVVUoNjuDAApwp2qaLNG0SCUlg5BwfnWxVpE
C23Yoe0ae15tf1VI+ejccxUaDo27sy5UyVRSHV79izEegCDIhhA2hgH6F8Bo+ur0gm4GnUfuMSX0
BbfuIMYOHp9SDrE0i4+A04S+jHRRFrpkH4iPQMGanMBiWfOx/UyPAmgh2mVSHNzaL+Fxus+SWgRX
0p2N0skBWdGqCJi9HjvovdYFw5zAEK13tYt9kdXzQd9DTc670XQQrU3A1hfflPC1qxdvRPsoaNA8
gD/gQ8eBNuhu8B5YlnQVFzyFVcau4m7RIrbaOfOuKrIrHjm/hp/09eHDTiYcM+6JGRqk+g4ww1+N
DwnFIGuc/2uQNBG4iYfAceV4dhtlrh3LdS0TYO78155Z+V0bMH0qqgOCyYR++v9msRuUm/hGMb9z
cRnoHqJ7YkV/smHfF1P0x0Czbk1B45AmiEh8xBZ5US1vGo0jUBDFO0L8lgAHWPHKjo5U0rbrIlNM
pUgxC1Lcz9v9Rtytcjj3qUh7hl80QTl33Zvyx+kqsLdoSSRuQsEAR9CAuHYMJFAhDAAJxpgPIGqb
lQj49X7i4cXqiuaY2uTLhlxamPr0PX/GZ7UhYHw3v0HBpuX8d3WnW3Q7VrumLRJdO3Q4JosTJq9w
2qhujmssQ+XqO86PtVVkN3ddPa3aDVx3GTnzZvxhP3QI//YXO/XKanxmNHrLlo2ZoLSfnWNEOU+N
lpWrK8FRsYg7NCe4W/sILYjFnIxkyng1eOgZgik5L7hodoqfITHNVQED6uEyQ5RQ+ugZqt/OjdQb
VIWoPF1k9S3DQo8aG9dO1Z5g5C1Qiu9unsayCK5l/2SL5DseFMlJA9aOgELkhm4zwVPvEVtT59+T
NKjQmag4USShLVOVKfS6Cp42bgswdiTMdHPRayss3yuYm2tkgbqbv+MTCI2gqGAQJpBrDiTti9E2
H2WVu+KYtpKiedTh291WwCydKWzKgYK+ZKSkOKFgGPEFjnc1UdLH7GWbz3y6ill5VwvAuekJhKmi
uIGk+PcT5g57F4ZSbDvqWC0ZvSFPgOz233rBhmWSMM6D2gWeoy2BQMFG59rSW0RI33uJVrQ9TS/K
gQe5pBingZyR+4ghlZVNEdZCIsHVlJZH0FoNsheVKOx96ArYUZroBipSTtq1ZLCAxKLrwzlyqKyD
G2KD+YdeUkGCfuvzJNJQ1PASMzbRZXrj5Ub8qvir9Xg1HYYTOC0cq5JzHHq80R5QoaHC7c/4q+FD
3KkW6/KsSmVWdTYdoH4ZYdrqiZIBMtAFiCVt0jiT0cIQro0ybuxg3iaQX1Vw0veJTGAylAnXViJx
70xK4Onk9R/Fs/4DXhOJ45K+GHBfagX2tZDeuViro3Sms/vqaZoSZQHq4ZvGvg6OVmZzdy65NS1J
c8c1XX4gezEIuSKkakm7G27A2v1ez+7+lQG6guioodrAd+oeTVisIzopEBM35bGy5OjEGnYpZdNK
TMqTHuWvPMaDB8qM0CP411vLWQ+s6xyRMOGYHy6DBeW+CKsGLhwKh5p61HkZcxP1UuM/t8wtPfmJ
m8s8Mr2vx7l6prgzADlfg+MdiY9G+FVdb/vG+S5xpuwibaWqIoPcW9Md57K2xbCqvyShZ6ZNORMP
UvaCfTyjNZcaiQYLMN7boicxgIZVaSc+o9C2OTzRd3UFm+KNHYOXiXgYQb0x73utKC7MZz5H7f9j
fZIucmYp1MkmhM2UQHzzIVpwebFFOJ2cDSSPYo8CdP4wYAAG8KHozOi3V19+gip5pNR15b+ue78K
fObA+hZKTYHR1ioGSayLsNv6g1I3saLGjWbGLQTN7AZFIPNBpmYNuV3VxxK80gt3YkxXVjQXok4C
CGEKewlehhKV09TnztbOdJlMWfo5Vt4bN+TWEzVy6mncl4wWadcRqSqv2Aoa2pcfApqmFkQsuGu8
+6CH9K86jwQkli1Vo//XmecvSeZ+CWEbyT6cxK0MzXKlGHEYaOK/dfMMIgCSvCFfEB9+bKCV/xOR
PQy10kKw9dWJGWTmyAzeLHptvAcWHB3KdLAcBwxCPKvMEoywEgaYcRadW31aVf7Cx75yAOs3gGqt
f9NNGAV+8+xWLtuAc3AG4qY/5PTVrh6hHL5DpZrTHnCluUx3LZJ8W9WNYrFvwQ/NvP7LS8Xai0vA
sdFOuZM2B8NM5uyDCylcejxz0J/CjcAySPnd1SgDUgnEvxFhk9S7f9cSedhBN1LTOWE/Uani3VuS
qzj3rEo1tSJMCtCU3ioPjXyrpDeGzFdz5pW5R3fgb+Japf/vygT3KXDTbKhIe2/oPYDWuELlq6b5
3gH5LCSUj6utN+1VOnIOz7lpUPgxWkCPwZyzqDjOEQl3qkqcgb+ASpexUndyNCVoaayZH/qW2njO
yNT8B8i82XwCF4zPDSNL0N+64qx57knZViH3yGyfx0cOyWkiwfRMyXVEZlp+IIzfyZdvvNm2pcDR
W9eIgLrphlCe7b700n0KXYgDSBRaURx+SAp7ZvtYD18k0srIxUrBWEQ+DQ6SMO/fSELIdaGxW0kl
3GAiwRSDLK5XYCw+KhQ4h2AevORnfHzJJ7iUel2nssN71HDVz4UZOlkkUWCLbGggiUbM66fYQ7Ri
4u19n49sFhRjPp8fjUuxtmdT9xtU2C4ip8GTflboZ/2NFYMLI0Dm+IqzBnA6weds1yQ2APHJ3F30
glM7ensj2sPXSXnemHMEOgP/6BVd7cZ09V9jrzv3QkH0LatgQ3GFLv3MhPVrA9hd4jEkg2UKr8WO
kTrkj6k2xMIUBBohR1CXuDcdlFXr3PgtL3rqAo56XtI0OytqisMfXg4thLVgFw9BP9VRssxiakxU
anp381Sx4rSgHeElfz8FEt/+HrTds3afshgFRszDdMRay7sh6gl+/QIDFEfJDl3EoioVV+s1Orf0
bqlakF8m2o0AdWRrEpoITzZikNAo1dbJPINF4BhKpi6q9KmqSsuvhhFkQMoCKKyPY6Jy+/py51Aq
dZqJGoJ11Qj4+L6tGRN3y90SrKVqcS/t/l4iCKkXl/F6qwaVHaxZ6+bEhXxjK2wrZfMH1NWLnrPo
j0XE9HKUGtKSI458mJb31jfS1wKzm966zJf0ouxzyoZOs+NFwVBawRimHrzBNbkBF8QK392iMHiG
z1xnUgGCEtZKm0GOcCNSx7kMRz4PVfSr5ZM3NkADFFSuMgng5tOGbeH2DAvAM72aDBWqSw/wVhTN
s2HCACj9HBCAqhN7isrdK3Fcin8F5RsIkZZo5/COs4tcfp0ShRbTsMuiCN77pmiaqhJDyBCOGHKe
QgBLFh7DEIwqQRhsUE0e5O3PYZtW52HvGTXM7eYySi0AKd8r/YSslVoa/dn2vWy8VQMtgK7cQN7F
Qi0ZFNjjcbQx5O+dLIrWJKEWpaEbx92TW3dRzr45q5NVi6c5pw6ThYCjxFMu31Px0MKuDwaF7fZ8
MmmoBxxb00S8aV0mODDokFConx71YtceGEdzbjK3QlmwkRr1SfpD4EZ1HrVsfM6/lHAjoAtu3/Pv
J1nOy4IwbQrX49EeFj3jQVxp7+Scy9hZf7+hieRDYATy43/YOitFEUPtY9SQgn0RmXA46rp5AIZR
ES6PB0xEvJTuGOcd1l579jiQmPKJkildhk0iN7XJ+ADWuvPKt0L8qlpvEoFx4XeXQMCU4jx7Brir
u1+1jGr6Zk+LfmHzgqcnEzS0JSj9NYqK87wHVu6Cols3Hsx4B/rhO3kHfjsJF6UIMUiq1N6x+ncW
RgueA72iULUjm1Rdn2jbC9jF0C38ORQ8maON0JfphblLNzosapzZjtvnK5hYio8VVL8wKaapHjcw
6H95d9OLz6TRVB1eIRkRZ/12Gd2tHBbcbxyjCWFJ1U8/LkrnVfFP/pQD2xZoGCaJBrFXKEFCtBxf
tsaDTFBvKoTKkW2msUVQMWvKktBjsfD17ckwTAw7k88mQfkBaczJ10SLwAZsAgaL+fJirzneEyAN
nYmU9nePEdkWbnyZwB4N0+vCyO+z8Hih5H0YC84FTo7ubNU/Y9iCgdQgDKZFNQN3SsoIdm3x1//H
6rqrKVKoFjulfkLPhANpou+gV2sVHgC2Ct4+lHvzU42cMCdb0EsxB6WBdbOZN3E3rdw2xU/mo5+E
iOaKUkRkRWOZNtxhaH/SYnuQYdcjzpNrvqJztAvR5jxIN4Gy1Roan/J/opz6uJtgHazZpY+Z0ETQ
wuqMGZGa5eDH8XFetNUtj8gUcIC+RKzNZjYuuwyReCt+53g21fiJP92ORZVrubzl/L45VmMBB+J7
XBzPVDpYTRsJ3FQ+ds1vPqjz6PJjQFKaEoUTTQ9iHYinp8vKX8GF0j13CQF66Mi7waaduVUssEs3
gVg5cRQbK82442JAfXBWEl6l0t0GIXyva+8IjEStTR93D/TbnhAsB4TEuNSzG4zI+MeywOXfzsAf
g9ZRRAhE/ef0EgI9+0uYZfcLRkDtZ4Zxe8LjU32BOOX56kwb7C0+PKJfCDxAVeZwIMpxUiQYZTIw
DXVbjpcWjFYGhr8+9UFcjhi65+DJ0pKU5QWXcx0vaLGobSlnUdGRJ15vK93U+Z4FtJ6DXDkgIVx6
B8otrkugHPjHIJ8UNW8GfzT/CQziLp2xqwLeSOcK4jS0+Q/RMvpET8xGqU773xiuT3hMI7ZHg6ah
rYGxlA5mPcHJCuRDby2N70ggELoa2fLmQbVEyS7WeskdM0hUMBs5wgWJG5ILUodlD68OE51XbZTD
V5fr1cagcOrpzX7mRGPsdaURMzcT+t2NgXrJIecOLG3+GRR53Bn8KQg2W1LYBHbP3XmQRTAZm+ds
2QETmvD/TNUumpIBDptUo+oUIkp0kJi/D55YiHtS/FE4+86ACFV8tr4HswCDFCf6eVUznwRcxFWc
rHeRgXq5C2ZxZ+VXBPPKEWMxIT9SLo81mKh3Mt5eNh5we1uLCbl3dOh569hwOG+vYzqEtVy+dGLI
DHy0Wy9FooBdjohwFKgQW6QdHNYN0jCMb2cBddXp4QGfjgiuGXebqiBLMi/N5J3azHCGBJ1pdisC
DVd2NkWu3gZJIvsrmld61ORLNJOrLCzGRHSJtjMgY+7gMKFtFOTEdem4CA/forTeBL5eXkyuYy2A
2smg1wJdKiIAkvZX60/lIMYRqMkP7I7i29B5pbsGaT4pw5H/4ZYBFUvzVLekYt3aXpvHFILjgWSJ
6omkuIYpkP1bTkbrJm+6MvyEtgywht8gmacRsENsTZHa/hxSAh2kheHEgAGmr9DFlQMxmIcOhz/G
EWM+cqSifv6eN2UlhDm6Wf6mObrz1YOKnhvHCqJDo7G1qj93yipTUB9VXbRZ3upJDxABrPdyLd4q
WUGNghPGIjLM2UGC2qmbTjQK/FEdIfScel7TSNkrctwEy1KhWdbJ34gFjRVOUWkY8q7neXQ9Amej
++SDxeE3IrkxuPw7uViFWIz/Rqt98DoJe1+05mkErXlR265/Mw0GaBxq6kIDitmFoCaQ2wE8Onak
x3L1rTGKL+OJ+4D9mgf0Ea0g4T0ElKNKaE0OhWq3jLGUHipmC2bbOn+KsZdZ8fUpbLJdezWVGush
ws5aCgxA/cqWxWOpYwqE7hlN+jIaAU/PNaULUoxhmySRPeGZx10nqk7EukZEwBdzHW+V+9U0eWcv
WpSrqFkifw1ZKxGzlxTOiIGL+PaDPxyFV76SzCvZr5ILb9dNKzdxnHAtxm/EIVgpGhIYpPY69cUo
MTYpZ0u8IiRHGEv0YUPTHenMCv4aH+8yrQEi3h0ebQndO2QSq9l4gW6WTnoT4FOtrZaLy28QXg88
5mkx/SuEtaUBNcXYVIZB4QzoS+5trIlnH+jHQe5IiX7EOPp+T6o43wKE5hofYmFKrTDqIyC6MXcy
f1IBXvn3+Y9seQdfjpu8uDJuRu+wDVZW6dptrmoxRohrJVsqPHMCZ+yToUeRQVW7zlCC2dMX0Oc4
fnRT1a8HO++ZM5/eI+yIh7xbfAPkECbK5+KEeoAVqBmhFzsFjlThyUArabMnKGFax03WKD+3hO0O
TOd0k8r6Tshd3atO+3wx8kr/ub/3qvr5mjRS5G6RvaoEIrzGyXeV+qcx8RURX3QToK6nUjupOise
YoOeKJAE4rcFWwyNGa1FX7q+Z/P8VM6jXQ2RNKIm/S9QO5H4EMKyWrPoln6dd5kaaowV5fcS4kTe
EBEuIg4+4tWc3A3t7NyerhnzIRKkJ2GH/zky3ykiANE3YKQXbeDlYrgrtp4/+XfJ3Da2ZG7cQ1uw
fyouXL/knlquL2fuwL0qVDtp4HqKh0PBRExoA8tGmNkbBaqkUdWDZCfjVQiYTCS3uEBC0MCi14z2
GfOFbLqzV379BBCu++1KNUtquqbC/Mxpg4apIs7pP65qE6g8uZ1k6AVk+pRlLXWZZp7LfFvrCk+o
KbpZCA3Pa/nUvmIrAL2r5nFgsQcNKLgaIzwAQS3FoaEhAuhly6Jp6xsHmU3NMaxfgIkXgFfJiCD9
WFz36VUuhE/KbxPbE4pdaf9IAxuZYX/HiH+i1eXIPei9FW23P8tP4jpKP//l5QG5Xg2JR0FZZHWL
Ivkve0r8zb9YJLNNVb2eSThuaQDR1Jdea09UDFfQrroUwZDXP9QMhVAHLhJqf/a1MyP6yJeKzGLU
pyXN/I6w0qMgTVst7jL/EgptpwXnQ+THdJavMjuTt0rTZLEI3pFXGr6ibENKXnZsMxzswEn8AV4i
IyspvadKjMkgk0L9/OWzUqi8ybB0Q3d9QmLaui0qKOnvvyPghCllTkmopWMos+CBizJGjVvsYXIs
PkB+ZDI3fEj6fFt9NBqP/k4NAanTQ76pjd3PqfcWGoIYAhBADNoUQo9DtbTrpR06sU2KAspDLJP1
2xOdrMNwdEt3LB05z2dyBO7xIyHdT9MSFpIUjsCRkqLGVxlrEmILJsDMiiB/A+wLXZ0Lp/7juGmY
jAgucN2920+/c+2tZHjx7QjKXKe52Nrjy/Ad8bjyjX/SjjSs7K8Eb7Ds7VMRCj9k6k83m7zqaYsN
gTN3VfBoWRZNBngI0/DZYx2Fws/fQRdyIJCojnKTgry6kOkttKCB+IzDot1SkWyAJXiMzIW0k0mF
gg9Pcdzp4zzpbezsI47sKNJoy0x/MI77BAd/LWSQcmQuzwO8GYYhhMi2wKJcv86pwbxjOHewe3JN
ioaTNDZg8VK/txn7JaIF492EGJFKbYcgAE7cfRV85Qq2rmUVK5Ia0ooRU3F8ZNPPX7QVhOgrS60Q
8Wq4+R1SzKQi79mfWJCwxlQrhNlVQakhAI6d5ppO2mdz/f8QPbsTTMX61w4y/QfdfnlT9OgWLK5q
DRl9DwPX0CtUTkbxSS5cFKdzV4Wp2vEe4xnVAZ9+0FtXG40jVKVgPljTIGIJGi8Uf36NfH80wFeQ
afApVuj2voG78ZfM0bRaowd+vQ58lRfcOUJa2mgfFgf/c4Rs6XXo+sqgTjKcwv53q/7DqLkF0HHc
bL2uhvoJRMxJX3AlxriIzzhjsDMdW0N5r4yOZEohKYQc4DVfVL6K3qkYEZjgw2aB+jtJP/ioHEKq
H/43PGoXi/1sK/Jp3sbLD0y4T1zF2WWkTg2zppu3NueAISLanpXnXebNQParHuHA5516bCAWJ0EK
LSx3VxG48OEtAULEsG3cRWO2NFKEnaeassSj38XMLMf/PZWzBPAYuqu9HZ77tQypWbbv/iwwaW4B
d9Mw2PUYwEzakQGFoD556P8xlseudS4qZt/JUKxYg5Fa4u3VLsoVKKDFFvo0CK3JPRyi3pEFhA5A
mJy05uPSy6fmU+XLcNus9eOJ/HP/0A6hNblv2qyug4Ky12my47e0EIKhf/8NzOG/tbKAbestpdTL
aLxReC2WNVoiWzBZmZltRodb1Uw68x9exX6/eyRKK9km4hGOEqIrQbfIyCFKkOXs8rztaVQTTvjg
uFqnODAhNzwgPzgBcQ701UIA4NNkhgKnkg3KBbC55U9izGHAZkBVhXwxFsZM14tMoHX/w0g+j701
SuDvIOG2jcYXIciG3/hcZkSglLX4V+m7xxfa5LwYcguehjUAADp+XGviChb6hqZ5RGIsHeJ8cjKl
Z/iCWddgGm09QVdDobGZ6b3StG+7Ps3NmpG8ugP/fekVkXCc2Eoq+wzMVEgfKR3UMUsnvk71Lszz
2KO4riJW5Jz3wc0Tm/I68MTus7dfml1c1Xn0GRP4pmtZWlmHvJIwNz1DapR4KWNOyrrQaevkIKSy
H59HOjv/Jlrzd3Q9f+b/PnWz1LBLc9aBRsHfopEM26Q1zW069pWOT/QvKmd9rLThB3NjctN598NB
S+50edRMcfWtRH0czXfxrlWeY6SgTMUmQNIRcNFKQwAKX1DUc0pejNuPUPTTP+cP5688kPa5cQ29
Dm90UMZybKgHilWgKz8kD+NGOqLwbtm0wlMNurMmD7vShWGwKA0UE3DolDNQrgjWieEFKhZiPD9H
L0cINebSpi3KKRJnVxtTEW9pjczOY73QUgBfGgUgI8NlQ7OnGOPuIxga6l1O6+tqVhty5fvivh4V
UKiAB44XDKFULvqWKM4EWKfdK3i3+UF1qaMdu54zJyEfg1+LTiaaKvqJ5cZT/4NH0H40lw0rOSrP
0qPoTMqQXMV7/6RuzEzKdMvEpQh4VPIvs7gVuwBuaqPyO+6LGjO6D8LDiTOYlj6a8b8nQotgMatg
LYw6z6YZfFrx5IhGDzZUKzXj9IrnAeRdgn4axp6nBIhO7S7CoXExDqS/7fqgTlhcuCUtAn5AN2Fw
71ggBkoVCPA7CuqQjDKQvVeY4kdv/scAwxgIQdFTgFFyDus8qv2mFQSRrYBihK0mNVNJTCdfaFeu
lSgI3VvPXoE3sdI/B9H1DOxFjRFlRC3ga/aiWJzMpH1bUa3BvTGoNdnHxCvoQO8ZeYfldi2wQ4tB
9LewbuehJm1PzaRRecCrveS2mrBKQtU3/SoHB+q4E1BANIk8RgBKjZcTUUNPprQCVyHZ5+T+NQ9k
+j/qyuSfcn8WPOQOMXsUG+6CS39w6QuVpjDh4Swq/YZUF/vT8PqHXFvm/Oebj4gmByWmlTnrTAwv
TtRwaSGjeZWdlpFuaAtxOxPc/fDbJ1wu6t43wnsEd9QJslSvL2vwZzl4rNKoea+urlmK8VfL4EU+
QdfdROr6CTe5infyG728Wc4mBYDeu3nC0Tfzc5BElPeMPfVt5cStG4/a53CO1ZWbkykV8dbvM654
th7mnt48uV1M6jyXZ3DZbH/8rPZQfyarFXffp8TNBlt50yilKFWH1IV0ehUT6NuWkz9uGulu44P7
K889OGyPH+QV6qm4YVQOXlnyjvpuarNxmaPhqzvxWZyDyjR/QmbDcDfLe0nwzw7XyM4uAiJpzcRq
B/jsAlraIo4rgn3bV8riEVGTatccwXtsUEJ0CVbC8OBKDzZpFPpY3ajztYWIqFvlqIK6GW2uJnlL
zfQ4N2mQHsVzg5pUQl9541f268MxtUWAWQPbUuplb3wEQ6+PIT5If7wcEFN5uFfgWuGvd1oK1m11
IRox+UmBeFBnIQ2H+qa7S1vEZbsTbRUhbZZWRLPXA/oIUFHEiqLhuKDyeTcznpQmSCCeuUz5RIyv
okUmlVsJOq8gCxwJ8/A9DAd0Ptbe18Uc8kaaDFcyH/1k286VBOLKq4pC0zqDKRWkf9aCfE9thASC
cuCjq9KxkxmWArwImO6DRlXSJtvjLtaBaJrK8AQCCEWfgf5gDPoAYekKDn/zdk8fzBxLt/Nwv0Gr
ypMSE71JXQ/76RKYl5hkLFw7hDnNOp1J6s8SUnGuWYL4SYIq+omoZ1UA/TSVWzWRYCvSUOpCCPg/
Deoll9KBz4aAzVnSxB1Fqrdv9fV+q9g+QPN+1bzOIPFXtEBiHpJLikRM0szaosoiTi1mx3+RThl5
MTP2mq27LKIehfR1bRzivbtRFgO12u9bDqO5iBJXFG+hNJIISEpwQqG7Z5M+RgUXBXJSqwj1WPpa
yV25I/wEcP4kmKVqRP6JSyM5JPOHoI+RPTKUv3ZSwNsGBFjmBCyqrkyKunZl/rZTd6rNlXJvFI87
BiC8S9XAvobVuh8F8hNmmvn3fBWMg4EuC6+AODoyK6p++ZOSDHPy0sM6oM5dqlOdEqr7WjjVUL1Q
hafvOo8wVVdGavj88cHuvyJscRsMdXdlZ2KiEKKcRaVfT/XKZxK+Yi/oVzIgRNrmyp8aR+S4ppZW
JbnNxMosgZkEuwxxrm4x5bdnK+OuRfl/AIgx/6/vQZwvx88LdERdIapMBfiJczubAfa8VQKFpZL8
E3EXB6jE7yKlu9RGZnxz5MX+wnuf2W7xVUm5TKEvMy8CZT1mVkF8xKejfeBzbbpv4MEV9kKagTz9
eoLqXHVyWGMMtPwnNusYnwm+drDnecWw9ynyNOETOiTdBQcmD1DZKCpfe3QemXLRX81YSY6175h4
3xcGgumjmDzjaUdgs7seEjMkycGbStiUC//oABiDy/KJ09gPIIxgqFDbuFgvDCQefN3dO1e5HAZM
CwAiQp2enGum1Fq+mhGYJ7m37pAniil8+o/fkDgSGDvCI1LhY40bg9EOuz/xCrnNX4ZvOTARamjy
t1A/kS3856HtVGif81eV4/1DtRkt18ChVzPQpe3or9DdnejiH3P/qarmCPPfxowolMjSmR8hq8c/
KO8shy6kNbdhGw/o1cirJDMtl4PBItGwawx154o/6mFmnL9XiQ4hCeWm2YzGmEdNYYMa1vJGp3ua
5x3MpbGMdZX49+A+pO/XHSmGIXrrPMKnqWt097EA238xUoOmOQ0hKmr11vk8Tudf++ByPn5wKvvd
QT69CVEmZcncyRt4MGBWovs9IUWpcmS/nmqJLX6wGd7mZANcff+srSPP4tJPw+R4ofl2XpDJHnpV
PqMzkSDmos9y3RU0rfUtw5bbt8E7axEwGJsJWhenCXkpoZeh5OksNtl4rdohoTbu33qIFfsgWxg+
NJfk0X2DKM26+PdKtvEeHu/rf72V4W4z9ftZrsUHbDsU63XQdW5XkiIeuYuthgx3CsiTbtrGrpih
hUvghe/DpgxGYD+M9C5Ei5KZKMVsgtfeJX9w7QI6eLZjjg8Qq0UgN92xx7PS+bLhk9dtueHy8iHY
PyZguXSKVEB2DYtsuzY1RT2V/2P7wktwHyAdeTgKKaJHbnKnzMIpPOk5YQzN1ue8p+07U9wyM+7H
1eInBg5+8ZYf1nVhmcrYQtEOeLS2s28+DahB3KNloJwB45CpfQmlDNJHVcDUwQCIW10tf0nbDDHf
EkEB6T2w5woDcpsGNEK6zaZM7XXaIVpKpuWSP4gcd676uHHBKjJPnocADTN3NjaxSFhN03U8LZiJ
RTLqQpWVqjZiPdwI1Rj3wNpOb+LAcoD3oWun7xpR6+wEFd6u07WVHWw37yYQqxfBecmHfplKyLgB
czx51YUomt5hUsD2T9aN2et6abqe2tct9CxWFLhcJb4qlJFW9ZmCrAw25DtZYkdAQuqXFWBtcJB8
AE4DSXnwTKiUdhH0jv3gvc4XJ1oeH9B0Q+QVAStU/IWHcjr0rTRF+Kw6jqhdQzTBO9wE0VZWhuPd
5xqsvr7sm/GE+aseuXh5cUcCazgPwbnCGVSWoHJm4+S5olhR0yMW5qtLRKVRhwA6QmZlzRimoC3U
//lryzpySQqK6LlfCH6TgvTap+7+yajAp9vEeEIp4zHrAm+AJQ9zZSybGDx+pTVEeT4tALNPRnJI
MertE5PqSXKM9NVpKh6VNUFQUF84539AaXznW/9kSsVlz5mv5lQ2wvEBYmDu0E9Nt9Bq0l+hQPLh
VVLKgt5JA3pvEB6zUNgcdEmGAToQJt1zZy0EsyAVhkYgIRmlgrdLW59kjHeZ6QJ0likMy+mGfgKK
IArhYlPl3vkmazq0pVzLYFOoHlvI5d/8Gi3WXr5P3cAcAxnbw4tq8X40bQvj2j8MVzd2JYTQ4Gz5
VMYkiJnFuz3RAPfo9V15UH9krpWdRhpH9W/aWygW+zSQ2ZxT3DVBPd4GhNXs2PV+VEZAQx3pSxK3
73sAavB39XuZ4Vunmjv8f4S8VKk8QR6vFKln1mtvBMc2wgNvPm41Q8x6j1rffBhLhlahA/rYyisQ
LmOAdXO9X2Vc0YSTsGvXGI2pp8PbyvRVa95sS0JbtFo3pRBQdthz7g1v/NusYSOAsukIIoDgsQ1V
A4AEuho75pvno3uMWXHTK8U86/govGF5JExtrZ8l+To4NWpByKnQ6fcHjC8MPfsoDs+nWc9pzLaU
uvmUlu4tSdHeSK678aJSIDd4NV2Hslut1st7lhRwidSJQw0la6hWHHJEIVimG9tqzviyCxN8ubdw
mt/VEk9GqndoZxqkhVDb9fWn9i44QdUR8QOBwcqUX6FUd4BHgy4U8om92rB2uXXX1NW4+XEFOMCg
1d6ZBGQXQ2UXU9dF2CqMHqjsBGWwbFxsAMV81ELbIW87KHCcx/6xzpkDKNaErhnkDu6o1JMkLAzN
uGEU+K+/Rf6Yuvg56oeLBSO0/ra6Tm9+DyBR6q514CmqoBLKsJSkXXOuv27Q1LGOwJBTHeycEsIR
HtmTByKK+pjwqArYedXPc46cGVkVmI+Dqazf0kZzTgz7i5s/U1y6td2wT+XTQLK6wV0vuiR1YnV9
MjcmSHS9Gz0Z0oNQFLSHPvzcy62Z1xlC/cwOUxYVUO8ICM0mUmuORX/xMhe0+uzvAJiwl7XmtDwb
qHpuO0wvXvgrKjzdrlB5OZrR9Dy7PC15cAycVQDQlLod8LvdgJLEC9RdVeMtpYlbhCDxDHBk1aqV
RLTjKAWwMQYrbR+31w8IM6MHa73jlpzN40pvlAc5yxF8VSWQ9PpnYC/QS7zBrEoBCh3/HRa1TAEY
B288oHaBALPZFeGcfUN40bf1zUydbfp5vCSUpftRZ2M92QuSLEhsWqCIX/KaN8Ge1M5Y0/TYx8FY
ua1Gna/17E04WBU0UiAKmqPZ7Nm+xE3eeApxSKI6/Xg3Xahnsgpgq+SoiYn/MVuUI8Gku/+8Gkbu
ME77CcYqu2sOd3a3MY32DberfUbR6nfFzGlCOCM7LydEWV9JXbkjSlBjLhi0PTESxhmzzYmzy3gH
f163qeqSyw57wHZqNeWhzCNHKMMPvKdoQsX+oRqw5EV+pcqkpDq402xP+8SdmOdc8iKwbasWN9T0
JteHLCXtkaY8Cvin6Lr5pNlTzOLu2hxraZ1x91xuiC8PUiyQgpv0UwMXRouG846OE2LpYNfHZDMm
vaJQUt6+jshsUM5l4XcZ5kRTnyTRknl2OfQJLDA5OtAKyfK1dy7469d8usSlZrNjl7YMpaymWwYX
8wRvAg+HHPPAIetownE9yiMbajmgxAMMm3OEDAKUQeuf6x2oaTAq42XUpuJKTBJBFwsqswh+maXf
EpVzuGExa1nHsH3tQsuS+YpESOCsYt9IPT47nqmfnlOT2f6qDH0D7PxZ/hAcrI2yTWUXpYdMCTqU
4y+ZiK8PDT7BoY9gEHU1UfUbGgq8iCToxy6CfQjd4Um5hA3YmY88fA1djZv/TEV1hhJMl9EvDglh
LIhnjpVmwCWAgq9FF9v6kQ91MjMW6UdYoBSJXl7S754oUB6UvigD+J4VK1ukzKLjVqe8GqJJgkho
9wJ0mJds2LFN1mUK3uogmCB0PRwe4OqLBrIwhoQz/Y/MOl9NI5BS+FcGC5mrF/spUdOSlg/WduM9
yLiXs9aXh6spVihMfJR4GOqU5i+hagaT1M9LkAYQsRFSk6H5C+DJkz/Ily96yAV3U2izpfB6hRNU
WOwIM6bP5TjnCHP9tOF8Ffl0C3t7SyIMThsJD0SRySRNJjtX/CjgNd14cvdnjcnygAGVScsCKlp/
KHAFpSvhiE7QJtYXIJ49efzqfPSdy+uInTxsxWp9ZQc7T7CE6DcRrywt7w78tkSgxk557FeQNUk0
SyF5beIR6LOJFIN5CL4NFK9hl0TQWI+cSMNpg4dNCDaECfpVvxzuCeyj7so13C15q+JGIuDjFtAj
8ZbW8stgx1kBF47Evzyk/DsPGYPmRBSqAgKAwTNEmbuh2rSXIcknxbui6WUY5saoa6fRkVL2YT3j
oQcvMw8yvG0U3VBzYVenfbf6nAK3Q+A+h9Ssl/DKEMvtr+LpyysObrMKhRtl6uU7kXsDe0KNcptF
R3LDi2u+4ENVmLRgjL0cxGFF0xPrZXkv2soHUPjBkjcFKzwkI1+wBrXDh4hzJ7G4U/rt97uTp9qh
ySa3O1CVmL/X10hnVq72ZRaMG6cr7Ip6Ll5xRjipH482mSLgy1lh+GiGLfkVbCtuMS1vGahuNITM
3Jj6Ua1yJIcVnPoy78w0f43ManfRqb4CmbG92kAb7RzEutS3SPZQapj4w+NK8LISL9o5l9cybvu9
n6EJPQNw22G13UQPR9in9aa0+/ZP9ZVPZGTyb4biZ13nFFZWAowdbKD1tWVR3EormybBEBp3gC1I
wmV/BXseeT7PBlOEr4B7IO9OqIOu/aCE9RHPEOu98r8rJSS+Bcwe33kK9Rl7HAVrBYn+tv4W1mSk
9OjajGABfoyR/jOSff25Nxn60I1c4oBlIBn51ksFnjWxL1lDe0CeyNW6pWZc0/IMylPoXXYBnZ0z
LnLvHWsWk0belBifAU1Are5y3tpHG29gi5e4ecgy19JVSf8vEify429jr8jtwvzVp3R8UHF+8GSu
ZJMbr3Es1pEPLflhU/wp81dLmwcztZyS0XaZbPa362FMd5U7d37YQFmJalI5quF9wVM6Rfnarw5L
DE8i2sPsGb4kkL2fJpTi5Q0Cmc1bjXEVnjzNouvj2vqFe4WB9k+tZVbHl45URqmaNBnCi0gYVtyq
oQTLHc4QXFon8VsuYhV+mWgjUpkDIAl+d7R7gMZrsjM8UdXoobjmvNVK8ikJ7WkrPUEIdxYw0Avl
Jy5KFLQc7A7r+r+4d/SMTZQMeULbiB1vwiokrcgGAgXnzJbLS9TPzp11ACFktA5g3Ho8pKICwwTB
3iTMSkDguBmgvx9BMPlk9fo4i/yL7HGAeyHzCEX/BdkFEb8cualrZ+63zHAF4p4eddxEv9p0flm+
2xiuzBkA38BM7/yxvCu6DmIIVB5CtvW8o7rWKViu0KgZxXLAVjDpcTHeJESerXZ6kOUIks+Zqacu
39jrFhOVkAr8MsYZEXZ1Cp59WpoGmmd5UckoBeWsWd9K0uAxsqB56/XpFlgBi/zdE7vUXBStvyw0
oiTc8AUtXXfDsCjta52Mo6robIvsSRqFSQT1O7Nsc8JanLTkYNYje1fUO7jP9yBpyPBPC51CO0w/
QUgnTEj0pBQZMNtWk7cqBkbtYSXLdSAO5PuVTqxhn2600M687tcvBeAkVWhlZunA9L+XrpgYgiys
IBSkiz6BusDUS8KjQl3am2zypI1ox5ZNIi/iEKsztYMT7jlTMyWeD7GTwbBPRHsAgm08TBhQ1CsR
unToLHBOoo5w3NvK95RlhF2RtCG0gkeB6ZXS6XkQQhn2QEcoJnkSuLN4IC//yRQUONKLnydUjX6B
Jl8naPtkmA7y+F0ORUknY5CasV0FN74HIWHw3yPUkF1kO2EmtGN7Q7a1ElIgG91u//1PlEWJUIFh
0qXrG7i/K9GHkpSinIakDK2VnWyOGZpcB54YnD4Yp1ltxPaZbSicr0KcRK9LhCAlvlhuR9vzNaMk
U0h2S262ZNdAX7Rq49zaiL5tPJalXEpRPqGaE+q+QpoCa1aNH/h3Q7gpv4HoP+ueKb7Fd5EqkOVx
q4WvcJSAWSwdsADV0r24WsI3pnpu5OSv8hVUjxnsEB1OZ8IpC1/x1I+iuuScpVEeowPoJ4PsLb/R
3+tiCbBIZLBL9oYSGRA91K936+8NNMV5OGLIV3DphjiECjQTvap6AHoAvJA2SBl/zu2v9TbWkRQJ
qGDWJLwICGOH+M5emyFxlDYZsHYOc9jgUKqPwpewGEVJb8DEzWk0OQiGTbSlQxqXPxfY5Wb09h85
ZazA+TKuKxRKsHGpf0JwNzGOOE28/+83wVo92CmrS5pfXjtd63OxCbuy3GTHpZS14/qFBFDkZ79t
uJlA9fo1qn7YtwQDcEIDFCy88rAHM+LRSva62uzTKL25N2lVoqU36ZsNcjYxko0ANZAytAqrY5p/
W2zWllShWlIhVuIaTdDvyhlRFw1MfgrUsxRLLOkNEez3/kSYWB/REzlmT16dgUeTMzRPu4OXyz5+
CeB9zWk0lrd405FTsjYRoO9ROmkW1ckO12rtITYXKXGRMaTBkTNhqt27fhxisa5XMyL36NzcJ3XP
AqojiGxKpncFKX/X0CsQsmXUYvWSYAHHWnQYRhNQWPbfdwyRWsGCPcyuhgoGQs6mpDmKB5CItaah
Veq4FB5nbCCE8cJML7k1Ej6YZfL1WBEZ+VprQPHGTeri2O2jq7lOZSxmiyoAN/c3yerOwDMOUayj
Mtl16nDPa2wk8lfmEPikvePckcivrf0EnUNriw0rO/gOpQM8fbQcpDftcrj1Z2tIK4rn1a47cACc
vEiNMLEfbQHiGvVIFDeFdRen7RyNQNPXEStHfL0PX4kGqZIiaTztMjxCZmIJ5SPtBXPUjDUtjV5A
sW3QQGh3D2WIDHN79uKkwCHPzjmHqANc3BoF93RxvsVLT8am1yVKhMRgrSE6jB+p9SbvXx9HGoCt
+9usadi4A4Y/FAjD9QVy+b69N4D02T5vUdc31FQI31snrjjn3Nv37/e9zlaZCKDVkTejgBW/ZICl
JmzJ1t+JBiJBXrB1s+KeSzjJJBciddU4yUA+8c8m2Binznc9/W27YmrTmvddmMewBw2bjHmsv5n0
BCkLx6DEhFs187SXDY54YZt6FelZWFdduHgj9CEXF6qan3jxU93QNrHG0Z2PwCVzeHE9f0uhllQ8
L4A8hOa/GLm8kn82YNqGebY7QF4nkK7dKmoO0QX45Nsm7W94syw6F95AAV7A8aOs08JNa5luMzCn
QBBk4AXyE9uAKu7eZB+8BPqcGheos9UlGGUu6dQhdu5tUVANPE5DGK/oY7+jJIODA8RV37dVJ3J3
qpi73Mc4KOu1Jww+pzKI2M/kxb4V63Wq82XFwmFI5sp0Z1Wz1elZk8kK+BqhovxdTQgoJWVRaMi5
toKlNB/o+o6RlVqphJHFdwVuatcxq1bgQLm2qNu6hZpC4Yw00+eI1ZVo23CB7m/WGLI8EG+Hiz+l
ubtAe0kfi/5cwlTLEyvmyXTURrGHn85BxorLVhHXkcTuJ7nqnlH/z+2ScoU+VTRf5RpHz3f+8IMo
OoirvSBMI0CMqjT5U3k6cbXuzonS7sHXfV2lTgwnS/K8NJWY9Qc84VO3PCw2znevw/T5AwJ5I2P+
yod2QcEEsuEI12usaEKyuytmQl9xWC+q/btH2UEGL2yT7p1O9wk3BC2zJQvAqSFvneTYk4dyemt2
pa+grygJeoOCT7+X038UhsaqhzPtCIIp71tWHNYxBe4BGgqEATTOxyvQaqeM5mbQcCg2weXl7959
LrDUbYP7UPMIwo5E2rSmcT6Ry7NKFhS6HkHLVZ8BJrz0d9Mp75jZpP1PkeZI48EGE88dSV1mj3V6
NJGHhdTwWEmYFyPiWB3RzjGF8FUAp9VjIUSZnSb2XRWttymFfIRzYyLqod0PRrfT2CQuX2stbc0n
miikUqMlImcNE1JWaRpgBpCxF1P7g9Mvqz9/s0T+e+KRDs0rYYr9uCy20FZv/h30hYwGhLv68bf0
kCmF7Qun7ok0cr1UkTajSyR/jsE3SkKZUVOs02WnRqES6XPu956Esss7zcT0sMcd47cpaxZKyYeB
lITSGRctQCU/bN+yA0iqSp4VH6idC0A+IP0X9JGdu6qLKYNgOSbvQEwNocjoGRPHVmUzHxgerXCM
+Fa7OrZSDfhOHmFvmvFKRVPRYLGavdIwb/xOI3F5G39BHF+vjn31bVtqVTrjcar+a7nS9x6fbQ5j
ZIP2DOXcG859sXt6X0Pp0TNzEZaM95i8EiekpUaVh1wa0FSONCuXqd73kWiMPqTdmlM8fZgkoY1R
UI6ltXb498JVj3ZSVpobfcI36S3VxmVRQHUJr1RtQTniEmhxSxIoZi39y/nGaEeZCR5p6CFYYvEN
CwnBlJbe4+Vn4vDE0kBFABSFlTg28FLMUzWrxfAFKQMlP/iIMzOxw1noM00hPxIKK/Z4cBprkNRP
bwCIFhUguU5fQPER8u0XAuCPJcokAIH+GO6LQG2dEcZltx6a5h24Ol3YBLb9q1w5ZHEQ//1o06zP
9IPs3686uj6IzL0tqVVbcFiMOJBCbk8pkNWxNQ94+CZ4zy2MpyWA7GaYyhdYKMA6/GUiLj0Op9FZ
GsruMKptJWGE/l5+czB06K+nyVyigNqkv1KNsSfmiLj9Ddv/0xBpIg9WzU7BKmW8Tkgdj55vArGp
AAZ4GF6Q6ZeItp1B9m/32MsvGhKLiwjTNfclwiVU5BTXTDZr/F6MyVGWkW+df5ZSJzCZro25GIu6
nlJazHWMhaeX6+3Bo94aQty8K4mC0ALj28jnzVy+8uuRrvdFN2yZuy83Pe/VWn1Zk22/C92rK++u
vT9Iz/qQm4PWUXIBAOFrtPaGxRzlVkUrYJ+07aLczmQIGYWejX4tw2wM2EYcidPVOH/z36WOE01w
m65iEiB/4XRuLP+WNWWNnV3WAcLcE7U4EwlGpQzpk1bChQN2f9KFUwBZ3+PQ5DA1k6G8FMESb8sX
zXkRPedLx7oIvytHAjvKiSAuMsmVfbQUKrv07rUyOF1lw2eBfnqvx0Ptn04r8R5Ok1gc4J5YNGop
1UV4eZgYGdlwZ0GJcJfFFf9w8nQSqzp87FxOD19uOD6jWvlHykqqWhofZgAyFT9I9Ikm7Bko3ptw
2xTIMO0wrz5lk6PAkFidPae39yEmImYHsyFSqS5AeSg2GY0Uf2dXOV2ohIAkZah6XzKNg5toLOtk
rsmhgjSxuHy17f72sEVj68MkqFlqnbNwoPsdMJUhaW+dDVeeMoQeoUk5FNKUE+NRIoylXbpJMMrH
4HdhL1k6j7drrjUchW0oqlAtAAw3NuSCbLRoig3bOC6P3u7lt6L2CUOiYCcigp9pWQVCeim0Ue69
viA2UYSrXEPNQAoVlyZWcpv8giS4/gCtYg4jd7V5lNvfUDAHQOezd3FBJxh/2oHHQ9cbKD5YOJqj
XMToZOpHK5n6sA3lVq+0T+yt0gYJLnyP0bcmUK3lXB651dvBBmA2Yfzic+n2DxiqFIo9eV1YN9YK
juknpH8V6o0zy8wS5sGTKOSPMwR9J5KFrd7OA2weItMf9Mmk4flEm8+eSpVGd1RmvP62LwvN8wu1
6vme4awWgFkZ/MpMHqI0OAo3L1DvQ2Ry4Uhr/dSCXSzSP+KDInrpvHaG/1YAro03Ws7j9qig0jo0
55NFRt3++KNALJWb2bmVeFAjvdRlMQZOoTR9a6k7KQAvyGqeOXiRr4YqFwLog9j6DP89Xz2AnTLi
nTLQLkZAJkHe+WYVKASIl2M/0RXHe9FoMMxN7BFZM8mePBniSAAgLtDjGcbLYLK2qVBnHgqnl+Fp
hcqSmU/ylERdtsYmaH8sNsES5e8xVZ+BXVeP+CdZokUmOhHN/9/PI07FhVjk4B2zugTQ0Kt6p1G+
uZD61H1JpvUONXQQgUoWH4/PgeRj9alYh39H2wt10TsY1NQeqlYrotmza2M4swLSMQGnkGxvBQ4M
D6Wa2i9nprbtnZJsAUUuC18vWveqrLdVG//qF2xWpfIC1rjtbfG2SHrzPTBLbLXacdXDYC1IBpxc
bySgc/Wk4f801wSfVZ+mEE/ERCVfHaJ9DhMoiU1ijyz1w+qmP7Jn1khW2eIbxo3D1Uskb3+vEu6R
5mPnJOw/EHapw4Zt77GWkH8++gfT7A35YyE2aL96ETLwbdsMHXymn4Hzz8ciwm5Qau7lpiPPSD3C
sM1BDxiMvvl4Y8ow499dIBz2xYgEpVWNdL0zGGfU9lxGQwPz1Fi4iyMfDxTgYZBBs08iRrzHc0V6
zj+lphRIm00318v7MbfDuX0NGK99RL2MwSaYlA289m+sXRxPB/th1lcM69yXtV4dx7pkSx0CE+iS
4oes4c8njol3+jSXtKswsWIbdMcL8vMF8E/LKTtGsUX/imS012PQMmadnBN+0q+w260Dr7xUsMt/
BiLHvAA2ngU1td5P9Q2RW/3ANFp0/eJdz4nlYsqrx67W2F3Rnv6YF+IitPl3zntoZtiZzgU7rqml
FkqqNH737mq50no3lv7OiKZ65twWvYNVOuDwiHEQ8plBNoVQDZuhVmW9kSQQhPi5y+jnRHO32zbH
LkfztF78YjGvdfArK/27QeudlD10G4m0udXfnjuKgKbPszJD4T67nlL9+ZWpbUJ/hPC5LTKk7lyX
EQCmIWBIvVwQOfwv63shDo1RItV59v5c44Xc2AqXYyduudE9m7/aAwjytSyHGBKqreP+BdX27wPL
sBL43QGTTVgpOiXYM2+nx2QrNUK6EXSxG+SdurKn+A0i8qiLb23ly/sF8JswgOicX9dat0bkJk89
fe68slBZ8CSvHJaOzwnmiNDIkmHKJF6wVS+jPFd58mvSuL0QuzUoU24b+u46DSR2NlKhsJ2uxZKd
V13HhggUr+hcI3iHMswT6ZXiJ8f5F5bIsxCMiQWlbLiUHJIopBB/XBolpxrOYz/NDWkIUDogVYGA
oj3IsfmyoTjyijUzQcO9a9VoFylUb95++PJV7/Kq7/Hn6HObQxFgVsbcS+nv8hQE5tHPUQLqz3LC
NBvmaPnLA2cjMzdXagb06qtbTE8J94lSdoBTiCEm3Jxm7GNB6JSzASUlzMErN1uVJeYDR3H3BFG3
j2hKbPGToYal47fev+rbR6b4cR3kEx8Wyhzp5irBnkEKksyAInRDxBVtWV90ISab/OLT/MSWiyL+
v99cTthDvq1kdNvHA57PBoPUiGUfw46flq185/SQaoPiDFzUy3ZetgVL7amDJIvHqU3gSyURVOIV
CeHMMFi4iGLxbRQBndRUOO+QjGPVuI+rYu8tPEFsCl1YvD42fd2NaD+Zzw6ByZoWPJ8niHRPxBSz
07Uc5zKJUUXcHgiesUzVd5xbvqnzWxY8HBCBJmmPsycvqGq/JodSgSz6M+UFUKmw4E7CBMo29LN+
Efwx6yFKv4mqpfDjJ5GNUsTCLvtJQHYGA9+KeKQjFbx/k20V+Cli2mMD73hkvBr6eN8VJk2hf876
BvFGcZRf4B6xFUEVldU9fu5QS74H1ctfAEeHkP9DSWl8mZt5Ys0A7L7F2jfCpYzWNFrFqAe7XMRb
L11YPL+gBX2vS7legVWNp6p6sdQR8CvpJ3OtS69jBuaViXEU2jZGOkTyeJtda4Kc1lnzHr0W/DGg
hVGHLb7Mjxuv/yCDvFmWc41dF/O5h2H4Hgis/xmzDG5eFslVC+YN4Vz10/ryNuV+JEKMYsSaJ16w
WCOO1RRwaOD5fUQoMilrOEVSL/E7qbQqRv7dwpeNQ0aX75yKB6h7cGSCU73DcfZUp4hNhV766tdK
QyPxqE92cihstw1l5XefyuJNkIOa6BHZJif5uX1QQLMJKDijyjXoE9Z/qrA34L1ySafAbQtqm95v
qOBDqb1CplZwN+0z/60rxu26sfq9TUQwxvnQgzmRVAh1/32aHD3tApt7Fl7/yENT5ETPNS2dOgxi
AQxC2NBi7S2gE2zrFuLCHXWczJkGeEWrFss7YIELle5ZMDTpRVnBBBNnpc131g8Ywum4Ct1Pwt9r
jBUxdUCoOO9FKGPTPWc6Hl2NZxUyZBlc+hcOdbcQ1tLAIVaqtCqMJBi6VIM2SOZPfMjE53xWyONK
4Z+VEyFOklXRbqm3w3M3q9y/fqoSPE4OUQbzNWz1STAWeMk5jYnZNrPz+mOAZ+3DabOrmBp7ItbB
GsdXHq1B9YpQkAfoEDRD+Lis79NHyy3R21cRVzjF/3uLXzkxBY9jroThE3h7I5EUWHcyx705LDGF
aj83rgbtVasOzvqCUA3UmBTM69dhWF4DJXXNYDkGXrpvqmhxvU8lH8/kHUP+aTnWhIjkkdj0hfbV
t+drHUO/57u54tv59y7mOYZvUBbbsH/pcSrG8Ghz3zA2nHkLbTlS/QiB6rYxR5CecJ0BxzyG+ZeU
XfwXZMSt176NRGr5wSwxzgqrPkihWmEcJLRnSk7f/gnHCsVbWKG7u5Gzlr+8lUiaUD6WxKPRKyzr
Urled+6xHKTVU8qBsaf1XjfQSxVLp0OnBYPy7Kf8hRMNVTgox+ysorUqtcHiV7ucC0uL8JnF7O11
YZEOZRvzSF+pCy2Yqt8RzfUSTTTNaDX4NQ9np/w/mmUr4FsAxmm53xn/Gey2i3I7tyz8kXFOQ5qX
Zw3hQ6jXFtGHXI0FIFlq7a0uey8qwC90e/4R7yKr/9vxgKtKAB4I6Ep6V2C7o3SBItogAbMzjD9d
PMUyjnEZiZjzB5LaFgGm7HHeTCnlTzeaH8N84ZPyfpgtOokXnZ2NJMZNc++faMAsnXMOWD8WkSXP
4hTrUtY1pyLg76yd8JiAV3ivuH0spsBXGA28PHEu/ANV/f9HO/jfuZ0OMx6KyZl1tfl/v7uYA7WK
13vjw8sg75KDcd6LLU4feO/Nke2hJERp0mdSHlbkEkq2ZeE5j8+oWFSwi/LEOyV4M2GbiX8+F/i7
R1ZdevtpjVEUcrExGjQMe3bJctGaOH+V29RVCaq5Cm83zvujSxE4yrQkkjvgc7RCH0J3CUGHWxxV
ONCcBvuHzEKxBqbJaJG55RPYJZUOCb10/R5fEjAveOgatG6uBzbiIE1KeN+nuhlCN32cz2PP6wHH
XbgA3FUTQNnoZz09AszL3pEUqjYQwbBCVnXkJWFybd+PqWMl1zBda3ix8dSvoCxC2pp8hCZnqw0w
6iHNhoavdnV5yZjSKXmr9WjXTlSu5eKu+E0l0R9u6H7lCZJ7OAXfuqmkFZURlaqqSWzO/8oXfWC5
c4jILBeLbinDjtxlLbSWvpQ/h0SQRB+JL8/JvZ58gdNzRN3myQTpkAhx/E5p45kgPZUKWDc9Lmrj
iVjfhBeYoCo7RnhFXXeLGoIqySsAddfudOuMclXeFiavM53ghPIzetiqIdSpRRPohMTuJrd9l0Xb
eLVY8waZtoMRNtHdt51cbZozPXzr7M9WHdbpxSlzwU4erU/zDsv7Nw7JMN6Llgwkv9Q+y6U18mwO
6eZVFRv3CKp5B8fdA6e+LquTsd5azBKXdgLQ3hRVFqPaTwcd5nuT/vD6rvDqFaXrfwwjH4KbPd6k
P6yMVkt7UjPnoyegxaTwqzcvft3nI0aYdQXVxQOXYnFGrPk1JOqVE/tCaQCoggsa9hKzQhaLUka1
rjIXDkk1oILKCk/PkRYy4W800PaNr8B4KMaIs4VFlzU+SUJCi+uaWkcV5Ul1gmupIVQKd1ZXrMuB
9O792XwbfYxLfUCu5b8F/UXiPFB2Z60LVQzk/kkqDxc5mdpV/kc6QAzvE+q3uynWcQLBKFVWwY9B
uJHA6gv2K5E2Ump6BC/35W8wKhU8Jcdgcf0U7trkMpQDrqGPCZx2ppxz5JIjsMe+iVPTjjXaQ82G
t3Rh9LhRPOH0hgpb32c61XRoaRFEekolJlMwG5qRIa0ruwP03UCReIM4X45Md+WmVPzoin09HxJ4
uTVdsl7LOpJcjBBF5VpCC53q6rBX7sdKyyQ1uSqrgObB8Fg0yLkngeD4c0sCIcys171rnhyoegrd
U9dZq8eQ9AW6klEuNi/OZGBcqAZYl/ib+3gnxvvuLwDlMVGbzJPd1+k3AJ4zujd2P/rEX432hGfO
djfBJphKj3RzS7d5wT6FIQUoV4AwqiUO27ndo3obwBwdXbxnp8qwFfN6FzLRoQtuEC7yxZae/sIl
x9yZG65AYF33n3APmQZAoUlgemLes0Y0z/JyC24eiF/amUDaFP16lVbYiQC+WBd7BQA79XO29fg8
qm39HIiQYuk1vdh64SmaM+cNzCZYIGngHPbh/y8CBeZblgkI8Eg/hsax9A8klJod0hkjXY1ucrnt
DjXoGu8hn1F8spz+IX+0tK6pRo3uTRLaj+DS+HsOMDmLdGQVU8X1il6CRXJBL6i7nrVBS5I09Zqy
lerzDDwYZ9aJgRaFvjDII1crv23QwPgEI3V3wPFhk2PnMVC+/PZ61VbMfPafTb9MxWYjmU3IVpQU
BtiZX/iqjxyJ+0Rkx8ulLHNzQRNIjdQLV76xCvwIVQsgxfM+A2jnlQswgkeK4VZbkNGuCKtf0JXy
omkQ2MQ/v4/gGSOeYfJLzbo3FlKY4N9qMyeP3Uhj7owfg8U/ndIN9FBMrskduDiNw+wLL39+FbHB
MBuL3OINKZ/O4cEuPIytoee4R2xoCqYhPHC/gGsQHaiVrSMEmiR8ogoLk1Pay8hb6/JTo6LdoB3Q
XbhvX59xPMVIFqh4B9pIY+i77opACNcLUisG+coOzd5VJgs2BDGpwOQvvxo/zr6luzQ0Uuegzwqo
OXo+t3QgGevzuviR6ecSBgro0oX8Dy3KyiBfNHdSaf5dq4HUJlaGj+7lrLpRDSFocW2yL+DXU3sb
P9gxVDE/I13VcBTak5rU0jk+R72Tw8y/bhUH1+t4RPldf6Y4cEVg5i3RF2x3Qri2gk3jX2mHoezT
AyY8UpoQRFJW3umVgfMdyxIzvIeElwiTl5pABJCiw7bAs6yANXPW8plwznKE4LgY+MimbhWhF3i2
EYvkC8I18bmoW5E24yEpIP/MDB2rPg/k2Yw3ojPV8ezdt80kpbi0RYJbXMbrSR7JOuD5hw/OPJuo
xsf437R57UxXc4XfkhXdQbXgvlBC6cnlTEtDvfWEzp1P88NUwZ5TZZLpYpEFiRMUs3PynqksGUK1
w4znU2uiOC8+jUwQAkKrJSs59pAMGY1U+cN8rKF7GXTCEHudu6i1hnRgez15cohCIFz06TeogeYr
+uuREvIsmlm6SbTWal8EnRREF981mb4KG5r/KQrlUNXaTDcPSHTDmfF0Fki2oMIaVEeF93v4as89
jyOisP2FqwdO9ZivSheGBn8/OqonqyprYV3j+XPCiJeQO3JOZCCR+awYjhIEJir9UsLiX11+WaAF
FBI2RgORMk5sM6rwuRtXpT7F1hOSoOdlOGrIO3qkNcANiMKDj9XMdfHzSYQCk5dcMIu1z647yyxG
yrYwxPHg7mE4JgS1JoqZoq4hsyyriIjv2q/5Nx5w41BmwV0BwibT4mnA6H0YEum7/bUQAodozHho
K2KEEfN/zYX8WNzCJSEFkerjL4gtio9J7idVRdBpCgk9GOxhidnlfJVaARi4MH6Vxn6Y0I7OdRNJ
Oh+Unbz8k07XnxY/u5ZB7TmzH6GJ8/TRVSQulykOmNCrWjkumbjt3Vb1tSzlogw7NbYErr2Ssl3O
RV2SdvLTra3uhl2x1Li9CUrwAI7eR/slOramYkjKzoK0B6pnyhy9cX6v5WxOZUqXPwjnPC12FyHn
hGmE711LyrSOpAFXxxQZJZy2sGrJd5Kcqcuj5sjY3s0oviT9BfahUA4+k5gKn1X3jmAXVMMJ9dD5
NX04JiD/wJ+mX/NTHhYS4pHhBPLDPhkEqurqO8yPi4qdgtiVXG/uf00OOsUatMmzkMcDZzKDPNNO
8x6M2jeqxvgEFZnqTRN+2Lxs5jEfRssyrUDxggTM4sy9CyGvHaGHr9+Ix6ZFFeVjohnOZ8sPuTQb
zIQP0rqcKrmqRLHg3Lh3vI6danRQ+WvQIhzYqqrZlFwjMziSUXkPn/nJdBgqmhuf4AprD+3d1nBG
E9fpMQ+GalT4ZvwvEWoIDKutzg6UKWr2V91IphrdMGxt/Pe8kf7LP3a9UYCWU3FHm50aTy9EEMyo
r2AU6Q82MRdBehEjsgulV2n7pAiV6LnVr4ySmMVsSulMfL5e0ZNwFQmicXJPcm8jf/FTGd5X5FWX
2uFGkOe50oVBczd6SPS8wziG+AXzFkblOtoxrbnInPlkG8UVLCDR5A+dmnT9Q+dzMH926dBR1zOD
noWUXkqaqpZdeRgehhNOyvrDLVEdX3n8VzYja7McUCt8fQq7YDFsaka6WMatHRLp5R+auhphBKHi
uOAkFT+xEP9YcKb0nshfR/PafaGHL34O+Vb4UA0O7bl/oEFa6vL3xfs+Cv35dHjWm9PmnXFDgk2a
S7vkfAV36Lm2Ue7OjWcbcPzCj8p58dl/cmEG1fTrVqZpIwIb258hJjtX6g13NXllNeyOXWUg1AWK
7LUuqbysQvAWuTUBC7PxrCev1CFMB04LE9eNZxm79zW7g/+qrO0iT5MKyMixvITuyVKoBe5MB+nv
mOJCTREZ/ete3b3/OPFRJk5bcyPtXCsUmT5Awn5sHv1cbtwBhJ0kdwI/4/anHu6by7AjP2hwsW7n
soBfeDrmGIgSQoG2K184x9HnnMRTwMWShAm719GxQUqVOWjLcDptK/BGozMQTJ4GMimrywVDiL0O
aKjgsp/T0Hzop2hgqVTDSRsyOsC9af13vPNQQz9mPPni5CUNDKlSNO4SNY1yLab5lo7Uzl0FaZF4
6j5PY+1NHUgAH4J4R0fwgUuhkE/Hm6Jx2o/RbywKA/djdup1GDksXi3fq7C/p4TD3B5u7DWGOVtG
idrsq85Af498E57w20HNZbeiHw+dZRtrCvdvy7NLDJQrI+AYbXTmum34ZmXYK491bF0U+8OZpe5k
C0BdfySSOmr9P/nY+QHesd5yZLaWcfugeq2ZeOfckx7Ji8A9z1WVKVcSG1BzYc3QbU0BcEsiDWd9
zRUPSFUcrk8J219+CgZOyxjcQ1MwgOnEKG8FaW/s3uPRoK/EbVBUdVE5k0xFyHwcrj6NQXdXR7f9
6E7PcZj56M543l24FoUn3yH4FSDlJUq/2iPZzT60lyC61aia3k7jppMMjdw0SZybQ6XML14O8w4y
wPXZItL18dfJAgkMH4hBGwragJA2UedxpsIA1Mloe4r11HZVggIYnqI+0f7UG4uLH6l18KjnMpGS
VOhNQIBVsFBGGGQ/6u1aMFGpVplbTq0CSmBqBBfQnPw83tltXf0PTrlj/DVwhaxnQ/xkMPFCSNNU
V7frSwuAte8YfWizd7jNu0K42duQ/NkStRpBp0dNM/Zz3wBweXLHVWyK/b90/2oCa+U234kYqJ+J
xyHQrON/xU3623YmqVho6NXKi7s8u/rQRNLd2vshbhgWEwyt/+LUFAxMdtMA/tOBhuPxgPKgS3Pl
l+B3oviXLLV9g63xF10AO03PoGtIMQd7wfGMJxywGQE64+RH9aNttO1bnGZPWj0UM+OVMQZ326Kp
c5mWMN7slmUrWelyVWJQLF0Hrv0kT/5StdQf8DCpUVi/ACVqcybi4Isiy7GVhuWrXrORZrBjg60m
etIg7ACDXMAQ+yOc/+xiWwnFjvtbxbXXXdLi3Ue1XuwfE2QirSc5+BH7le9pG/CkO278mffwM4ae
5ajVq7RxBjjhSldExkD4fWPKknlCpq9rAkKqhAiBOxuYDPirZJDs6hcHG8bIeydgwyQYpSj4Z659
qaIPCz9j4/335FypGieqETjF4Q0Vds6tKgrYDEA3iqU4BLp83x/HIKWEXj9QG/Je2gktf+9Zg3lY
SbZSNqKUJeaRle2ifmzGvNjGWdexWKR9hiwZGpgZdB7kdQRQ+OzTcWOGsH4zUcV67Hegp6qpPMNM
nE1eta8KuqpQzhIy2XrtBRXEUM4eFItI/ITFAiIQaY41MKx2B0QPPn/+cWtcc9cfEO+1LBqZnS43
dr9Mp2sTSKwdXswLXDkbBxTPjGVk49qti5d6mseS7RmauHh0Rm/ICmcVo4HPPcZSElweHiirltMx
Iw+xqGKCUgucNEeP4YqpZDOJmS2ZjEkv1aWlWCNtP6DDUm+tyOJuzFEze+R3Ip9iubfwtwHcZKRY
702Bgfp24H0oP1fEiKKX94jMyKGsg66y4axQNIyAtoiGn3/TcMTEskyG9qEEzADkO580E+1/GgYM
lOhrhAFeVzeZ0UyXw8K5aZESDaZnJ5LM1LaaLoO+U2PMT0uqZ+fwQF+yw9q8Y+pXQ/SyLdMNGw3p
1Tq512imfaFadbmQve6Fk3OfBb8KSvYjG7cuN7Ddhc119W15HE0TTiIeCSOx0MtFzyTxG3R99mto
0OYSojMgSCjs+SaiG5Ipu1OrtYkuphAIz3Tbu6xSCP7rRxw0Qdq1B4C7MkVjvuV8O5LDMD/CNMw1
kK5SMq+zkKc+sA5M/aBzHyw8MKxdfBz36NlC6W84sFTwpwNeQCCImb1hJ7OzVJDxl2y48cSXfLXZ
Deipdo5b6CLZIcrpyQVTG5/KVCXPKA1EF3UC0Ka9yh6U0nV+NYMar/9ywFmysKDfXtDS5rnk0aQs
pFs+XcAzHWV5Uk6Vz/F03HMNlMgMg7DvRoMfkDIIkink/3bl/3AcmquPblA6KcxMIhajgAxrWD53
w+SGcZR7/jUgPTqY//0AGSMxELGn9s3u0vFqk7srX+jC8BC1LfvUqhlZ7CXC3mp9ExenoyxMEnRZ
H42TY12FbiBupvW99S//nJmFEHhIQgrwMRteRFgAC74KIi9EGXM1UZy4M8MM5pZW3K8MUnKwKIBs
pK5QuxPLv1PJ2XhSFaHRw7rR7wCxeODcVUm4i99yB+7XxGATDf1Kyx4ud8xp3dyQDt1ypqhTT5IR
vmS/GFArXQgANEZf2VwzXQlD7ViCP5gYQAIx2/tEbxxQS+S/yvYTYdfTbpHtCC2qOcwSt5HFW2IZ
2eK1MhnBBzNjL8p2+EaA2lOemN/5WcX6IZMDDA+SbAyRWFGBcmOOD7rdv4KfDtbXm9FIBV0S5E4z
uVsJn6vUk6/1N5u+pSbGJJf5yHvXniHwd9MDtntt19cz444vdQ/Ud+bl1Zw0aVSNPep2dLnLUwZF
rtvGF0JvldzF9U/tvEo51c2vMOVZNtY0P2677U9hlpuEJ6ZIfLu/elhIUAQy/T8T219mcaVTcm5y
4mv3HJdaUdlTCOusJO1pOMdH+cPapONofT8jxK+rqgxCEGnId3ztlPzNIdZVhG+Q2G9swkGvIn+D
WX1uEpcx2iVgl/7OpOZN/vphewooq6ivRCOVU78nJ5HFChvkuoz+371sUyPdSqkLUZvx0IVZYZg0
BfI4IMqm5cYolRxC7mujEzJUD1pCoganL7IO/DWqjjIlrzFrkv4nqXyLD1heM4QtCKca3gimDqoP
UDqW7SbxNU0rp4rGpPFNHpynHMoyJvtA4imUMCRg/5C9RoQHqlmAVnfooke5ENuClDPbY0+h+NXs
Yr+NAjdWYzLSogtWiHaH9Y18EC/IT4KIqzRj22cHB9NvjwGV7rDrZxWFzdArrhc59SlG6QhJ/zm2
xXLd6s6vZsmX11Re7FcuH4WMiTA0eWHqbphwqXLNKt96aF0bagad6Bl3jqB2VknNmgYxecLCZ1N/
KpS11Q4LPGUFqyfR5/fEVSIN7p9u/5X+qD6KSRTlbPO7Nl6ChlUJse2T/Wc74SZHBtiy5lD0bJok
Pdi5dAChZrNsbmWorKZ2dft8teI4A1LN1gBhVpSywWstGoMW819TgJm4iGp71XuR5cI76i/Ol+7s
Fr3RCiZqR0738PlrXfx/SGu+POWB8uXHxCof006y+moGXtPluub7bYWHgz4nope8hBXNZnghfGhI
3CHuCdhTciTgisWH/L1/y0o3O3gqwxPntJpAGaQihqEY6AOwLUif86wXzKabrOeBQX2q2frRyG2s
/TjgkzzYIY+aRTNvURA2+NTVF0wZ7CHbReBcX0KFyDSLzW+qxsqERuBjjmevTC2eECCaUcQn3kAq
6AnO/ZsMfN4sqDCovtdiGS6EM3HfPr5cAGmMlzR85Afjs3FjFs6Mlo1oUl1vI/5uHHyVd2xFt7xZ
JH/frkCkR9LuJDydiO6G3ZUW81qdtCTSGiHRgQGSCHx7Dfy5Ub70BrQDkB08RYFV/2Z+4CoxSmFw
9cuYDXDHhwU0kIxD7KeXWGt6Nl1UFfjZbBMdyRVU47+yda+XVXkFxsMuNMnfMyyVpCu/vC+eS1t4
Y4mho4F9hMErsNyxbR7yHB2h04C1SaQByCVycJSBi1mqi7XBkVkyen09Pcrza8zxbKlssYBzCr8P
CrBv3xGk/lgrSjSvyWwpVCNNIPXh4ct3KNHOz1spuSNvYOBdpZ0jljoK/7PLs3ud7k0+Aj/0GxWk
dlPeKCNUVrIcD5srFKzSHQF+tjh8qapTgQlWMUFocfNfDIXhTcK5j4yKOxtbVA4FMCXt1pXxofkI
njc3j2iMYik3tzpsmkml6xMvNh49Idg7Iw8WjFg0NsfEsnkswAvmQ566ZTpjub9L2fQvFFU0mayj
7k7SlSgAVTv3GDUQl/MYoqyYf5aGsqMDDakPTxcrQG3Xnqo1DGyuwXAXq23L2XGPNv6WWTJWbCPP
n5LZTx3UtZSDzEJdJ0h9vwfFT3FN0UIPnZJsOW52gGnbMDc1aquvSRU49AYwfaC6GImjRIc9e+xm
yTCMiaN9zRr5/DSluEXhhAHdAzRQn0X37q7qb/fi142yozpjeEgzREIgr/QlFRhWPgjA/zVNHlB7
yBE49oOw7FL+vFyLykcVQ+KwZCJH7Wa1HbA8PP2OEl6eoN1uNA8jGW2LdYQ3BB3Irg73KDbHTL8Z
axTl729RHVh3snnUmjPUCRXNdYOV7HFcPUwZQzyiK1ZH9hPfyNoS8DPJaOw5wyYjLg9lSyRWTqN0
8Sung1QMXxoXynYhTHv+6o5j4vahlFYeqGnoKkaDewNQpUmTr4S65di7HfBQaJWcnIKbnRJaQgkV
gb37QL9W5Do77mwrHqdV6IBohhhKnrExrgaG1ZSLU7qDvA0FpdzWFscyJ257Vp1ncwZXVIHi3wox
Kdb+3+DBAp8SAds2WRRrTTn+VL9cJse54jV5oJYqxnmNHl61YF6JbSF4LZMUf9tQvGIXYmy0sUWe
F81mocQZSMNNpXtC0gI+vB5DFT4iygT6dcfXAo+QvB1wzu3t/7WEOAl5wBtsuvlJsXaL1WunJdC0
ESYL59wp4S3b41s4AHOaw4MSPbDMwJHWIeIj3QucBqvTGsENiFekfbuZp4/Dth29PVtM7Sl7LGU9
E/Ixo2bsnPYabGxtFt/omQBCrC2M11GS5O9z1908FVt1oYrB5sPniB2iBiyS8iWB1p6/j6BJP0fx
HYHPnzea80BxzwK+Z8j9DkEs8fKZoM+KRmzn4HtQST3bAdvVxpcYIDv65jFzBa4p02DNFDKVPChA
ersqhST3z273/yAi4trZFSE1s1gbaeKDLk27/ObSgt9V7y3TZr1SVmw1TY1eySA6uK2JQFKoyfV8
Evd1ETfGqsWEkB+5755Yx5yCdArvPIpEltp1pEAXUYS4xPKhceONQAiQH4GKWERPfn/nNc0OTEAA
5IQAhcpaOv6owlD+VFLr9tR+j4CJahkIkFrINusSoSFfhrAQOlnn2tj/eu7iOJoKJNVjJ8kLFdqO
nJG91taRVu4yDN6GFhmb65XEtvv9CXJ97+VrSV03/lqCjqtCgJhER0pdlybvsPWeI6hmXqTNWepa
qUHi7f72SRwjWIGelfRV1l8rLc5BS68cVKffHPpf+XFyI0swBpEFTLriDuUjVAtGkfGpBlbsRU/H
HbLWLnhyQd13QWy4iklLj6TIfPW95Y4kxWRO8+HezX5yom1AiiQj4ee3bxc2WxI9QeYCa/iKWjQW
h4z8HDBCjph61hrGLJeiQldP3LepdnMfAJURl+0p6C5bTME/7UuI7hqhvgsTwc53CXmTARZh/6zb
8pWtoMPNZFHzYRU/jfsF19rqrEB4DDSSp/28csCZWT2eknNGetWGgqvx3AxzJS5nCj+G/lthnJdU
EK+8QetRVfboOwlsa8dueDJlgvwOfF7tN9hgYElHR0G9y0acHAdodobwaeU6Wy/Frq5na8f9n+dh
iQYv5zau6hWA64Chw/zDcO2VDnb6Fq2nDlDp1e7GxjZ/z5raJlLzCrOHfEOOCxby7ixOWNYxGr4h
+0kx01jme4Q4A/osNkptFEzvZzkGfNtuJU2/Z5J8V5QIFR++F99Ft9emg4zW5xglmqJjFrpuOnPn
t4uWfAjeweQ9YTYQDjAxLt3l1BB5fCcRR9PkhgHW0wmKto/xXsUdbFTNQKSmPZMhVNBfHyHh9o4G
DtgOr3rRwH5SC73IDKoOBIXEdq2FUwzZkpfZ8rO8A3i7+p6BcyQtdpmm3muAQrFlzmVB1O4Cxy1D
n7Hhd32dtZ1G/0ZM88lHjUbiB7oQih1c+Op8rqhmSyzhsQb2PUnzdY1AjBmozuh87gVsNLBBFDr+
8HkiWqcdpLwXkmAooSxMyYx2mS/aElw9jenWm4sT67FoR2c1vfcSmNCbjRjCyqtKyeIT4ecfB/Ej
0oFWhHiJW3ypqx/wyTke8zL1kHez+GQNSKY2ZfhUUNeqt5WtRHqfaGKS/1fXc+ZmIwnzo1O+Uh1U
lz9Att/pz/EYoL1w4hUrI/7qlaPCfa56u9ZfRrHaQvzzBTu4b1Rn9vSZgd6EREVgdKJDNHbr753h
CPz/F0UoX83j/QydNfPUrn3pDK1mO6gyvyDI17TGITiun9BS/F4MnEAu9SXLq5ZwQFDxzIF7FY3k
7Nz0ZltAoOV6anzuNNjs8FNkw8NgPUQ1yUe5b00wOrHKJ14ZRz9X04gh648cFQkm0cOkLpBle+IV
uKr8zHL/tV98FuyhepHcE++vKc6bGDGNw4zyZBayt9UHYK/1M9g7fG1XcYjVkzQxOT3J94VT30Iz
sP2OekAPkheQWcaeH826bkmUFKJ5LfiFXbB6w5EYtq7tcljcUR56iqEx78hzW3rvH76bb45GAjkV
RSkmjQNfGEq2FnC+zvEKCIVucA2Up65KUWwbrop1OVmcn4DC00B8PzCgeV+bLosti/FKaD7Tq45n
SKQr2Rll/AFt5m/bgipeSEt55mZmx69l1OguB5XzuCZvUO1E5qyUqCGzyjsnyZWejbAIpS18w7jp
CfdHDkd9V6GJx44M/dfwOmRvecdpUYNppf4kStVc1rFxcLysF63ykw3S5y48EkglQmKlUy6xEsp+
hu/iVBqaFVdFcy4N0putg1wVEjnZhIQNNqjTWtOLxndvHbLycwpW3Alu0Y7ZZLGLCCOvusiGYEDq
J8gXrVuPb6o23wb01hpihZUCQi1Vik3TKXW6HofU0NV8DvRkI+jMuMbW8PrjBLHDb6czy9xTSMf6
mozQ8Pt867iN9kSInjdGVflifBedO3Si7YGmUtbV7pJxuEx0eZIPAW+UXUlYbXop6CnKMb6kPxBp
dWajWNm5WjfS9HGHjjd8uCcbYVVEK7MZMfd4lxzsBecdx6K28pIC/Lcba8TSrJakJjWJ6Inxq91f
RDRHf5ozQw1MOiB5frAKDhWEgama10VLFSWjUgclLnfyIZvBSwBdsHR3LsopLYMr4RaKpkqC7myj
nPIMlGmf3Wz/d6ZVJGY2oMtWB6Zcn530atpRYAx1nBONCm6FPB9JKBqyOvGOl2xHZnGnbHDWtPNz
keFmXEx3Mzx+WgkiqvP+72chcMZ1f3kaBh4P95uNrP5b2S1YOujyqTn2yjNVJLKTq3kEXIaTLSO7
qLEMuSz0YYwn6lzbUmc9CiRW3sEFl52uh+AN8Cxs1qz5uESoXeDIHWKudDjd56L9ftjCP2knJqKZ
ANX3FjW9MDG4oRIOf2v87mHzrmUFgL90JU6sNrBxiSpn61XpU6+iuoxk2mMvidqBpOPBT99BnSpn
0eoo1ivZcya7BzXNw/qjqbn8UDdcnjEb6PrqMPZ8g2b8rKl5GrD3IzVp9NHvfi6nLVsbVSmkL3Em
vgbEAV5lsgnd874vGpH4+9/KP7B42a9cEAG2Sv5zxY4eSa7DQJKXiHycmWScqjuZDVl6enBwAXBg
qGPGa3YWE/5rnl6MmyLWxwb8ecG9XcHhRirflJs0G8aYCGj12xMZzQ4ZWuf58MruEnHZo+cNhVMh
7PdDEdR1b6yjFqIqbxdx+OHbGt3Fes2jLDP5OXQR8qe56r8CcSa7SHW1wOZ/Qdqes+bpJReaZug5
Nxaw3BQtisRewl+EiI3HsSOLT6K1NHzOJzQY9ZssKNOfFxhKN3I0DYWfChnMJE3WtBJH6yMOf0cZ
Haq4oUbxWK6WvzRQXaI8qtVhZ/bazLvNdNVcjDd/TwZUAoO2iQrHg6jl+OFFe8Y0xSOMRImUIOma
8Cj6yJ+o3Bf9zLYbgVZ1/0h2+/eRTnFKu6Y1Ln3QTG298/1HJHcYOY4/CURHeTT+8Yh2uGlyDsKc
hOZ7aV3I09dsaSkNaG5rvhP36zZkAqRAPDxYaPt7bk7WRnMFIjCdUhdiAkOI4p89k7DPROsriXFB
HR1LUV8wOTCX5dskw08jW55JBsEghABK0loL6helQ2ea2uW6rd9mRQhYKW/pgD619v9H6JT8C+nm
HGqRbjoWFdfM273sDG8upEck1ZchLdLcx1S00dtLJjzHFdRTp7ZLsoJDQWYstY10+bnrX88UX2ww
R87rQ1Kx9u7XhXOs/NwgfpTyWsReiBri+HCuEMAISC7W3WLjnX8mxQgAU1enmJBDG8+SQhTN9X9Z
0p8yxd+3od4APdEVH5m9aLTOdm5FDgN9cX+quDNvLHR1LuGSQW9tQ0SnWWTggsFC6EpCOfnaFJqG
scgYbNMva53mX7CCjEFo2aW/9D5udsTDNXGuN6A5Mb0gV4Vbw/VFAs2+rFnrpriliEdG7MptItpl
2iFMgkUJIBt9hdPK3PiobEhmAoMTaEMVRLrpN1ELgHP4asVyxxpr8GHSq5F1rZveovCIKGB3FlON
7F30bQAfZlT8so+ZH7h211sSTIlyYtxbxVGj9kxx+IExu9XhF9y5GBf8RvRudZAI54saUzRtV+Xd
knDpt5LHvzG8DBRMZpedZG/Pc0djn47UKA3aNZGMjj4FykYgVpjkcjNgs6E5aMJsQUr7xLN1OyWD
SvbIW4tFTxU+8Ilb1V5l5X8/wkS2y/1NqZhiMiIi7vYm9UdH4YZQ8iJ9CAEkKtSwFdCWiVWlTUy0
YcW8ZLYr4jT8YzblBGug9bkBlMx+ndc2YyFuMGebToPfLk6OU5yrlh4O1WxAB/2VROkFJssllAch
2ZheJJjHjqRF5JmZC8SH4zRyOtjAyndYH47RiwUzbQayh5Dk4bXwkwO3cOS0VSVScOLAImGdVlqz
3nm5C5uCATChZCmOQLae6OLxCI1axIdNdTLz+PE1FbM4dOj0YQaTdoDbhUKzAfLRZh3cIKRD5gcY
AK7QdVVjYpkDGf1BZIvOMVaNhmc4Bqjvl0rczYXpMWezmOkWpE9fwRIXEmiIPPCBD01U2TwUuToe
QCKe7iP2viiyd2EP+e6MLK3zoIdqH9cq7ptIFzxl9ufarWwqgBmmXR5ghSqFn2H2sWCr7ogGFnvd
VD2oFp28EKlI1U+wjasLHg0gDShNICZa9KZ8lmrKSa5sji1e27kBDCYf2hL+vbppa8297CAn4C4V
XQdYMRfeCxYKg+DsYjHlj/vtiBMHaWoDV9bTMnbp/j8l38f3HbVhycM7vz8M5RhrNAs20Zc9/yU/
wdEy13rz2pZ2fdP9f1h9T4z0Ms/N8bzXtZNImF99iJB09++SCdS8hmImWHNGECvuuH1ZYTGVp7kW
aS1wg7W3Np8V/B4cqFn/Uw2VP0dTVGwSjv8yA17od4H98HRd1lUMyAkCMPu/TY7Gjab/hrKglmqt
+5qxkveyZBQ1PYH5UtNHS6vYeTh7/Qy6f6bpe8RWOnwwUWGE9qjnwz6R15VksOclB3xLEJgq/jvt
kS0hYmQ8lpgMm8N2CEjwiNJ2YNqcZUFK24qmb75yMgW3RCSmwpQjfUbCKVmXO5MV3UZK4SnEb/Vt
l3SemnpGsWUY8rbijd2hpFYyWgadtfI8xx22gBo2TU6gAK6hbuSXMo3hBw0fBbdZoe2ej1ncjyiU
ZiL9yIfzQqKbrKZ5qxUCMx9B5eMzAgF3h2slvf77SYNX1fIm16LS3Cpbkej6gcc8hIkjAv5R04mT
zSeJ8VUC0I9n5MmhetN1BU03uF7XHfpbsjNOA7saW/9AzP7Z3XFjBPWM2KOAa3WgYapkeTaMj9Hx
xFcDaAOjZLYob41wacWjz8OhSGw44fyxJKH6veHuO7m2hLfCNFouXwhLLks+zTKSci5z8CHADtXf
BApcFL0hdsfRaG7eGkQd6VH517PvUcG5El1KzurYVi/PiSiM98Zhqny2/8D1Y3FNHJ8E7I1eOVyj
MbNPJ5rKHD/sl28D/ScFGwZwYoC8Mw4xtc1BU11xtukU9Qq5jSOTZ7whbX/EEUT1THS7Q2m2yhdc
Ffq1nLwqKT622gxB//4Zi+HT7hq4TIu9bARZMyMrLBXN96MNgLRT7Vvw/2q2VqIC1yYe6EF7ngTc
7pSfzf6RHF3jE3jUTUUHuyNGuBfpVNqxy2dumVEdJJq8uUPqYzwn4UCYkG855gbxJfUg91nek4f9
I0lo9LoDkBQU6zSTziJLaAq0l8FlOeGf0lTFriQ1iwu0/Yey4XKsnpbF60hLT86lx2iEBTBnSucr
eDUXEfJ32YfG3Yx5FcwX7XwnXbNZmDXfk64IlwwkHsxFB9Br6bSIHypHqsMdpvKTDY9YmOSks5bq
KMN/D/DvayI234GuZjLyi7cN0SOciZYIoYAoTrZgsnRaVrpxVk2Sm3ENxKeiw6oiptO8dpPCAbwZ
ujmfdHQciqP06mHG+kVijCXSgFRGLSNK+C0PfBxBh81ZoiTjQxPNdoCfDS8PMJFmJttz+anbVd82
8zrm/OglpU+LTIevt+2lkhBm8jlopW6ZPzruxx9AL38CcubruljSIq61xtllowGZbQio4nPwwKO7
HNCRnHlmiuN/JJWrfTIo3EKom1YLjyIFDEPP8d4dyBr75+waPEgoVK8icAgKsiwJcj7xyoq0cTEA
R2akvSQupCfT/SvGOu8ioX7QMFWuf+KsDWtsERgHUE8KFmzlefnk2VWJ94UKnEw0AjhXYzwVGFIX
jDeviRlgXda5RHbh4Wv7CFp3qryb2T4/Wu/9SLVemSe8Z8ASZ9R1ND1yNCp9eB6WXpnevJ9rVwrK
BCAEHIX5+LFMJj8RsXG4+tz0jzZ668AHa6e5/4lz7KQoeXCSPBHcLf99zIDCArqE2WPxMeZtZBhm
pDe0QcMC8sfzl1eY17Sv2vbxYlbZjlTLfa0okCfM70J/hkCSZblW322udLSr31yKHRyZ5yS1LS5E
542MObMo4wrm0zW522JUV/hejGtdNWsnKvQhAKIjSv0NZ06T+tiBhjnTZq5ECaXipSyt3Cot38G5
x1u+ujWfR3nXynz42S4HDl9jHjxZ/bFLmALeaTFdBOWaEXqhk8h7zbqFNgD5fkoSFEhkAE/xr9P9
0Q8UWPEVVRM8idXdCENxRh10QRZVlNFCxjmk6469VJwyDGIyKphWUiRE4Gaeo4s39qncMnzSpp4B
pIS0y8D/vPTcKX7rqcTTM/WPiQLVXcEduBe1AxbQz5MEeP3NU66o3A31+jEGl5d7n5lH0xbVvm5z
NRwgH/SMjINZ6uuPR4SH7nbamhm//R+eeyPXmzDjGpDFXXU6mvmvu8AWcI233lFuFYgC+hZS3K6y
g0BjMTPR+UyNL7Vd7InSyFETkgcP55aFHrDe2HP5TY+0SyZNkY+IPS0vFK2kIkX0i4unM6u/mASa
/gRqbWeDwJXa5U6Htp20NIs2BMGC+CoS7N1UOkg6cEFq9xW0IdlGMIMWaowdPLtre55qvIakQEjt
B5w6edBTAr6gGmXyxOuLfh7R0mQVGe6Cjy/PNkSp4tzqZSVAoOcV3Oaefono1sR4eTglCRplz9cl
pztIJQopTSceFOFVoZ7qpbBolfVluyzb3SNjBokgXHu2u4/aBxRQt5Ge1QebOQBurg4NKLWayxRp
/sBVrkRAdYEzOoDQ1HUjFhsf/hwp7W19Kpz8VEfosIHsMMu6FnfgW010qN31QaosHF8zvOACcDQ6
tKqlH2K/hUawqwI+MZa/tWIuksgc6z3LKBoY/ped+0sfeE/6vSbZlc94ABYGRCS4PK99thMXc4Hr
j+SfSadwgfQ3m6pIFpJvN51I1EwB6dcKUIi/W21fv9oRq1uPjRp+6cG0AwnH4A6MD+j1oj+cYIMw
AApGY4w7UGFFWbOsTP1Rfs4n4G/ZT92JWn577SAkIcJNHely2dvaQpHJ1j/Rwugj0fS9HC8eQ1h5
opKnJpLaxyodBgycrpEMvEsFpR+1y4uOxYkpONPQnKxgYWv74sSPyE9JITh0UsrGBuUzYvOsRO7O
4nfyN8ww8rkMg5rEKDBwbSytuxnaZopHt8yY/JQxdwfRWH9y2bLRMl5OckANNyG6ta1Jgv+WbVOL
ByiHkaBRYj/2OYPmQnAfrrM5l+zf8EGjH8TJFO2jMRFqBhmkCghj5aVxvDShTM9lnv6DaFC5Iia6
N0b2BPA+akAvNgRRn+DKYv2KwpghrEXhGwVlMxt7adZx25YNaC/1NrH638knd2KgO1LBgdKVon4L
mmY+20nnQqWQFCAAz2KIDJh7KtYt2dNPQZv1Eq+vHSAEiNpV/firG61c92AFE36CCqHZw81CHyYp
GtChQh/9XjhWzPo8GebuHx/DQ9KhdOQDI3g40jhz3uCzTFJbQ2jv31w1/9YP4V97q/rMP3nITZfo
J4LpQHZDrmzJ6lMK1tO8FySeGOQNdt++OeVtyVcEBIhqHDeBp4mAUglVckIGQtfosMjKcSplNHkI
yr8A9Z2HmodPQmvpmPNULRYcNvVq/wchjyMInpk8wz7yYP8EQvKCnKhyxFpwz7TeLSHAAcOMtm7v
2YKgO4LoL8nVHpnQb/5doGd8TnxV8clweUAn6cMwGbQ28NuyFyUeRSBaKQ5dAuXP0AYUVnPqswGG
5jaNIO2did3wgK+2RTVmNhBXmOl5RN3JzLLf+h0vrzk3vJzbj5ti5ntviQx9MBKpkEEOSskVmnzC
9SFkBxs6uvjhXv4xTyOnaJhuUXnQkg4WX7QJJmWyelPIpRQlFzgvhBv09JfDabWyX6qWM90AnS/y
UD/c4hfY+ycVNf4cPo+spTdeN6QwpSwJ3+uSCvYKyxbysYIVP9/QUBDmdFGRoy1sOibqm+e8Pgb/
qkadYJ60+IvJ8fXsbr4Lqsii3gom2L/Pg25sK7h5saykPqL1YDG+HAfJMFozLbN1g9J0Ekn6Bwzo
DSb2O1aqqLgkyikFK5gWP3YgKKjh3qJLBZPLfNwPttV/DJoYf/rKPiMxr5ZR0xviZ/caaky9BI9r
6EL4ATF28N4dxu9MOIWYkq1c3r1Qtx+4oOVQsQUxt1DNFxcVWnjM5v+xNnou5qWpbeEwfFH6yZwa
m/bLbMsJYkmcgXqa2pwcsRTIZCpAs60tfTQAD0q8ZlDR+c3BuSDIROqVrE1qJsrd3DMFMQ8vxwIs
Gvcp1hFKJmSxQXJhQFrypLgYaEl+Zgq9LQtWkH9UysnJkB+d4n1auPXV6UdRFSgmS5IEoIfxOBT1
i5nHvvTgxH1+I6Mf7dqNpg6xol/hDLTiOgxw27IveS8xAxE7Vf6tagKeaED9z8VmKX8eH670wZxF
TsJBMh+fU9OJuINwK8e8aY2DKoiVHnmOCQbb8RvfUj3p+Wgz4XuiECqFvdKhFrxQXAG+A3oyfyRp
j9E9et3valNnoKz4BzvwQztRh6efWjtbJxtOUPSpGos+WaIeOVsLUfRbQuqDkizSBkHBNzIpUck0
Vr06bRQKfvB9HQ1nbPK/pYzn3gFyrK8RUGs/QpmnR87XWCNI2np55Z9bjfZOLlIFOkhcvs9WSxFU
Fpt6eN22H1DMF2TYl3ucJOVLKZ7gi1F+jJvxdb1i0NYDs2pKa+uUDNFZ7k//DMk1Rjfc7efIm71I
n40mVlrKxGWH4LBXY7VG8mBRrfc2JSz04jyp6ReaeH4sExK1mvBl7vBvuyy/H1d1weFlw/HoR6VH
JGmtt+wiRsy0Ak7YW8epZnTKWYHXgykLcvn2opieykMajgoHkETtvaNaiEb/xHqbzUpwRQwWFCLj
Ur6c6r9X5urAJQSvmS8MVVZ/S7WOCtAjsbF74MOYOtg6KQ6Hxp6FTfgWiPu6yv2Qs0upuSpSaOtW
0wqWiR9NwxWKVJwgv9X5LKxnV72VBrygG0vBv7B0wtD/jlquLIDxfj0cofIJsqpttI/GxJFjKc+C
t8INcnH+LURTJdK2rS5eh9F3cLgLkvizQD7LLC1wfxkXq0sZKvRCGOB5U6kSKuRLpYUCOQgkgxjm
HpI6DSMazbCRQK4bGl9TF/4N+JcVNb4QO+pfzfl39nOZcH+9fqkcmtSJZOAjAlgS4ktDV4SrTXJG
xy5H4+EZgF0XWgY3z9XnVfazhxXV+suZDClV6sOPtuglxtsyaKlZYWcIHw1oDbnxjzbXNRGKtYag
iMhZ4XkiNO9CQ/StgMIKUfaObK/4VfS4J+jWnC739+uVEzoZmkBTxxY1fOJHR8E014AXAyBXwpnn
X6vOdCAzUmbPtbivh7GUrk50IYh59qXk/4mHGkAKqgVDqt8DVqh9ytY2hhtNl/8zoP/uxbSoz5WM
ookYzj6eQDN/EXsivFwr+1Ui58qCfzkYwSfV5JyvoGWL7qlCBQCWW/0Wfs/MS5QKo5KytZ6KvF2g
g/wnKwbkGO5f1L7vqwRTHgxE72a3a+t2kg3jZRw161ABSiZDb1JmGNffWPw1nKM0d0UqNT6lPYI7
4jvxTErSq6YVAwP/SKfWKh9DnvQrHNglr5IterdshjCvp5+99YqqXeJn5b/q26CEteY8OuHtikmB
RBoBgXuLgVb5h8Bhu0cN0UnROKpf0rtewVH3oGmttolIC3YdE+XD8ij7w5BoDNS0+tkPQV4BJe2b
tYjTxcPMECxRtGrVg+Poq6bPYLNkEWvyTTuq1BsuHAHeRwuhAWof6ffNWa9v9GNZs80LRfBIrVrn
VXsAGADo9RhI9uqo3ZSj9FVBzUddJJarc9+Udont+EplZixUYK0EnDiENHQjLu6i3BZj6UZ87F82
S2fIwxkFBm03ou1Cn0cRANJZ5eAQOA+aLIGDrq+pMbpjLu8R8sNwIopDKHCm1nhQFT7DwUouDqOw
RYBw+TxuclpRuDzyu2AWLQtcLN+cF+LS2kb2DetMogBaGLfTf9rw2azxR4miNkr1VrfNl6n/sLCu
3ffCcTfTuWs1CSi35VwHBUoQbhIg4UDYmzbHxJaiC76NrO+qdVwTzBhjBsC6u/nt/V4my76wtIdY
H237z3BVZENT9Mt1mPYjC2DYenfmuMfFE4pcK6pn+k2fWHWyWzJym2dYSThD/Wy/LW3tliwAMRbe
5TMFdoXj3KNuplDzFt+VwIK0qHKk7WMaTT/EhbdKf7LEUNKkRBHr/e+ac/AiBkaltspMqPBpJqzO
x444mI9e9fzzfgMLDhDsEXcWtACOhuEy7PHkDSzuYBnISdaI3vQu0qyc0gKG4m3DBDmjMRIodzak
FefztbX3l1bnSBr+D8z2SEs2UWNUIAwl5EEOAbCbHSzD6IpBxbVZiv1iQ8Z1s/AS1yAx/AsZfnPS
+OWYX/SXjRaI63EE711oi3CvR+VKvwUPALDf97jxR2LnilDgMvmMyuwDTW6MzrOG0Fix+KfOCsLi
zp9IzTU3sc3J9ck0RJDfBM9O17g8p5p1G+ARsmKsyFqnYZO4qwtWB1ltXuXPxjC5wgYS5oxwqjHl
HGRIJDEB1zoQKWrxqboX/Lcmwwpq7Nj+j7XrQ6HYw9uXtj2FRtLx86+wYV48dM6wF87jcEyVs0dl
KyRoAiNqbemFTMxW04p2Mr3d2lTwT+BQdYGnI8CIsBl0FhOc0T8yz/OsLOeNY1s/bLvxuzmRjjEJ
CWFYzdDI3y2i11vbgNu4pdSPoSqw7wZ9V2PhxAAu9M0EHw/z3U+rYfq2utoGC0yzYQJeL46mIOZh
A+FESWrkj+Up1DHPcp/Bcg1LZlrC9YB+GAc/CvHtXHOnyAoQ8tYIpCC7v8Qy/6qRicygTha6C+2b
ezSvtiDofYnghCWxerkK+uPC5ocCdEG3lZlFVzuF7Q/kot2z1Y5DDpJDUnvy/5nxsFJZAeox6wle
OqMT6O0NoTtcTmEmgsDr/n63uNzyZCaDpTOsH2b8iPB/jepb0Fp14s34IcNhaeXZWHnpGWDc1o2X
JLu4JgqtpZtbstptMT1BlrzkbSk8a+hF9pRhGrQcGAGgc0gBX5TLy3aKm1aewQnl+vIRdX8eLdxa
x1HPtbYMcUziFX1tKf9AsnBpFjVkaMCA4qNw4fVrP7gMeXslr0iNf7T91+XIQCv8ap7308lmPVDs
ck4hsYv8+VpW49FM8kqEJnUUyZ8vGKoRSV/X3SU99noZ5BPjz3eAk9kyZXeB6nP71gy35jrlVbW/
HNQCQnuWWtQZCpLm5081XlnY1oKgtxGLbd/xhHpDLQ0RryehajyY78BFWfTUYRabHQ+lJqrxQoEh
erjDYRq+zIazQbHzuGH25QmyJ1kHKODnx/qJCTArPmPto6f+kid9OmQgPoJVTgC/JAeta2bml1zI
kIXjwxZhP3A1aYBq7rmYAn5zaFbQEIKWW2c8WxgLJgklEnTToBxp9w3DniZnGheLrV6LPe/dkmof
wST6SLMIzw+5voitkyNNGSWYh479THv5kCP7Ne/+2CpjO2IUwUf3RM6/rJ9ow5CQ4bmBMnhu8W9m
LbK5bT75/Ss5riC81EeOiLb/zgQ/pOF2Um9QAoiyjGhTHVkKnetXvXAK0r/lpMwxU3WVMhxo1Ewp
ixG1HTf1XT8IGJqSMgb6vN6S+jfJz1nzDXuvE7RAJ3iSwMs2obqeKIcs1D7cuDcOuQKjyHlHCsu/
D0BkjhVEbMznjFrf9qfhc2QcLRBickqm3VocVaVhr9UHlbAc4OB+8NcT8FHgZ8mroE+IcpuYxupo
eDaIzWFyyI03CT6SJJyypguw2qejTsBboKmAxPxr9kUXb0ja1xm7YtVjTZBT0GBi2TpWTsSBydLm
n3YMIBDOBlI+A6rMJyGrOqKqu4pS4jG9x+zNVb+GhiUBhkrxNTP5iRmw3RYf1gQx7163gUb1bpzY
LgUmhZfJhp3i94q75CiiknJahvphQY3oQ52wM34ZPS5vBx+XoijjH//NzLyjO67KDAprSDNxUcBa
jMr6kEPOJAJmpQSbK6qRCc4shlIGISLaWDa9jC6qB3vuZ6EO2dd9lVnHrcyJl7V2oo5fbnjsWrEh
FwGdG5hBSfXxBiBw45eJFzGZSKM/sIRJe60kY1KL2z+MA9UKXgYgSR8+hyxZiDCC7WPdwFDSU/4Y
NfhEXFrrwsr6JUugyT7LZSM19TCXSPPzrV98lsEu+BGQf1ovjgr3lXkG+CP6+hFxu7wDmeuBfoyd
+G5d51JeNgWkdI0dw32I5GkXfYCbq4k7rhEWyjrJsCKmGTY43gZt2PQ6fQUUQp6e3qWWu4j+YQPp
KZUsYNElW0pv0A6eJQmGi7zg4xFq7I2YjYHg9kEm1wsEqOs8h/J9eEMcCuA+bufZujuZ9qhnnBZx
1wegVYLoiLWkSHk/q1CP45+IIWgowO87Q/HBDnWGV1VOeOMTye4Bgm+wVA9jU/VCrMUgpKku1cC1
7nbJ7mdEtc92KfceOzeJInSNWxLmg3TulkN+oYlnSGX/VCX39jJc0kH/5HHffpeKWH6hqyjKA9gM
zIvEUc0miPttTknlpMkEzatqveVPXb6Ox9BKlsyZsxYAbLsHO46P5FxdBJPxZk3B5kWI40RnpFZW
z7XrzNxaQP306tjul6TmqqIt9NePyy5DcxV+5DwQgF2T+TxStlTFLlY/+kWFCOOHB4U9NnNhyGFE
2tjvdH6PMUukbKm3BaORikuCLNOCaXlgUQU9UL8XoeQzgxYkBY9tSRKH5s8egVJqF6npkAUlt83L
Ihtwx4tdcwA9HBDiSxBFF8F2FbXw+l6G2iSvuTuWeGz+pn8ZiR0CYMikCHLIwSX2oUmf/Xq46U+n
7vk/FrVd/b6Tsr1WLNtcy8P5zgrKz5D0k9vcHh0zTxfEKiTeN1DT9oRiVGfKZ7tegtskcCiHM0cc
YzPzHbXRMigIzg1ZFJ9WneWG8jfA4cFFjjZJXZEi+cJ1M+380TXcG3cYYuD8NdlGZXvCJJtYQ6cb
lusiO74F7oks1ABgZ/tWt8k9BsCIKGltPQDZQcGDXBapzWIlEeZ8Xffdw9ieocYED2Inudit+7Cr
EWVoPY+AY1z3IGs2ztAOxWlCx3tJxddKsQNFe6cy02TzndRvSPgJRPNKEP2iOq6xNBAjQ7kRor0S
vJNuKMF6WXzI4PpBoVWyL3E40R43w0ID2esjBty1cgWYVJOcodSrUbi22fuh7ClofLHfjSkOFtvl
2EH+6VNg182ert+ve17/wcSP7WJHy/kDHhVWhmsw21gOyYCVXnk/sErt3IU4pUaFEk7YArVkpV2R
k77JuGZgBFVN3OwkFf+F5ZUgdPJTZdOZdu2uUsNlYHE/fkD0mFt3yEkKLh3LefdQLZjs8DItXV6q
KU+aYizAB9gqqIfrtFkR/rcqrbbXkHNuHDgViWA4PZ7A9PhrOZPW+fKN2RdrT5h2KoUNt1TUtMzs
mhUSy+3rD+x60+9u21nfSNi4OoAU2Bq0BVmsiWN8QvzQhvMFAdxJdKGhYeJn//xVIDfvZa1Ws18Q
B+qfkmrTWaZ6ORCRAx3wrhlGHBzesiFQ5sU/LNidgRMHZJj8tRpEuSHQalnKZqYtl2GUIZeF07hH
5WDfUV/YqwCe3c1VyeKPZlpLn8L5MvzYN6zsKEQCg3vKMZotevnqpEhpKDZTZm3aML5uMPIKtNTK
INjx6pkbEz5gVyLEbR6TS/QvF2ocWy9YOBVLIXjEuumlHBYu/rgsfFIdBtOsBH6Ncs9/YlJLahxw
0+ro5R0kcPRKypw6stxmS/dfEmiHxQPR3z4uK2trUJnvMb//dD9lO6ccRapUbXGmJ0vw34CGA81U
YoPNKsOkUaMXZD6RSkqsdGD8a3hDswCBtq7Fllm/WO8Pw7C9ucJ+oQvKoVhO9EGI+M58amKUNRpt
q0BaeQ6BDidTwLOJoqU78VaSVoQVMrWRF/kiVf7jZpbQ1QnIkGH4ZN5wPcJpJ0sU1T9Wat3Q3hei
E/ZSNvCyL+H5hEHw60MsuMvPwKBWbj0ABPMfbLQakDjcZBnOf7zSgn8UFChzUt8xlLZ8OLljn6fp
aL2UIICtevY8W32et9Fhpxk6y8xZ4kP8UkW8j+X1EHnkzaF3GKjdhtIfh3zfsAMA6GJisZBEuN6P
BJEKncDWhD0AN+1Mcy/ppQI/PT70R2qX8dsG/j+O9vHnMjlfUBR18gKjVKGd73Qyff2Z6hZHS9Rc
YqkCZxcTYZ6orNQlqtwuR6XgSVYRHHc/0JOHS14I6FW+MJQFJbqj0kKu6qVqyq5tROUZhrKw3aXb
H5b8AHv26i1GP3QdQozuKR3UiEPGKH5bPirvT80LjTB1lmYGfuouJb9yDpRpsozk0h+N85+be3cF
GCF19hm+82jZLusHDkEoSdMtFkgbH5HsfFwwECvfOpy/mOdN+tEFf9VkE5z7TrEq+k2JaPJJOntn
sFWNtreXU26wArLqihSebZxKRJvG186Sjc+7Rs10JONn9ptdCRc9jjhGD0QMyAB7TWDoqRJP62dP
nGjajpqkOP9R/3upKiti6GRwJWQNYnqn+DIqGLZvavzVQ2xrrBEJ+m2+2g1DC+ZWirNIUkGeS5rx
dpRkTUgmpXidN3tJoY8ATzIR3vBY0wNOtDTK4MYNZhtUnJUZxWa/adWrnrIEq6OhBmhPByIu64le
o4wEZDbL8FEn3Cs55Aais0ogRkmAcgdCBARXRUZRZDBxYI/2DwiJMXYtvSCXmBtsXyhh/nEilAaG
QaKseNe+95X8K+XphJqGJlEFkJ6i6XF+wOVM/GAiJVYKQe7nGHr2qejg+j8bZy9P2iEPJgvqUL9T
39NFg7p4Jt8lkAgg5siQewhYdBESTK5vkOE8XaTo3zJLSNKoXTsqydEQIUGOiEGBxHP/VTWrPnGK
pBiCQB5fVgAvZe4DgeqM2DPgEOX9VCCQd5nQvAUxtMOIvkjsqdsc74MQySj5CPG5YLe3ZTC614wb
odJyYEmr75YVR/RYrW/l8I9YlKjmgUna6eT8Pp20GSk5trw0nrYgnMHK3L9yYC06IxQkCx5X0Am3
wYi8LQ6SxJXZc1qwbkiQy/nVGIVeF4AeYDsctrg7u2XtrNSYL+VjtTnhsUp/LFRS0eKTUiIquqpJ
VwqpDjX+EWe2Rd7WnWG5oTNVzmf8WcnKjLb6an21aT14olDnJiYi6TKXVYTRJaKGMNsHt+n5fS+e
ttXEwMvYgGtRT2lM3h4vWRqyzubxUZe7Q41DhkvnnFO0m0diJ9MlZc5cQqLGo1MzE0FTt/kM+Xlc
KkebB6CmitokAmcMkiBMBddjuLhbvScpXTs3g4guOmxD50RxpWFKrSujVwM9qswyw9MquhHPpv3v
ks+FXNHjzcD0xsgSiPAoRkLx8YEK6FYslmByHoDPwN+MEQ0XhPIBpkrJY+7R6hAKgFjAADzAb3KE
B+lqOp3WVkMJBgvMaZZVKKKeCqyi78JvH3BorcVylrPFFviepyHRjYF5IZeNoPF4jtJ8ksxFOap2
hUdbPAt3pYVDxcQ/dYcT/N/CD9CwsAOk5X7zpzWF+83tY9/rye57KPA7IkU3DeJtl8XnaaVzS5T1
E/jX+4Li4w43x8LzdGSwEmDX/Dyw8T4A+dvox/U38WYg/RQPHIngXiRFfDu580E5xsZ72uFsjpE4
+tdEkGjDxQQqtpHxRiJBibenOTkSlxwgBYBMuf2p1NG7l4SLRsSN3/lPT/a+EAXIhH6Gc8Xw77uC
kfo2s4hSPeT2T0e9BAS53z7H+pl2dnTqesOhB1rNZ8PDuMFw1xSHunw0rhu+jz0b7FEDRDCVHXG8
tIIygmJMHaXhTG611y4nUMjLHv4pkaQLeiWZEE+H2sTstSslAAP2uJkZqxMXh3sM2la9g4qda44b
u0mNqGDU9vJy385O9QPbgdadCWM+n3Q6ULioNd7K4aSc1R25ORe9Rin0SP9RLNB2WWPOo9Kpazn6
3J7GdQ9fWIAZWfTF7bkn4kA4/2iXMylPlfkmIdLvHOPkCuZNrBiocegHEH5qjrx74Xbm/PmQix67
HqLiass1VzB9HI8xCiZ5MGc9yLxgMHDuBKMP6lTTqoHQ+UquLUZixeZ0c4KvYpp0a0xejfufGHsl
ArQ/Y7blAPrDAmShJikswUDm0wX+gpm6d+FbGt+lVcB4QWFfwXiFJ8s/iEJue33vkjJ0maN5Ebrv
KNjHVP3pcNIS0a1SwLEIRu6IvV/nqQodzSB+52c9fsFHYkEmkUlraWMWWE0EVHK1/fiGJTm5/BhY
jnmhJUx5TiyZw4hfIhxGOHtd5axrLgPfZwkPyWkM/T2aSQBxxxvIJD+1niDOcgebe/l20nXazvjL
I3j3ItwiRGM8c5MMJAF/c2ieCkTybQNodDzY11F2YjRyTm3yM1sYaDAziprKXjr5B7jim3avW18n
ZnLArlzzA/W0pfz2qPppRbHskpTTiyC4iovhbZn3HMf71//JoqtBe1Hz5clx6nq6qNaGhfISQzV1
hygJPYAzR0Lw3KOziYL8aBL6myfE+/rFdvvYjbvmDnWiNA23IVUXEvWNTmJ8RPNDYkEdwIi+4+Wg
D3hSL7rOzt91JnVTsdY5p1K9yosr5JWxDClrbMCzbCe2plTTyrueKcgPq6OBsumyp5KCXicHix2U
U4FoJotKQ8OzN0RxQym3fnp4O6b9bslaZrSH3z9cy+JJPVaB8KdekG1El+3aenls3LnOR4pHR3Fm
zAzDXuSJ+43dEa/wcEMQVtPSStbHXR3ynvf8wt44abL5QXRMuR9E0qbYcjVtxJLgDjHC31Oh/GhN
V908+uL9+1xsL25geRY+0R8IkmR9PQDmjdObGMPvRA/siHPtnlNaN7ggtaosX6kzZM3dt6snW6Mw
n/FfdmOzrZDgC7Azh4Gh9btGPAX+oORgVTXZzYMrfYcE6Q9+fxLD09LpjsvA0hf8TWkMKYp32VN7
kmX09daHDXDoYmTZoq8wtEQsqNYDxnMBQC3Lb3n2AnbYk1+yyR2OXlU7N4pCmRQmbSzJPIeSZ03K
oM9A29yDnexsX9ZVhGTGYhLEuyerisLHL+ZPTt6m3PzvRrb4UHDpOFd37fCoutXxwsESFqPKeg0k
HYnW1S5aXjpNbSblG9ah+iKrviP+NzUQUksr94t16zu77W2SzF8OfMa1DKiUBubPCWHnT7E1GNQf
ovnIygFPOomTQnS6BfeGILl3De/uQsjUNBB3k/l9MWfBaaB90lw/UavwAGqCYwoBmdVmftqId0ok
hi7KC4vNXVG6+3/QhUZYAICpmMDNqUYyE4AVWsUZrdZ69l1/nfbFjeHioMyrYSoOWI6v2y/KU6ll
ygbRqyfTcJV7iYTkbQRWJ2cxyG2gYfI9V0RaAtpTkaDKWRLtG+cHpttckUjBQ82iuDWYWdVWiAO+
9V6P7eX7Ov/sLS4C30yYCOWskwfM7kGQImepL4dgMWm1DnzS7IcnWMl0GelmTekMjyLQUTxwvFWZ
0LpO8zcJ0fpR4Ik5CoIJgHQiYcaH8zlyXg2ILVX/nbqgSfrpM7SOYsAmUY5RyVCG2s+pKHPD1x+W
JchkOSqEl/GAr0/yMfcA79uuDiLvVACFWQxj2cwkk2KJ9I3VIiWax7ZSKo6wzQwrso7FRBG1VljR
93/WqdOPJO5B+UEjF9roBssi1drypGDxQWo7/fT9hxTTNHGTD0EopDmPsVSknovp51zrr6p1VydP
2iNlUGzny8XppG3yG+FkVaRiIH0vohUbzdvhFA51rMQFv47FO8hLGToyxdIe4Sc58JyAMO3k9STh
tfXAiUIW+PCilTNaahcx70jOo0WYi5iFQebavFopPzr7WFu1/adjRfrK2PTMy+kH+8ItHsbhgYlZ
XbHRywEIHlyjlm0x20w2G8dqJVvjpV6dlXZ9TIEmmUgYf8up0NrBe5ZMDxBGgk8bT1SE77WGpk54
Ijb4ZquRVX7NUHAf0xFRHMgZIUrEiD515+PaTWzGx8Vc5OoaeH2ixH8tNHcVtWahqCZ1tXVF9jmE
B8wZ7se8mKRFu2HfSknf0U6x8Ozf1D2Yo4GfIbzQSc2SK+1Z1wnhScPc+ScDe3Bc8h98dngCtNvH
mzO27FETnO36Tnp/uS7Qgx9Zy1EJMvjn0XFCactEStXnlnqhYYvCa3gLc3KPgpLF7Kx+2wK39z+X
drF1t4DxHdB1JpmpmQOEqxgC18Svs2RBWLmrJkorb7+HhnaGaZDbAoeLpvLnz18LnparSikT7jdS
/u7FUM1UQefpmWda0Sa24ftuBCt9PCMAWOPP7/UIxmZvM++EP4XvS+XozMaZI9v/Xi52t9y27mvT
IBIanC/OjdPpBsKB4t81RQ81N7NtcYBa/91ePbz/LN52urM6AgkNckxc70TGPXQSnuX5tDH101Ok
pKsI+YoQuwH7oJOAGA8yOZ5ENWHz+cyl2cY4tkIpAbTS2itPeOU/56kiappx5pKJkLCh1n91I8Nz
7hypYtAwL8pguJQsaP8sS4GS2QMGJZOLT1xCtch9p3+94NYj+zea9E2E1IY0N5/s3vj7pdcrsMDs
D3TkixJw3lhgegP9xNyN4OFt84N+E5+FWeAIgUXM9u7/HXJuxiOfJKLy0eDaFJX0eOxALZZJZ22L
8755nnXavQWC1QDi4yOejNUr6fBxXRM1E60UVdggD5/isdQOl2B9GlDv7ACex/5utwLLdCii1YWT
BH8k4W4aQfRzqYX1tGfUEPpSEhDx/hXfKLP494pv5Pdxl5gHwgSB322Kc86nDhn99+89J8u36+Rw
AX9rgjAQ6KJHPznP3p5DDHhpKRqvflmyvuZHdOszIecv125pcSFuco9739frMOFicaV2iBQ6qafB
Q1/kCuCciLBuGOZkJU7iqNwIG2RRv/pRMsJW22kFoHPmcAtjVkEjGCC4EanXq/JmfF3T1EcBa8Xo
azpHlMhZJCEnXRSvHQ+MvBoMC3HJgO4kOVyy2E3W0EzSUuW5A4y8NjZKOMsxepDprm2WZdgnTqHi
34rCmISvhFbvVw4TUSMSXCK3ofO79UOQjsK31vRpt+6+wiquCUeN/ZawZFdcOX48oe89LPjgkp0N
M6Z0LBYHEjqfp2w3vWhgz50N6ZMUnZprXSu6ZZp1TgNHRFgLTcK6vkb/S9a2VT7jsPosyWpf+trn
X1gIcESVUyFZE/j1GGqA4I0B/iMNgs7nxgiToiXc7tJik1/vjyabD4CoRiJ8FbJSK129FHiTUUxW
MoNkT+CUkSqCpZf08ZNB4936nWHwqS9vgmEG+k28MHeQmkrzP/d6V9kBLIEWQIPrgmnZoNUR38RU
YlaNf6hdXOLaNlvMjEsCnynUGz1Nv3Lo+Em4EzuR2TTzQUilshnC5vJ1unnlr4VXMEDoWBduVAOw
uwAOpNp1BO9Yu27K5NpbWyytz3JaXUyE91xgOgZx1Q5n8Rqp719mu7Whh2rp86HvyP/LwE7RlmZs
Q8KdPrzkZiF1bv/fG1tzjNrBPNa7q1dFJoaXUBMO0Nj3JfpCddbNLhxOkDNi7rt+VZ94Mi2VBNok
uj42SKkfhOJ943dQhyAwiiqSkctj8lFt46a1pLWEB5xFa6DcXeIJWft0iqEg6/AHSVwJMSpMYzOB
Y7H/dl+5hWFUBRBLGx6mUaZ4CT8q7Vw1f4pvvhDRdhOmiREwvCCtY0lazBUBKkVl7dn2jjsq8kaF
lEQKBArc1HeMwxcskbncseRf1UyFNpiKUuaRj2nAw9FSvgiqvVjo7zdOgp2LxrX33+8DsvTU4nCt
IGf6+vRSfXOwVeJUvs0+mLBM00NZFHFIUiV1RePuLdvS1iSdOm2wbx7IvsUiY9j+Ej030Y6XJyUT
hQuDXj8O0LTom3lElzIz9RyDH59lHvnX4t5Hrgyr//mXn89wvrAFBExI0uAs1kqihCdv4L1+J5Ok
2craNslY9lrUhQyrq3E5ZUqeWQK0DR9+8pJwsq7zKads2sqDG9lH65N35sHqSGvMClq7aFJqCZQr
JOZfW0uQWs7jKMO1n6BJVwLxPKwMp7y2mB7oMm3M+0cQw/NRiqFdl7L1pVmtS3wiuFAUDeb2TDdZ
MDhsl6ZRMfMKg21ls/ARbFbn8S3PUNG8Ptbo1YUVJq9IJ5TZ5p+r5c+ZUqMd+8Aa4j9Liu/QFemT
2BhgYY0cmWHbiEpXX8zDqL8KwjysktH3kS3SOSyQUqvgaFKdoWDeGK5R/O3tRV65JWE5aQxC8qC3
GPoO/ZgUvjlIHO9xg0bpR0Bu2NpUzGsARLjthhtC+OFHeqCrqHQwz3KmarYW9IwPzUIp2wzZXSQv
UzUdQIJREmoXYYOTFG5DAABbWCBuzrEyQFruzLSOXl0VikBSAL400Iyfq7o7iaq+w/oGFTj0Ar1F
xNy3j7rAmkcgjSDtjj8bI96pUdidbSYgcxGWdgRmX+knd3AjlW89teSPV3GLHROdZlL4XqhOXKH4
F0i2hUJtQGzNnTi3Dg0RAEdYPW4Bp2eAancGiz7h0OnQ06zVrjNg5IGZOQAta7lIkHnDI/QO0elF
jnioIZegqkUWECZsHP+DoRyavDsvhjf+yNZK9QWcoso1dSh25ekHfWYODlP/ZzD2FFaND4QOWfGV
FTxDMpEn7BVIU+oz6KKhZ5seJCjb3qZVdTB+e8Qj62/+4LMB41TwP41RngvsvP5Q3NvpgW6LC0mw
NnZTUcUWn9Dm/1W9noe8uBgRyNOvUDmCj40QbtVClYo66SGKGq+oTQv7nV5n+CxseRcPMvLsS4N/
s3CVWXYRYi8oKt3LooY9Ha7ZO8RQAPRlmKYHIyaVCrMdvl1yHPP4PnMobJNwq6W6LMbHoXVNDmFc
0HMcrUGRjJS1CwHcRgV3o6Hh029lYIYFd3nqhFdNOZ6B3m86jjyVQmJXy+2RtP9cTRoDsd/dfiSo
5FWHTdlKoU+nHW7CluOke5pzSKPKV7n9HfGtmuYUCy7yyXKm2nLFKRsUiZq149Z1ptyodYtvVr8S
fOL9C1q+MaPKoFgRpXVgYxP6X5y7l3i8SfHQ3lWJJLZSRS43E2i+XYgZeBaKctKj6D/XfjUDhRQZ
lYpFf3nbbjjDg17evu3znCQvfT4cDy5OZaEe9nzkt+riMpiFoTu0f+L04XDr1D+9r5/Bj18yFAt7
AfzR1XIQrCJXbUV+vq+n/ffNrIcBrhGUHz3oPcTgMN8ViFGfYYSG37QvOjkNWBocsp1cwbTuG636
7GLLQD+KvbKhYJ74k9adQ4IQ6BpUZtKgLkKzrVkJNIpDzvXpF8ELQZDHYyG32cFJB1J1Zcgf+IUZ
Y0+bJIyYwaSaXD99XHpULhiPcN/c/fHsTHd8svACL6X+RbKd5+Xya7SmYZdSyLyc9Dk0K4Voko7v
PaSqOYgrh41BF9wcq0aLEo7mkoA6PWBBvkmbN9yVCuQ9Lfa+BcTZoKtKrqezM4EOMgL6cJiT9W++
rHJMIMTW9wdtGracMUmLMDQJHJdvlFa5yfeTWXr8Y5tdw9beWbXhSfwbISZVOejKuIyzYhSR3z1S
B+nStLw/zv4Ct56TJI/UWbdno8lwVtG0wD4XzLb7ig9iWxNe64tUq+6Fc5sWjNxSUlh4H/q1qOyE
yL641narmlus4iApb/dSUo2uYAbKiU9pU7ElOH4lm7KzDDI82k8UXKqeldWjLQMFUGSMpZbZKDpQ
ZXHnXGqbAPhu9dPlLxxjx+STgQ03x3CMgD1PnANAQLbud6aDA9siqqCw2/6uuIa2BlOQp5YGRohL
3ySYPg10KuhNEWW5ElUKoyxV4qQP7o9DFF4IQulS4pJ2f7ykecWpij00LNw5+IQ10avOSqXkCjZi
lvLkoW1ik8NU3E+QRDBqZqa/k3tkann4g/ywk/fRpfo4VLY58KKcYbYmaDptnWrh6F/Gsv3qXK9G
bjRGl0C6A/O1RnfE+jSi9kjCGMWH7dkupC9D7Jd35djMQeMDXHASZ8lYpoWx/WGlgy/jts/WCP5W
IoWJcPDy2m5+WbCcPBEV6HpYEtjze1WpDSWpEZ45w+SnUHpiOFu45V3ZHbTgpXLcMICUgzqscdTN
vI0mMuYqIZDxn8ezHVx+wAgpepcYiqpUbIyjD4CK6K9WHp9W4Sj7FAEXZo27CINh+T+lseSt9VMz
qD9TjBxJXxGwwZUkXp73USk3mssrttY7C1Qvlp3fbwUZHWU4jYWbjFQYp/31ujlxTEtL5Y3BTwuO
1WOz2mP2rBOb7FytCb/wCSbSveVLJe6ydD+kOAoRS3Ha5iC2KyV0SAVdCeNLmOBQopmWxQWfp8gD
U/IZ4SDRbKoeCuQ5WykUezYTwsZRhXBQiNdkvzoHhOybfyubMu0JaeWelNh3V41cLZluBrAixCRw
PQ9As2TEpvlnUCvlASXmagjco2navoPmAqL71LTus2e42rRU3H3vfLh5Ig8176cS7bgIeZ60Qjsj
dKZ9tpmb4EAPHxGsZ6vH5+wR/IMKdwV/hc26Tl/QcXrtCHhcYMHKELEPISoSjVKuDz9TpYYzUZ9B
FtadFWy9mkvYmIxlvOPuhY1rhyUlEsHq746Y8SZf3hz2/9kOEuoFinPHRxsdagwHSBguEGX/YVv3
5LSYFWG8IRScCDht88BOAMENZx/OK7OlTSgHNEQtT5vjdg6OuvyiS5mP7mwlzM+CvTytjbwlNr6f
lz59dsOqiP97nF2rakKs6+BOWp0YOs1OlTardZxehQ/UQbFivStrk1zgoOOvn53+QYW/fVg9RdKX
XiY27Oav6JNLg7qsSIs4uqyTWdZhOPApQRw9JIocbfsx3BSRoZo38DTZ5WRjSPcF6leX08DmJIcA
FXYxE2KgaY/RqLkRQJk1yAsJ2LIiCHj/K5a1LAqXgA+FADy5OekMnf6Dr2pTjIYOJvLb9fbLUG72
L6aL4XR01Jz6jf0YwY/xLmWG04Rd58qup8Bf7/fpFxV7O8NbgCcopEj/1wr+GsfFhS+3grwLdTiI
j6atf59mXMBjHnL6Fbiu8GIP/LNy9J2aR5+fIA2Xr2lQhDmuWVAMlkn8hBbXsjhmgexaImoKsoby
ceJrodSXNqggQCOEdan+PIppKquaZLCpfMWkCvg5ZgGGPoDLltfTo8rVatMbWoKsnNgCK9mB+Gbz
6WLBNWdsojgA5AjaZ2/WI/Fad1R9S9E3Av6gVWfYziruPvaFxm3vxDGcdxDs6XzHmQkwYOL3xasL
cbbNUyDgFywrrKrDpBIm50ubEgiWaW2MUFJBLanKKHGTchAZYa/f1IzxGZ83bXS/V3qDoYzEuoZJ
gsfIMdAHhspe4KhD/nhCUHvSU8k0fZ6AS/8CqFIM59t/9SWokmdZx4+fjQ3TQp0Q1l0vPdcPb1an
WoL7wcGMQY0IG7uqK6lJV7g3ZaqU2m9DCBRoYh8X48QoZ615+QiUvIhYrGTXBxz6CjNer9cZ/v+F
P3ZuCmoSf1gnZGVRP+t2j3xjv6oMtVJIlf4kf2M6aHDvHXp2cjBUivsgR4O/tC2sUac8e5At4Z3s
HXLYtdN5KlJ3IHdq5qAks+ImY5quRNHSwl10M66/82TQ76LJevyYHgg65wKHThHim0MiY5WV53Pi
ip5kRVjYiaAhW6+BPeb//1DoKatF/IVhVO9vb0E40xsQP5RSGXVxYuLV5k8TxPOyZQFPYt0qdC58
X2pYBWh06uUs/V86OO8TKndTSUPpvCfmyGeDI147goVt1ndO+ir87VIU7hjr+7l2WQP49o6EVWhs
Drycc+nXrU6FurkI9pGc1e+Mxnjv1HUHtjK6jsfOpVrq2PqdODN+esFZsBbyXQheBBMSQQupj5xt
CVi1Utc2flTJEtu1pp74ZEDSNiATZzKWIs7XP4wZLEG3Q3swseawlcGnijnaJJJgcZdhFybVuLK7
IpD6SBfBNiDLsLWY3FnjUOKraGxQd53A2lDwiTvngQKGpuPkcjFFHoK3R4V2SDFXSujS9nBIw1cO
fyZXHVWN26k/+ZHscWi3uHdaJnDYdDmEdeG2dYa8PoeUNwikEs/F0Opu5CUjHLLdVok39Lg+0tyo
k7K5HBD4L5RpVDhKbPz6Qx2arbHM2b6BogZ2EpgpyfTKkSRTPpO9Lu14UwXqHElUk5z5E2O/VA7V
WxmSlyicetlDtgNbm4hrT26ePDZYhm/gCiql0JCQFyz8S4WyGGt2mmNP7aCtmfmXZhK7/EDea0H8
dhKnRwQPZj7hHwT+6cRV3ptE4eEERrvIKN8TazfPVzOejoEz70bg6/wDprK+GnVy8HV7FQhv9ITS
moeZVkUVqwWQXAbwyI/4/RpWH3y+aKy7qIuO4XJGNRjFUZ0x6Lh+iblG4UTAQcAGPpo+iwl/8YVu
zfwSOF9r/HISkQ2bcMLVQKJV+L51jomLbiMgCpq5b8JMnIoYHf0CoSmUqayonfdmAdTg3RYyfhLx
tfAFVFsWwJX29jlS0ASWGUkltQ/uzuUkCikkplwTIsF0qaMicPahFCMZN2LUZaq4ngrvfNzbahS9
jaERgUHnsTqYUekrantjwQEU6J29jz5/Q2omFYBMmfgKP/FfdvbNvCLQmiGSDMAcXELLK6qnVcx7
TkbUeHE0l1Ije5TWsZjP+LY1cIutDwIlxyqLrAXmgLCsLy6B5x2F74uu+xcbsTYgzYO3htrWwwoc
1KK6jpIGZEJfKlpMgeWbpntELImMFqynppeKgNsAIp6C2b78vKXasuJIf4pBh94uricYFeiOBMpV
jorlPlF6aZmf5yfqqfqlzb1mk0l5XkkSCZmYVNIEKIR77gJM55T9sNL2Gt2n2SVfNZdfGhBmRMqD
xTKGJun23oI+EKXxQwg8tXvk6dJIpOZc1pUlenNj1doj9+NctFtOEHN4ywmTJRx9BJZZ7fqdovt/
ShZN5FAmLbM/AMrd8AH20fmS3Ii8BABsFYLoQ3Y6fELdFX1OB2oMoimUBIAGMy7YYS+T0fCHbffx
T4etKKVgPv7neEDnn0AiRrRhEBOFIjXTdNPuNZ1vDrJNwFuc1w71gKitWpmO4GNV35Vrm1AZ0o3/
aZuiKjWxGrQEDrTqnwz9MJCJ3CQoo2mH3qdpLP8NgbsehG78DnYNBkiwGIE35pinA3w6kx3ogj7G
lZqzBgDtu7hiNCAVzcrrgKdlUMdNFGFnJeS7GCot9gOfaem0Hzt0bfkKbsl1Li4f5iVwMPGhmRlr
WhJy263bqFCdiDkpOcD4Gu5mG3nHq++vVdYlcuPuF2d8PvK90yuUxRjBhKQFrLhRd0NaX9QHJD4J
pb0A9yBGaRIv9RNjSM3gJ+FF6kNaWgBA8Vod1Qx1DHkcwgn1Xa1bFBgWJCo9iZL6fWdntxqpYcrR
ckCljVvk5BKer9D5qehroKc57jecJOAKjX7I6lLABbzkEN/+YzFCaZVj6VPCh8AMzw17Z67AvHDJ
+qHhdn0/q7VxqroEsA77huUjLZcE/c9fHLaLKmuNcUACg0IiyECfkNjCfGCf9nF0fMEsNT1LTxNZ
ksGozr5kp4pkH5p1jl8xVlzTdWYfq7gq47AklGTrQTm4kmMD8B8UabqC9rJ1+wZapIPV1GcwQmYy
4y3fA09k7GJmOjZ+XcqvHeVk/U3tx6TMKsGey8jldBmApCacV15wGNWID4XzRJXGTFP1Jq6YFefb
j5AH6Bt0wBDOojQt11ynJGpAnsLw6Bkm6hn9pRnjRGdVg9sM198ZfCyab7LNRQKLsAcdVDJVTnfP
OAQIC9HWQ77Qpkt+L6Sim0hmLfV2umiumfA+mazuYXUkrsxPUxRBIwdZ7Bfj0sJ24A8pXNnbUV7V
hEH1UAW6ZNpGmAtQ4JRhvP+q5oXdZlBTiXJ0qLeE/9H9AjUQBx55MWW2F5jkdSz7qYzRpwvJnK/f
6WwM9bfbBMLBe1m81QtbSI/UP+hOKj5LVHHpObxovZ+V/I57ErHf8hExE31EW7FbWL/Wv6s1nShE
EQJyHp91TRXLqdA906jFX0iij83VHUcGJ0KKbMi/JiJeWi3+a+qUfyeLGpfB8aPDNi2ugpnFDA7u
DoX9a0YZ0vnG08opRseotxELOTAQ9NFEAztcus35b9paDQjTMyBcvtZo8c7czvBHfL1PCVruD3s1
7o7Z5TxlRvGEoixBQUdxE2GFn4Ng+irf8Sd7GFzDavtwcNRB1xtEeeM1ZYm89UH7WNqRbNHESsCI
ArXwGJgfK6OqOB9K55DyNMEdx6QcAOdSw265mpHl47Vv/ZCjCK6w0t66XxxzPK5kaIiwW1HE56Vp
1FgCUmTZVBfy91Tq8NzOnNzd2V9Rmf/Ppp4k54rsid2crVhc4n1MdzHEK2uEKl48XcV3r61a9p68
LPIKQGSTumCVC9mk2xSpNQylnGkiaotHdadz7vxx7ee35lBPiIWNeaOYtgtJLl8uVwlt3kzldLOW
ADeyWtasqQ4eosM2C3vNYSJfK+oAQrny90U1Gi3WdEGOHt3nji6kuGmNGmNGER6ALq4gsdpv089m
TCHIm6XxKWi3OmcWn+W8bJH7ngr7MJN7RZAUs0XIg3eKRwJRUPq2rKjONy2J0xcr+aQm1qldinfF
wS+s3SXtTCR/yqXdYM9kleY3FGjjvvn/wZoBZEL9UWk/Don6cfPQ6SgFzXCzFHsiU6/ho+Rb5RvF
0G6bWPlwiD8KDb2fHPGur1G/z3wbjm0lCU2v/OjbMbkMTe9Ur8Yyb3rNmqEYO5qN3zpLZUfr1jN1
1YPhAvuDQutzLIHB5YF/5kChbqAEx22HIRnIqc0j/4w0CxICQXyw0pW3SXI2QJzXgmxaZblf2QM9
/ahjb6og2hB91u8L6qzc3r9gKHam7+InACiWo2Q5cz8p1FoTCiTGf3u31IctmZSRl92rE5YNrgaJ
pKEqcBHVRpO8pSLPm+a7vBUMkiw5ZQ8xcBnbfjBF97e3lM7+jZBT8hQI0ZJcKjXhDu13wWlHvBUK
MoFpGS3aaWp9K7whI+34X3LYVWIgkwXLNEW/iqmkkcVNdpgl1IJwGGAbuWYocBYgs6eYSxNYQEhG
F06gSfaYzpRR5CylZUcUFNT1mloODrOeoC0htTNhLuae+4kLGYzELRENPSETcexWD+THZo/IUxmq
ujw7+tKQbgrDFT/16CINwXJxntYQrZILVzl+3PCH8WVDQoO1uLjjrzkjnpz9o61tZUcXIGjJVzSO
8Imd4lHZdvJmp0Y1iW5XnOh5/DS46noM1ebaQsq0TpDGbe8sHtzdOBJSUwevhpgCfAAmLz7KoEfD
EL8S0H5MDcSBJHi7zIni0/bQqb/x7DJh7hRKWM4/qf/J7Hwt6IsDfAHWV8qKKHeb3S9caMAj6BQQ
Q4meGwpYCacgc/JYM1sQUcnLZfWVJwUPH1bHhtwSVxx/ioam1cC/nLuAIC6ixzqPiFx7KPfIRyxM
rf43oJm513Oxby0BduPr01szyTyrzo6NTvkhv7BDXE97zEUibhORJQFdkBh3f0hXc2q3CRC6wBzh
DYOzywYGf3bd2G89ttCh2lgOHmvY+gGW4TYQmpa5qhDfW/aSDqDV2YYR9I0HLSTgHQhO6JXJ/okz
8kT4mMUYp9C0jZTFS1iQPX3TxyzE6pzlEBWdg8siW7DpF/Ck85/PYjYfP2gYtOsPgYcnN5QaRqzE
N/2d8SH1I4Yd1dG+GHuJ1zW7tnsX2paclSDmSNQYSqXpzKM+NAcJg8lcL3BvjEq74Gz6HvYwd7lR
KKY/OhJYIGY9U1USd3tRR4UWP1lPmc8SWDlwMwONxUFA5umr/glDTWraZhP4pSbTk+VVayhkOnve
rlys8YciEOVx3iY8nhqLd0gbtKMZZD4qx613eOeC5ilLG1QOiaeAt3nz+N2mh2oCxa4lXVWJkdqw
r0S9ULPDop5139AdoCQtiBIcSXIy3sF3dAMyyMoDZsNbte6L1BPLvoBbcHYxF3J/DK4fGmLhU7HV
8vZ1L+moYASXy1ieZziTL0kwOgjlRnKEQ/Fe3AKMezX5F+VhAxpLCaK9kjiUBqzqFBao/m50sPZv
mLgjCnQO5bQ/dlOsjXrn67wkC/GjVWSj6eRhxe6lTGxY6QWUpYQzL6MkXrnWIm+JY0gpLZuHZt6M
KHIxLLTQW2fUOw3Y+SEJ8QmoH4Y6kG6R6NvCCje8VSS6+NMZ8jd7CwZx0cUyacnbpC/RXJd/187Y
1giyux0etIu3YqRExo9SU6FNvYSUbL7IHouE5senOlfApzwxoPsS6RsOxCijdCoGgAjoFsthDGFP
cBrGGahC+uALSML6RklgiOeZw8H3zm3HKVd1CybQgnuj/eBNDMHVJwQSCc6Em8wCfXwQwokq3Rib
/2AHMnSes+rOQ9L4dJU+Q+wOYqUBGcI1KrCVebNPEdEcDZ9Dn6Jg4hs5asYk/1QQsxhsYeV0ktLl
aAsusnS2MARbCQBvCG8pqZ57K34MpiDrlHCVARI+Bxw3e8JBuaknnx0NqEFzylvr6QnXsbu2+emI
rR4wvi15nwfByfAgvqfJ7jAXK62hHdkGVntqSaJoZbGXnSG/xYZESMPgZlALXHoIUa8IULYeyLxv
WsJeb74HBJJa9BRflpnGmUVr3brh3jWgdUcdHOmYoOiQdcmXxcEMqYstWsVZ5peIicVHRHA/PUT6
cAz7VoDtGON7HJ+EgmST/boIVOi3SAZj3G1ZFeTJ6VAXuPVcX0m25HNp6LWi18dbq/GsyS1o4754
eNeQt1zJCraQ1evHmdF9Jg4gwRUE94j70ttJ8i24afgFmneTDN+UIvKDsRJDVKY2T7ht+3fWQHv9
2f+UJBeAvDaWhjuOD8WKxnoRdHW8CueZMeA4UMIbnxovKJqvwpI5Uh8aKMlVTihflxaw+nPqnu5G
XEiEZkdwj7+U3RFHf2uVoFtSvPNCa5qpCZsFB1IVRUuSGzZrP1sB769wblkZH7tlFL6kYLpToqER
a8ela6JHPubUVVIfsg3X7gxQtXyA8zi5mO4oQsfxlS/z9G9OvLtCPEU1xMyblKKO7fwtIKTRFf9M
EIc4tuK22Xd8RLfCk0SkQmnu1G3wbZ89xP29ditWrtbeF4N69eRyvN0+2ST2q1rqhSZtmJ9VVqQC
E2JraxHuGZvqwIwPmWBlGl+tqV4P57h8ljBMzjwA0mq+/blR/1/zSWp0pB/iOp0cWJLrHsSI9gab
1hentevjj2CI6htFhNIj0Xiyad8/bIXMFAnS/l8w1dtbGCJ+cTErtLeXBpJD21F/T+PrbGSMmBNl
RAn7/9MBN5+JWUlgVJ/feXOlVxEg257PixMe4FHVCwoHof8yds4OLicYRh/keO3EEKwSrTlfWMzj
OeyKI4g2XulIdp+oS2zIo7yhmMrevvWd4P60s+3DdtQ2FHfwhxPB9WP66gse4tbBVM9Ht79vhAGu
AdpRvi/NgC4PWrfaFTrXHdF2XQawUchQw8h2zcSxCvIiSc4w3DyVOtoG115Vlj4dnMjZDF1nmpE+
LZuPuTzilhrMbdnrDvuLIy3jICV621q74Y9ZZCVS8VRp75/8tNKhohGTqyiwDIXd3v4qjX0P2d2T
Fs9u/Z8wZF8Qbijs5A/+RZ39xiSHIznV6+lDJFPXWu7Tm811C+AxUYQlGL44RUFiu0WX91U/SyRZ
FItSEDP9Phbzz15zeFDiuSvPuWKWQM5lqzkfJKh4jjXspGtVZAJIoVvOtguzop+qpmrdSy+Gdfa5
D7WNJIfMHWYtlRpkHJagYA7NXgV/HOm65+o37gbHwZ7naq6I5QzCqoRd4XtyxxTpMGVDPetIME7P
m2icYVH0Vk9zCU2sP6qtVMtJBhHaQ13afcYWfJpoAkn0rjfuqE6svf2YCQfk+v/Y7cWwt8vyoZQ0
F6wMZIqeTbNTdkUWaLzBx9xeQa7eK8/pDPnu7gV4J9ApxP/qEJI8dq5mSd3AMYIDlwzwavWpBuSW
Z9mJPYYXur2RkG4T3Fu0c9ktwCsDo4jGhvUwzdfBuR3PIxOL8PMyV5Vi33O3/Nd0+iM4BPYnr0Ib
Rhfdi3S1ERjM2biu1TenTbN/Yto8twHRenabEUxBY/xJzmrbPbk3UkktT1y3RyXBkW6GKBd2jW5k
Gj1K1w63V6tl44vq9TIo8OyyPY6C6jS9yAmsTj+nCPiYZGpNJX6GiF+oCI0MmDqBHt77AVilyZzU
PClZsaJ5+b4zUACpRmHOuM9F0hfe4WVohrJBwfy8FPaE3X4EVs0ESmS90TM9/vdgANjyvo1a0zAy
vmKLuin38c+duaNPCiLoMmZL6pm8L8CIwvnhNj2Qne0aA19RQncZtJFuXOaO08haQkESGyO+QfDU
sQRdrTovPGeTXhzGnDAeDLpFx7n+puU8BNxuCZ2IfcwX7ubRiQM0d1bvUEId7X2TYquxqZnQ9L1h
S2rW3AGbIh9ZMG5jEfMX10LJ28cK00XquT1WpxnOKWD1jXoAvS+KmHxSwZnrfsBFqyEkWxXESa0I
RYugp9AFrJHTCDdNNrVT70U9B3XEMdCaX23E2TFmV/WE9NW5LzHjHdcy3OmlgORIMC6tARNVXhiY
fxQI7pMAqN/4fYftuORm7F2kl4kQcNRAS8XpZzTa/ICvmB5MP4zMfBn/7825abLdoQYMm7Nh7ZdM
qcXnVQ6O0RUslNSGvdMc0IErWNkZXTTmvMopQ5NUgfkyPxDsqTRiNw2ikZBxhf/j96BtgOtan9W9
FZPXN6V76/Ruilw1Dts4T4ir+MC9/sNhePXaTzPzFL8IxvkkvH1y+2qxD2rIsLRF4er44WwNNcl+
DsyhK3u4+CF6EnEziA0xBr9uaVmRgZNR2GdKnioSKUBXeKN90vnlzKCEHvMSE8u8CoxkiId+QcsG
tuNz1yeQJXxG4F5F5nvN+sHXTgvMJyzes99oQkZ1AJYRB9MOcwJ1tKg5eCBihtWKhZJyVS0dso3j
yFM9JSlAO11db9l2JrseYRqZtFLXEb0rnr5csXhWLFjyyn3V1R7NXXGQBtB+szPED0e/+2H8An24
8vtOCEKbDCUFEGZL5uHdJI6+XhWhGTHc+yVZIK+TEnF0aKFb7mrws99LVj9tf5tC+Lvbwdg2rB0U
o6AkIxY3EIjl+CpP+Ni4hu9L/QJ8FuBrt95xe35kAARHIGs8mmHDn+n4YxjhL+lbRC2c+QxRmUNI
l+lWmEKqo4IPa0+YW/lB9RB7iKJFGST59xVa2wip2/S9cd6jTZ+FyV7kJObU97OjnfuBC2qrRt63
jOJPuak6JTq/G6wxCezUysqq/JU5sACJ+aHJJppAWv6ixa5Mop3CvZsiAa4pJ+M0FcAnV5f++KeM
PZ6SSHhZff+lOQS4sxsxNHG6lkH9dGS+OEgpXIOZ871e5/x07rcyH75QhTr/phI6k1e6aGrs5zIs
NG3xXyyczEj5mCcP2unk8Sdf26wgSSi/goF799Xe+d+kH0I2PGN+++iqh3tCO6Du1888ZZVohkuJ
iytnSq4xjk1DcXWSlO401r9VnzsmvMuoLmQqhXZHjad90m70ifvefG391gXqqGH7glBDLbslqMHA
OiHgd/XEz2Mwyy94Mf72fqoPKQiha3odcdUW2owrfriMhgoNKJ1D/Cfiybi8kKlGngs4SbSJEgBe
0GpRYN3JoUrZvf9GPW2iojcIqdd6B8fqEDoqVlFmoqWnC8ks+e1UVJ9Q8kKCkv62gfdDqW2WHbws
1ZQRvKgCbwKfsOKAIJGnd/0JfHCZWlcVIXvwAKOyUOMlnYsQI744Hpcs/Bn/vznEfnXw9iwsbwVN
mZyqw2/m41WzN1GUk4cRhMO7esgKdl5Y+rbuQl0sZ9bUGuDzqdbizVq3ussTI2KzwHJYjRJY00iq
9ivHpGm5CvuOEsAP3HXdCQewPrjO6Uqcy6YvsmLVgYxP0Ih/vrTkvZrzCgelxNZqvhnewES9IjBz
xL37J5qFH6kR27U/SZO8M4f9XQ45Xd9OlwN7cDUkQAiZdhF0PgyQEudCoKS4khIS3sRUi9w4nfHh
Y/t0sqYHhTDUuSct6ZzJXsjlqIdWPS+AFQld6R96YkDyl2eyo635FGwbORJmcUMjPmyp4Iai8DI/
JEWfWLwYJuLjg4bo0YuD5liGlBp5KadF+AK/1+uwCN92NV1/FPsef4kQxhJ65ZyBAeykuWyCV3QZ
1Ao0PkLG89SopUbr8xBlYMyB1xO++1oKjlU9Vq5oRXAwTfLBu9/dSbkND+YgT2Z3UY3CzDKe51J+
eJRs0tRq/34WMhvLkNdj80juCffIHhQs7vSKeZZshC54PFSS9qdJ6PBkIi2EFfdD8QDvb5ijbMbv
hIjNlYdpZEGYSBb9Ty7mBu03t8AvOFeaDD2hIqDohtpmrNZO8GSELRHIWhJDgONeGodLMfx1f2mH
3XzyyrX77h0gdgPhcNzAykjuln8q96pHU6CqAHGgD1oklwoNTIbjj7qzUjH2feFUDXhm3FAG434T
w6gJ4Sy7RlQVofjy2wcqXoZU5qwTW0bZ4tgZ7PTsuDwZKdu/Avse4hh6QTCT/6ToAITP2ys0FTIT
8XwymEMVyptaXQ2WnqFREg+YpE0CJqQKI5laEqZE8mizWrfbodZAU6qBwqxs1nxG7EE5e5xCa8hJ
xbKLxevbexgNPMQbqoYN9mStS8pxiKrhvS0MeN9D++eeqkZp3QYlnyMmn0H7jstXR8Gybidw4G96
IoEmRgFv24j7OqmqQ0pJwpjOvBIjtPNXjGk//YparDke5Xzn+nrauo6eDLV4EooapS9OcwO46glk
npjWE/M8UuUMyY+0nSMkPW2DKC0D4xMvAn3/CtEjnIBxzgrWLz17rSE/6QbEN0uqsNSMGE+Nv1rN
epnl3DQ12pB6MhaW7CO8ZsmUU54v2qWvTfDK3opN2ywMdDZmFlJ/An9rkq6VDmkzFO3IBfLM8w2U
hqaA9QvWW644zi5UEgGjGSKoUrOIKzEuIaZSSCBrl8D3Bnv3p8YF6vzGFQ5hEijEW7JQOsu9p9ZR
NrRh9L0gytJbb0BGYWjLIJLUadPsnz1HGYwKCZmFEm29FQhmFfYXOH4uzpf7X3UAmsBqOUeEzOEY
SCp+B2sT6tSKbwD+kDqPeCJpBEstSpYbqCEhMNLbZFSJ4kKJ02C/BFub93dSKJy8Bb6o1euhEzw/
vf4oDwH4VJNyaGEpTdwTXGVTtLtNjoY1CZzEv98qBGt9uubjO62KJJJbJWO5se4bDLWdan38LcfR
q7kCmDPY9SGEhKy1fkTa3NMKlREE0KmJWzBG3vmXIew2EygHI6JQYm++97thwBWT3lB+/Rce3l0Z
bvnHohjzdiuufOSUqQZBOFbHeK7k2UE2TG6F3hxRN8KVnzZ0DFoI2iAusmFwpB0UIensVBN26E+A
Opkg83Xt5P3d+t25ujcvkKRJIuXFYnhKVwGcyv6ZkXPaWV87VKAn70qSr5ighGe8JFdav0Ssc3Dd
sZRIy0pVndgVIG4klyZdwq+uZzb7jIXmN4sCD/WSUUWGuF+CiSROUA6m/ixHWRwoXIB/czRIARpO
ENYvgIDYiAukwOrzFLinjpVE2a8Cvac0Lsn90o/t6Prna/rndbiUjwb46LEWGlMP8doFEUsIq+mg
+duzYOK9vK8UjNOwaGLF4YxKhhq/tYe0banfhMYzR+6YJY8sTK+BtVWlEppDCGqMGEB7SEcYeoFM
Q+duZFaMoPD/4qX3OWu4L6qZhSP4mHJOuHtWACVVna/WqExun43WvCH8n2llXaStyr9q5sRG1n9p
OHYftDowxF+02BL6pe8UOPaWTctPGIaMlc9v6+YODrnITtjxV8H8AvTgGfFXtQiunienKL1dQCKw
4faQkMNgfYU/5imw//QyRMQsw8dFFL39YBEyrvIGcFmWnZZWlY8YP7Pe5g99g5kV0+EAO1gR4t4F
dqWqthkUPJtHISSv/9BiSial0LEnUTyEWboRfjGdHBE2Ai8gIfvdm/EQxomtGTw6CP+f9bS7/Gbv
NLgB5u88Ll29EDnI6SKnYMVfVh+JpVdqGNDetaqFd5YYLClI+fCdpXvFAdO6cPlwH/WiqFNAfJWb
/ESFy/zZcBuq6B+0Yycq4L/m6F+Rg/fyfP5x/SRhcFH3uoTAs1hZwcGEqD0I8wUUnJhALTDWrTum
d6zHSbd4zK7sD/PE2oyPUZQGDcARqrxHayYv8+OVpxVW7vtBHBhjFRIODbqAYsHbhrPsmRiNXvz9
iWa5u7/pyEbvNVrmcSSUZW0EitJ6xcPYLv3UAGZ0UDeUc4O1ggI7oyYhW1U1y9ug2GJ5IYFaI+oH
lZXf/9OfUDmlt64NiNi9SzRGUDnzaLo0YkNHh4Eyp5yBb6JMV36BA7JAEIs+ax8jw+31FgZ7g3MP
PQCNyP4mFZnZ27opwQvwtJ5I4hJnMMkJyg9F1gST2+ovn2IjlKKUQt6LUj3052MH6qTq+qo8o7r5
cAz/tjKp4TfSffMvS42X0cgs6K+Zx5yBb71p4hMXDzMnMUMKhhAC4g6QqDmDfUv1mn+Km2Xsezfy
Dznr7RRZ1uQOSvMH0aIfQwLlu4zL6pue94+l/5pbOr65NyHG8mGhcWR5PAl1MfNiaa+L2wSEF+PU
XGblAHMO2NG8ESwM0dgraOjh6zYiSVK+u8BFlJb27ZIIrkx+DNHPFqwtPYRHiAGguxAsyMj6bTuz
v4J/ZbZoUKvDLcZHjBS6g8dlcyXtjUlirps93qRQDtw5jq1tL5prHt4/CobLMxkGXN8P0QDG8gHx
ti2gb/6UnFK8nO6CxQFv+3xSobgSYn65RWSfAPlsFhq/3e7ClfT+S0DjkwLKujbY4xTVfbqSQuvu
S2BvgN57+/09y+EpYPWZ14B7x72FQe/5To707RR+M4Yisb53A71CvV+EGMSlU2K4wda3JWUAjY4d
ypm1VIYq4q/kFWjWi3QaTKTlEJDwFyqx/K1SZBvbzqspw3/JXNTids7AMsD4pZ69ULayR+geDSB/
LZUZoxEJMVQZxJb6RbkDXDSDeM+qqkup8PgDrLRD7pKXlmqC4wlQEK0L0YxeRyLkIZli0f9EBNPL
i96G4GB2p644M+mPRz1/WNCZR68I/oRjkle+6qKoqYZf7PtwuEoSjtPhIR0skuhwZfw779B+hLZ8
9D6NUHHoxGeablomvyKciR1/4jSSK7m0FuPazLLvW7vWyxVAYOZu1r6DYBIUfYogaV2xpxT1LooS
yhESC/m2EB+jrxRXwP6u81Wk6f9RkAnUNk+Gal6+e85qgT4yx86apQST8BjtxYXKrD6yjV1FnLG1
OI4cHSRnitm58UyhpAb4BgDOuaTnlc0MwNrAdTI5Xbp/ZtUXVKWFjLiQKIWVA5WUfNBWpiYko8V3
RpFmGUClxEMvDtkV2YYG0jntxKnigpTirrkQ2Xcgt4yr1/VSQdqlePqZ8YmpmwaNPbRQIy0SjM+l
TXx5FNxhkhg09jRr4/v0RFK8LnZy9QjSf38yBQZSJEkf80CluMEyNWDklxIQepgK+kEbp9XkMNfO
+taMgQOsLuEkYqiq54CvGQgThociPwBzRAUvBbxpPGF4eBJJ4gt4PE2db7oNgK+22lpRQMr66Sv0
egVrYXRoucPvDveoeZUH3fWeeIdnq7/Kba8iHKpaLgSRQeRagN5IfczvgtXnrIBk4bn2/wZvug5y
TtnvNNC21fJWraG9JIsdU7/IjjWhTlbbeQ+5+C72IBW/m8DMXOdcklixaYtIr5wW5FEICf6W/WEF
qd4ac/VUBPiMGeMhy9X/eM5lK6WybIM9txZ0V/4jj5TslFEDmqn5BgvpRW7RmKXAwnyv3eA0/VKD
eLK1dGgRwK8asdTE/URZr5YpJJL+ALMyBRAV3wxmrvCrW45r8p3+D1ZQfJjuil+6KUokhzEJhOl+
JJpchWHMp0xIU6LlOQ9HYVWIJP12l1Xv+rP3Gy1OMmDmuCAn+tx+hPBjDUXHb6NBBgNMdJhlLmud
7MF+OILizT+gVM4ZGhENxxsnCaqwvzACG56DGKEDaTRR/VS8WJWF1gAoDZEF63Sg5O5CemJUzpEO
I8i1vgfuakd+ZmDtiKnW8CVGY76q8TZdJEf8m9mlMsxRLMbXcNm1lkwLnUznmK+QAVs4o02wydzf
qmpNui4qm1/KwnhU6f4pUhhnebevIjsvHnPAnP1Pyi1+4/lMQOi9OyzPFUvLiwGrMCXsoia824Xp
Nw1v1Mvmk2SXyybLiQ1kPdiEEQEpJnyc76q2CnAyoxncUXQEQ5lCa5bjOBhJn5OeioT5nkUGo1CC
NZs+k7yG3FW4qvYnqJFJJTGPOKja8NUqoy29q7rbhqG43IMNaHv9HWOtv8Yn1Xbt6otTH+mwVYEV
cKZQMmYQRMN5FkH4rJPE3hOdYRYHTemvYAEgQRgHoQksVpXqa/6QwnO001pPAWS+t45YQW0M4eMa
o91B12Yd0BeOS/jnDqy1Py3SUbb8W6V0kyBrvwNpI4O9FPFrnqxVgUGBnkXNgUjcJU33ZTnn6aqq
dy6L6ZvYyTn1G4H6QQ5yYe1041Kwuzhmmq6dk0FDmKdi8sn2KjQQ3tzJTbgQwqdGLgpAwNfQi24f
ARnsnmqX8M4Y82M1uZiibqvooWTfQGQDhhMQRNZPnHyASmBgxjYp9ANxgn/PKUWO+hyjSCXftJvX
ohXIhlKzOiZFLqthE+kh/yi0/cAkdxtLHGGGykkstrBWBh102JOsRO7fMiWInvFc2tUO4LmlOQrJ
nkFAcP5p1ObLnGGAWhs4i2DvdmqIjEvx1eNd1zfEOl9Hg6LVpk8JJeSKbhDksbQmUS+GcOIykv05
g9ujxjCTj/QCT1SFNvoyySBIm4ltXklOrdI7ZKGoco9oHpZt+zV+tZJxjDNgGZsm6f1QaNwKvgjO
fH7JVlxHcsrR/DaDNnjAcG1gpytEfXB8YEoQoAEQRW7JDc6Y6TJda3v1VxTZ27EwX4vYUHTPwcLi
FRX8tJc01Oue+D4jYxMBFLaeGndQCRr01ZX4jCOlu6MucAjArYSXqSWK+rpHo4ZngprhWYJsrpmo
AcvQ1TqIXn8u4f3cnTl89VRP/mR6I0dDKGQhCJLa/HcK5BrzeDjtgi2Mx440DtoxfgUvdpOwvaOr
9ANUc6sU58dFMCY2zdQiEE0sdv0ASQBPhqV+HCBmUZLorstFoL9LO4vVHpKjrFKoOVKhSyzlt0C0
I31ofl6fBTDjnzW4iSpKxv5YHlHA2UEoChvwGMRShz1quOpUKzkjLfsAUwon3I4kKnFFTWLtjxGA
CcZUNCLvtiB5bjGP3lnMUyv8zd37qaJS1QbDPnW4dJL7etBnlZrkVbplFK8mxxLxs6bOjpNpUQee
weEp8okcWrBz45sryFDGmBIjVWarGcLgDdgGfbd2Xi1+8coirtfQAYc3D39aJeu1Tc0VvhjIHGk1
1W476d1UvZAI/nzJew7wMwuoVmxT153myglKVsCMblhNZvHjdVibCGCuvb/AOTS4Q70lxCo/Sflu
pCf4+eEsKMHo/9WYvfyHU8rEBhP75ZqvJvfjrFO6eRLhDHG0MkOV+sTyjrZaetVfyKjQt6lnqQH0
wsAM/62ccud0C1K9C6q/k0fuvQfIUBmBi/VLJzdWztfjP7V8dHnAQzuNgVtUSoFJvwYkodkt0AOr
tRrORygk1UYN5YnphEkZLT2X11tLVxHcixiHz7CHtid1yrHDVC2gkHokDU9YrO6WwkACS6xzT4EK
/K3ffK3ZWtKZIUbOPF4Nw05UNl98qphgO2yxB93cWaUAiFQnrQ6FgwzRE9oJASmEkH5ScfbLjG24
2nM52y3Tc0jF3qgJgR2l9rVhry/SJ0BTsymQhl0XzpfgRENxEcDZZcAuSa3keCb9RIEMPNULGdgF
GAeMq/ls58WuKEU6sy+BCxopileGpmSp7YJnrFoka9PLQuZ9svusEh5RhLcEn5EFiYfRG4UsGJ0z
UX8F8dwJIpATPfZlXk4kuM2sHWTsKcV65vEDexUu56PTR0Rzltf0hwjidYB4QKpbPiTzEXXhO8R8
lNiIr3pzCPW2+u9W6KvfrdQSH6fileLXOF+6IaqDyZRIAvSzz/8bbUgJJvcQA85FbN/2uZtJKlfM
xLHH7op5OhmIZeRUGy83SFKhwFYkSQkqwhRcij0CfRdgLowhtUa243M73ifNGHcsTU1KMYWtZG35
cRgO5+roBfq+cz4zw7v+9HWgGvqX5PGcE/mirQUsu17jdlcr7+VXL7a9CIt1Jm2fnoKGV2Vczkky
AypYAgoZO1FA9cajJ4/6mT0vWrC4OgnNvHWjjRJwAV8r6WFLh8xpt2kRF7RQv4xyOPnlCKCHrJHf
lKeCZw4qzeK5PETcrvQMJcDlhKF1SiDkhIfVMHEjWXmxV0G5HeuBzZ5l9Ff2j7GzTTroaSpytcEx
yXO5Z6LvaOSS2l35dOgIObTzf1Q3lUxbYNCUgY52DYn3V900NFCYjsDlnApXIVl4ZDwwyD5OE4la
JWldwF/1lfKKsw12E/7xmysvBVZN3T3xl7wOBxNLWpjl4hfIV3Tr9lNjepbLEnUMJh1BBKIdloU5
8/DfSly126NszB+qtdo9lEYi4rVbpeM5WLfu5SugAs6cVkBMwnwbd851GqlYGPIlN+IDWMGsBHtB
o6Gmqfic38f0LppWWL1xtxMiASWCsXEervN2iV3N5dEyou31RG6GbUMR+sHkdFfIHF/vb/lrHVzc
eLP9tMxifxqDaMFzSdN8tKrP9EPj25zJ+c91LWvuYuxiNQ/olO922mlLevBpWCwcJS+Vk2uSrPGC
jACWW2whh8v6iqJR1vxBDNzccIo+ukfDxhpJ+F9Nmf+DykXsAFsZzXg94QQ1yhWs8qS+yLpHW3kA
wBufL1Las4NyjETAxjeGfOO5CPhUIUVEu0b2TgoVDPhwfNVSvl96qa8dPm6fSbUBG1uYAlNUYngB
3/6YgvV59AiY2+A5c21w2hcvMFbHbTDIqDxrcqMh4+WkilzB7HLMoA1vmrOK0xO684Ln63pxcojp
RhoQS4SgURNpW/s7CX6D7455RVwxZzLb3C0v2yWDQ3RADKmxJRcug4we1kSnzwLKbFqEdMo8T9pl
qcvNBWM5Vv9xxvj47n+jCjzX4w/H4WLaXfdf4mWQCpmDvq723zGniF+Ew3AEXDxeKTaV0xzkTe4Z
kgYA4GYy9EfrRtXr/X4nVhcS0HRLAl06EPRdjFK9n/xbHWGKjmWiuZ3fFPOKOPuOzUBjBkzbJIsJ
E2fmJKZYcsJbgtmAdfylhofawL5DCF3WVXCczaWgmqUusS6bhiguz9rqObGaOydzA9L8pM2zDVJj
w4QdOjGnfYWChEuI/xtT/4vcjGWn5jDDcjgd+e90pQFXostin1/9rfzVjrZUgZLHfkbwtd3+ChjF
i0bS+gTeD+wqWRJDBu2XeWwwjR6evNoWgxPRlNdf3YKPRx+k+PVIJ/lqzMZaK97T8R4rzRUUnLh+
JtHGwgpwgKTmj5pl4Er8fFijtpqaT3u6Gjsf6My7fK3Vm0zbPKN9Xdwadt85xCTkFVj/7DoA2oQo
5nA4FiD1xj0/QYHVNd6bf/CpiEy5s3PP9vMzx2k5yZojAOI/iBOxyntLGD8QXa2/w2j9fnSVk92K
ZMe9btp5cMhW+s+0worAx1zSPhjmM5zLP+NCXK9v8pDcsa6TBVuBpnYM+uCL0N5ofoWGjLEEbG0/
2Z36q2D4V2+MO3O7Y3/WCyhlG5pBPu59YNP7qFHphUTUKQht1bJQUs+aXqDtkBHBW55L1vMwQxi6
nMMRPGFZgB9GRLK6qpvCLbPUr2yWidH5oEKXAtlSzm8TD0AetV8FH+rsDls4Q2VMPp8v8262FTvu
VgRpRXejRiKCKUlabLoAOWIDsKjLef37TeNrv/LOdMd1wR2U7PPro7vhDVhNvrR0STVZCiNAdPQ0
XBQ4fj4vYK1inEfFNEeLLh5pBeVqe6wTG1b5xu52GptmIPwGAx5FLypJU5TT5q3cN0wPi2fFLSOK
slajpBdE4DxqDhbccc8wVRIBn8ZCcfoUjpsf3RK2/ecXX+1TqvZ1tugz8nzPMXge1mMeEcJT9WPz
weim2WiWkk1jO795quOC3rtBwxw9yNN2+gacgUuR+u78ZM5bR1rrLyrOtZPjDAT1MQ9LlxFAONnW
nv13kvXcXBLUwLI56/wCnfzNv4qRDC2l3qkagrwcoa15s2lpAN/SephWMJSN+omJDoKx7zCHKRnn
Ckumxftqb509+uHNKBiIBslbZTu7dD5/PpZWzHekrnEmoNeEHgNIjCDMVOExZQk882QzT14ZNs2Z
xFUMuxzAAfHy89LGWdga9wp3DFNg+C3TNL4pmpQJaVAyMbcRTvLmMp3D06SZyJQZ22KtyvhZ4mSn
BN/wV7H/ybAQuC8keLev4EmpWpeN5e78JEOKM/qjWamdzTRIDw1FJgm566sxr3hYejezyrA9NHRi
BrElyooiAZA5Y1i96V2vdoTqQHAb9SoB6nlufENThuWpncYOr2N8E8bmdIUNea13cwY/VmKyy469
pZYWCs5cLoJWnoeun+PB0ia59PpfAfjoWe5UUVjknvveAaIUjhB09s7TkdpILUWZ70wG9YBzg6ts
f8SxlYDCqUcZz+xVSgDNtQRa/1D3JwlZD8hjVwPmKF9fiKPYoT9P0DLaLM3Rn8Yf0D0HGZK6BzTN
BB7J7cO++KKyAO5I/vRKB6QxMgOlXD39pOcAj1nJt6dzV3OrOP1/+2VlKlnmahAXqA6s/B3+Vqps
WbnuxtQ85tVDKr8j8glm4VFsCXgojpWQ0ViVMmOpIKYICOq+wtw8ei8ksciVDmHynKIr+Abcl6uY
5RATl1eczaHqPXUh8+DIh37D5Ugbn+rqtWlRtYq7efD4PSOflJC/c0cNlbAR+k82/1aDxKPXMAkM
WID2ag/yeQVSM4XqDZbIsVAk5YVFzzYyVej45al7Z58dejX91Sdd1UD6954i7RRAvFbNiPE8NLhZ
2mg1g9RA7T83v00NjBhaUUGbvBtfn3NxmGPSAxTmTjl50q7n+cnPpUpGLupOG92oDbbTBILzQSHL
0xcDBn/zcxmF3w7KQPrsesPeD7jJovBPFrXSc3BrnZ8Axcb94VsClpOFoLhYnRE3IhBMHPRungxB
jv2mB6o7kpxap2mlV0kQIphExe55LjXDkYJLOe5+9UY6u6Jf68WOBXIZD3vMZQIdWVrXslWIIhvp
xZO9eGWbm0iy3HzNm6WwvRxs/foU/BPqaE4KgG6PM9MFGUZSO4ih1a1jYIt8rTR1iHqu+/n88AlZ
v2Psp3BqjwvFGooRNipYp2XT5HmSdfO0YvZv1MQi+hM2pNIgoEhqS2HeTaDNzqtE6l+3dy3vNXW6
pOQkPRBFcgob6WX0HmLxLEPQ/fN6wsSEmK/+3/ZpI58PeBKO+sWK8ZFXBI5+o3NYOwCekSAwjezJ
Cj3cfFkYUzPBnRksIGFaW6OcMT9jQELnQzI+0xyAf6OS8c8pu1MVDXEHlvQecv9jA9FJf1117x5g
vR07Pm8Oye6ISRp7fWTC25PKwHDVjIk8p/VDIPxmIn+luSYtCIeVZDrPG/svaCN9djM4JsaSscgk
UY7BQnRZhPPeZXgxjlDnpkKkw/clRdQ0ESoHMxL31CU35+thNkjn42aUjTrntlY8Z31k5gu/0FT7
GUEDy06YzhNMiVUWXDW0yL0ew5V326p1QxVmWvb90U6DdyN/qDB+aR0hRRWbRg8NzOjzTpo52HSY
PacoNR7fmfCmU3PFooUhrQ6Nlwiu/pheAKeksB0mPobqDGrrZRuzPsrq3JNVnZGAH4EyFha1OhHY
46QSkMUwh3Fnz10pwUAvXMD8ABPBSCnwWoWQiROIzDaVW9Q3uHUSY5sulbuD4PPHBtTQue6VWHuF
Mms5/ocxWdgZgwic+P3rqvRiFSCSBZlBnyNqHMdTI++k9F7Wuq/XziVnJTfuYNvQoIbL6Q95jpNe
OJajezNJrwgPe4jiqcOaXyufDPncGn1vNV2ryzQ6orzW1DTj335dGR4QNE2BNo7vWdY6WQvXEQoX
saA75iNZBROrw9RwtP9SR+R24ayjQct5s0NSVPdHGQvAnrwI7kvX1QN7gyDn9a5SgjWJNZDH5GuT
xf4LZwx8Cw2gclN0nQeS/xvyou0ajB0snH9CH6KHUpRhE3hlMsCEEzrWfZwTD3O10uNOYPozR7vR
/X5F05+JiPRADjVC35CZ+b/Mz0fkRVfgdWKyWbxrLCW/x+kxJX4GrsV5ZQ7yxHTNwlDuFwyDBcoX
u0SP34T9D5LwL2KqDbq767SNvf2UrHoVhbHzuP2ItdFa4c1LNJfpk0b3nsZXJDhEzIKn+0nLgFiz
VLuMcVvy0YYTvMgHv77W56y8cYdrCpAq3BPEPyeDIZJuVjEK3uMfU5U6PqYKmnud+m2VqA0WIjNb
mt2ZBCumM1RvrKqkoXlpMfGxz0uHSVVNjDChRNcYUsd5zKaGrCAMRszvK3mJ9VljlbGKuDoFGtG6
bNCZtmbaojuwZr9j1RR+1n3cSXngkwS9OhBgMSbInSo8aD5Sg192lz2AgzxDREcEAWDn4IrMFRrv
1d+qDI/A6Lo2GoYFkTg/4Ux65IaYIlSMImvatnUPpvlH+/JcvAx0ax8CNeS709OV8arlBrElJOSg
yuCeLpAafhCzad2ZBiqKMNWNknp+XkfXrq9LYxFoTp6mrqADuiPzv5fSOWxilYAi7OdbPAg9wmcG
Qs9sK5zZE4jFxEpYzVPFsZo7kjVgdkp4sDTdwFJ8G2e6d0fhOqop+n6qSeL19wbZNf/cNbRHYfQL
S9Lx0qtwyynD0fY3h7SPLL3mnppW1+gUGBSHtJPlnw4LspbFdu1kVSrZF7AsjZVFizP+UVWiY8fl
8QbyxGp+ymD1fUkJCmDsmpcQUEKH42jdUzIeuABYRt+R+Zp+/mVz1sHnVQRORCvbikBQu6Dw2vxk
0CNaDZv1CzerTvY2w3MQLImFNfkniNEEjc4TW2KS1nEzmEVxkRDlTfS6Se2djG1k2Dtyg1Ba68z5
0JaKWejqHJojvsKd8ZvNEs/DvIng768pp18tR8f95AUEkKcpHv/fnq2xu7Z6jIIiXdbsIE8l6hpq
BbqAH8gGzSDmo/muW6vh0LAsPjSgoA/WoktlcvTUuIB4/aDSd8hzhJcdgmV9gd9l6R4LacN5fx86
CBvBtb6vP0CZsZIEHOiXqxwsd0r+wJAN4teMqpxlDZ+1nFPUlXaeeQy9MvxL7s0u6ko+dKWf46R+
RR+q0VFwoyUnGcyu2yec8k0TDmqwuH71OBufQmQL+E0ukKxNSV22IIIv92fyH3IxOS31Ppwwvxn7
/ywE4n+6ScYF/Ndi52VNa8ZM0/DOwX7NBH2czEKZYs8oeD/aeDwkm7zdNi8I5ERKcRBjl1eS5vNc
NSIhi+v0Yf0Bht6KNK8fcqt//JnRj/aszlLU/COMA/H9K14LR+HtsPaPpEPC0CUYwJV9jvY90X2d
4r2gEvOiGhEFFcDSyrBGJ0V59R+a8yc/tu8CXjays23JRjPy7ypRzWu0kAIjKAWeK3km+MtcqU2u
9F33NUTeOtKGEkxVPJsjZPCgsWFUbuPLDi5VrWt/4yiWl/plYNRVoF16RY/98B0rnZIOK2A6u1kq
tbXQagPv0JOe0kmTdxqO8FthSTjPPuo5dNiGQQTECR7V4yQs8oIIsDdZ+m0hvZadJFzYY2iRHfbc
Rl/+AzT58fOQgUAJ0Jnheh0UFui9xuASZ6yhLiwpOlcGJrSQMoqdB3+hS+RMcPfPGGrUaMIiukdi
5z+cCIDXSFZJepopuP+h1XmB+ld8KKDhWSatqraGKE7V8NX/CV+JYWFzq9+WO3eM1AzSao02wUbl
/VWuIkIYOXO2TmLQvQ31iQN8j2HHQl3bcbzB61g2oPzw6AwjT+H+m00uMC3VRPGtlJ6gAzp4hyNc
EwNeD9dsl7EVRm46iox5CnJoYA/jNzlAqZ1XS6G7ZqPx0/rlrU4KnkFuJOSCUge1lSK1cY8EuU4V
Q8Z0vRuUMU51KYOhdyNK1pnQK1jnxenD1gxqrK09BXxWOiSLFHJ28adpfOvXqT0c+9RcxCAiEQ+4
aQLFoGmvFkMvtKuQN4hds3no5JeMIvQzLZRAgMsqtSxQPmfM9N4osMYIcCg1V/xE/RvPt+YKWEqj
CEXnPmZFgs7jr2gzIB8VJpa2W6Htt3OhbNT+hffgpzmyUJhe55tck0rRGHSuFzuqeh5swMUwdGmz
7iegDEZhFMvq04zzn9WLVU2hBJgJPAbPqWhEDP9Wzc6IvQtmbqiGeVUdmEWKPNZZChl3uy+QUIB2
ps1QyEo+ln9m+R90Ce2JicFJZY5o+FPnA7e9bDPdX8y6WBgLFc9VDKOrT3MCJfhNXX43VOh4rovx
KKQq3Cn8pbda/NQPDNr+680EOKeYM4V2i9d5fHl0Hg2BgHQhQqHMY5ng6Pmvt7xGDblG+KnKHxK2
4bOpjE0iZtBM2xI0GOBMNCYmOqXOwPkslmzijB9FvfMHeaq8pIYljUHHYz2SmntHvjKlojQRz+h1
1XDAu2lU1UHy5pta9cMvuGsHG65CtNC8fu9YmWZJ297V/JbRoNwZDCYEYwsXwvdoZQiJIsmxFEQ8
73ftGvIpqT7KtqMS5lunDs0RuZbPmSbmGhfbAAAD4qdzbAQV6AW12HoQoP/F31a+5KTu6rUj0Yn6
n2K854YBYsan8EFDVE9OY2nup6X6O5feoY0lijxRUcy520cAue1DnXExjTNRBEyF9BkvRW/qv3h+
AuhTsgylM+qJ8YR0CHhRorzs1T8YrThWvGPvQ7JbJPPtXgPiUT/XGvT3cQMwjNIHpYQCf8na9I4i
zZB+aJs9wbSQZDItTsOYn0l35c6/wZCOQmyMGukiUn7Y+d/ierU/wbCwby2G0Mp4LneI1GuHPRzC
/qwvyGJrCjO7s+1Yj3oV3R95Zk+YQZA4Nkc+NAAMQ7ufNMyUKN8K6X3mc+VPa8hon0Zm7g8r5Z+Z
vCrIDCRt7mi3w3TtO9PHg2FuyrmDjykvCSykbZL4dwDhqc4xg0QBi9WT8VLTK3oV81/ALBfZVibc
qr07A2MOXgKkjXHIk6YMN5TDBbbgVIKHzysplpHWLMKVAcozUIFzUW46iDgYc0y7/8EEh/xcCoUr
A+maRdxiF6S0P9/oYpycM+Rv1lk1Oq4Jp4obJSUhLI9yKcJiWCtFVO7oWTts0+IuV7hxgIfTpIeu
h+h3adX8z7mEvKO/e+jO4fWrLVEkagYhErEuw9OACWSCcp3Gu2xK4kPGq2motXDZHgQDvcZ4406Z
ZTmfEraN2/xsvpXqdLHFx3YgrV735DOlcTAtwG4wf14emEPF15xPqr+7DeZf4Gyuq/lTYfLvAC7L
DFqp8PoUxl1ZDy0IzoUw8HJi8hUIVCL4NSD6OxCu7kfD7TV0UtllvCZUeyC8yKLUA629fA1YJ7J9
gtITXpAYuamY8r4ayVFV4d45PCX+Bkqk7piDqpQaMTGQycEIbwbmo3b6kNsjPxxMBuL0VuKdV2Gx
bYEjxLtUDADEALD+tVFavkO+f2oMwPPVVNZEFHRcGlY/R7nXdVm54cKlYU7TK2MBMyjFJWy3smfC
XbamSPQAIFzXyjiOx+m3NzxvfuooND5q8fKFLca1HpKMQOdMbSXGxlkmuwGoimsK3EF9SUHCSlXh
W7ujIMSVA8yXkAgE2aAD8FKiT9xJi0KzQlMUv9ZxdbQJl8DqhPfkqhlgeKPSeG1Y5ZD8B4gVw7rT
oeQfE3mLT+lt4OASs7nWzu5bZxVhptJbYJF+5Q2ZYYSrfHwVzKFCcNUIrDZscL2KmeyqpSNo6XaC
W4SQSgBRbpmOU+nVT4KNpA4OzCn5+715E3yEJ9Ul9803BTBbDZNvvK+8p+rsxXb2qzdmvi9QMpYd
q29dJ8gpgFlbfNBuq1Zefe6HG0fAWGN3kpIw193PW3bQ5AuFNHXT11HBrLLTzJ5UFgJK91dcwuJ2
ml+3jfnostEHVbOcyBAR6JjjTIIpO7cFQLY8H384xkkii6M0uZ+yHWB8zrbhoIyJQ6aqOOG41Mlg
V13y+jLrcXPGn4VfiM932B3H432JQ01F/hNVxZPUdXWtcfBht4qlBRZhdz7doT3ZQ0ms6S2lwoa+
+6q65XjIwd1GyVxBOVUbdRFORYo9oSbfx6xIwXQjQlWWVkzdEyq/aILKHG77VlfLF+IpaGDD51cO
KuQGSzhbKrK01hnTHstQCk6reh89Em1qXAKYF2HNp/ICQtd7p0aygv0O3+cytpj509Kug+fBMi74
N5krsbdKAy58Mj8gtCFLqgUmJPfZJsPW1A4YWEI+I7GcRqecGrvIkofTn7P1zx5508xobbQop2RG
GzG1LzdS4ccixPIfJCjwQXEcG2TCdhEqAvmtXKmxl6jMMLkUYr2Hc+hhfyAyP76qKmUtZ+C9JZNp
t85MOEddA0oqpyNRKRFoTjzCcv7p9VhrHsBb+wx5mT7l08XB8d3oKW8CA0J4TqL0ZBYxiyq5uIJm
Fs7Dlt4vFzoYdiLQvDkbyrgQ0taa8iO4s/m5eU9KbCed6Jy5Q4l/qKDaFdFNLnuBqnWlzyZuXe2J
kVr0DFPPCwoYi+XgmzTBKstx50PZmCv7/Is/Rh/BvznK6IMljWp8/XisXhZiwvXpRFh3AzuZG5to
8Cd9VMaR4OYS5rRhtGLAR9XSSOwgsXnPWjYKoRup9wQpMgB4dT2txgLfGalL9cw/IFFy3hVCle1t
V8WfWnNFW32fU9D2su4AmnF/u2ktYppsoSqQ46/OJg7xjsadUwf2ZNK8zKeXkYDnCVUAmgtsvPdA
BOsEXPeYEbjf7rsXX8vqAoXwuVUU4M9sLypCPbyBBa4tn8ugBaJ0idXc6r2rKYf73L0GC6bM5FuE
+il7b6H+0GHzNiIYWyzw1aVU45iSH3wAiuePXb9g+NH/EYsD4mK9xpuVEA+ydwRC4v3kGShj6s6O
ChvJagjSidixG7o09rtQUQQixhnoLxoMtqs9NAxV6CXcv1o9MBO1/36nVnXW5wXCV+x0VIeLUXrg
5I0/klZZJXePu/yqDFlRpHOYK3Fw48SMQPZakRyrttu43EBZQMTsg1NympvMIfWLR3ZmymUN6hrq
VAZJDH1rXtJjhJdJlj62uYXrtBlc4efwjzM12xBIGbsC6yQOUrEB19QrTjIyrLCatUVJwijobxlE
K9YqsUWdHpGq6hpuEKHK46Gfh5i2RSIQkrf+J7Rnu70sKC04Q1JZEz+9KJfHJhjMxdSwYtDooZVS
H2mSbmFW9pimyPO/XvnH9pUsinhIxO9wMUVEW5IkRVIxZlmeQ2mclkUG6aJsF8nyIRReo97B9HuW
b4zbBmhIVDPEMJFSJlJ7MracJFQ03F+hMoRPC5xPIfJjEUXfqvzAN4lUwtNLHHBuILEy8UkjkiRJ
6rG5b2o2oQ97A3R7MqBu1KV1DZh0ogBanindwYAFgpLweyQVxvNRhk53uVbQ4pi1H7J5RYq5uEYp
WyZH35Dp1nnAs7CvUWbF9NLQrgAHHKQu5gCHHK0YiPQHod7s1ok783jDflLa6y07EZtqgTICkoV6
EIHjRombH0zPDotQN92uqvceQYeS3o03w/2UruhxDQ/zUiSgLddLAznEt7GodpixcCAHnTdWQf62
M+og/ZtLYnb7N7NatEbEh/X2xYQbvRzj3YidcCCoKYCb7Niz9a9NZArvumYhm3ZBEdmbvSHJtyaA
rgNue1+LjzVvqVg5bf4whuXTVK5UzKxQS7jZ5YizXdDKjwMXTGICwI170eCJ7Kr8fiClZjW4GOI3
W6w9XJIiijCYhGnOQ3ALRWZM2MRPSR5PZnW/MV5p4IkAFHQ3E9ybs0Qjyn3ipZibj5bRY501TeXS
FxQ+2060CoC1NN1n/NXfYyhngG9pEqfGAA0uqEhPT0a3nvTR0Y3715MK3g4ld7vxknRBwMMDIIn0
Jd9Z4mjXf/WmPYm4+1qS2IIYDY23KicdP8QFZoBcG1ORDMVoiph4QWnU5koT1FBhRmF9a2u4LeYs
jXXm7ZxO9JxnLKE72bJKj0CyFiTx0CwOsY3KP+sFMwzAlT/fEa+Zu8PooJVl/uiYQm+IfiC/KH5B
EwrS0C4Hci0XQmKekHkPj/USFfm2cePVJaClyLHTl22fNPkAilacrVOlyjTOB3YvnaIFNm6b2ooJ
gHymB2yqdNi8b04/nn1O2+IsNHSJWh/FD2aJc52v1H97tOBe2EWqZURqADZvVosugwwGbzvgvZYQ
QB2987zF6erOt5ZKA01+fxSxysBjDJFO/qtwSgJ8+BN9JRmNmKCp9BAyI8ATuv0fw8ow/LOBpfJz
ALWAeYO8BjdEWgL0x4jH+33neR/LL7KotlYYJrv8j57pVripV7RAtCfvHx/0sjmWZIdKWdY8R8HN
GWGmgTpRWjcpwJu0M0Il1QUOqtxHOtBAZxtQEjU4eLnSkCGIRQpe1Y05KnanuGpuFJTjU8S4c2zU
UWDPf4bVBjc67o0t3c0V3Oa+uNweFDgB8XTXGqcwBsk8wZYhHfr/3zNGuF/wxLOE25U+GrsC9GYZ
Qh5yu5uOJQGOzyZndVV6f1e4UvwVPXNljx4ZAr3k9j/xhYYnS+TXEWv3rwDkBIthUlU1TZo6tQOD
G1FrnFF9bVT6P6TmnoRw3R+56RDTSq8vvyPqGxUJC3wU3M/hlBeAN/DvnjHz+Thfkpfk1cbuW8QL
++4S4AxKGShxoxVuUupb76/a/BtxhG2nKh0ZEEK8I3qwoI0kZOcmFViBZB0fbOXK5Ugg1BrOHmb7
+SRfnKfEalOct0MWBhruG/K2u0gBwbdiCRqd5tjUobVwNn4/QiwOCxki5R56bnzLiB1sx2jpoOtv
j0LgqAfDq5mKOmJNzJakN19eHa9SqX0jA5haltHlUqywtViKEXg7ennL9xpQdmxOEcXqhvRdpWZ4
3SR7gQjYyIY6dY0KeVXJ9zIGOR7UIRQ0RJvxQ5gkVz2kS0wOBJ4GM41Sng/cdUdGumukoTv9WSMO
aMtOkQbpMAC+LdHWhk7RoDy0WwkKnqibqBXrqEW7gcCfP1624AWwGyZkrBLFCFhA3SaubhOkFBYo
XyKpCRnUHvQi4MKCwFRt6rJQnSOzl22XzNM+nEZ7datXFOdhzFo7zcykcdRvszMrq/vXIdzm29UO
/RP0ijCgsbPyOA0MsBgd0tFh3OVYBU2g/eeA2/bfwoLYOnrFh9DuBO2o2tzkpJeZXQMGR1M5Drm2
aJWIRZ+dg2dlojUAJguk5IWcQ5Rw2iNiK2kpO04PeHwYyYYDmHkZKN2oVCARs+U2+3MgzAPkyrCg
7VWbMtXhvkKeoJlYfkAmGO8eS+2vuZ8KPuFq4APv8a+goz3NUvS3N9HXcN01s2pm6W5TBseunkOg
FtdPKBre1jEvT7ShJPzwWWTjfkFm+lZVKKnD9N3MbOHaB0CTi4kmq10CMpWdLSET4MiOuG+HTQs7
VzAQhbskKAxzrTli88TrVIIv0UmCC5nde9YCpGzY9KBC2qiWS0AhDEY2vRpr+QlxM5mUfGXBPa/D
EcWYwuATwb6vsrXjPapHfj8e6bGBmJ9++Pl8XqIcWIYmV05FoB8AANbpRu8G13+SnhYNl5TdXmiv
ONCCN/09SFWgZV/AKLQIvtfht0mLeMa9NNePbxyHcf0L/UUM/sbN7dfqjibRDDHLarMhAdnKwYyj
cvbTRlyyc8I4TdlsjjkdjhJi03qSv3S5mzCX/2Dj+5Wv6q0snCPoBst5fKbfB8t54fKibdF9C6fn
ZtYxlucEpIzHfdgmsfxjb7TRGVNfv1+Uj7l0sLR+U2qMz9q7DXiOCuhdP9AYHrUtrFLO6QfxTxDL
T0r3peEYHBGAAVbqcS4KR7SZsLk5FypTFsy+ZWbH7MMTJUOClK4mLBf0+EJINWnKpW0E7Qg0N4xx
agYiVvtroZJWmcnYp8eDhZ7JLQls5j8mvImt/Ur3tZM4RbSP0bHjKHWSy+1siZI4NQd4Sa8y31Ng
3IQcDnpURRbUT48UmZTo/P5Wm1+/i2znUNArcmyOWaA/F1E/ES5/mLMx75LzZJyGvG3HqAMcWssH
H1tDzXsekvH3q2Jjsxtj8XMEBUg18TRRtFObzTY1DyxJql9ezIC2khk9qRznEarZgRw2xy1JvR52
5HR3JE75a87xNsrCt4ablXX4+NlnJ+giiyyEwq/pIiiE5p0wyhifW+tF4UdbPzyS0P/vw3tCdWwV
kh8VqD/YSLmSd3ezFSc+a8WbD8y9KnAMHQo/0LvCmP1kLyu+hkRsWq42BVAdr/Z61eKOUGM2IFdt
yOYvxR0lnoRxgC2/3li8O+Urkf9D+R2npho4h/CBZprUPxyvH3RX/8uiClEl8es2gHWcLLOJ32k9
eU7mF/hLvuJrAJNWrkxYuuoOnq92XPW2cyH/KmGrVReMmtciMFL4sq7LqoV2X7P6P4maGnP+sfTV
in5eiiklaCThABT12gc6eZpEm3XTUyslT3vtoO3YYVRq3ascEGQ719ER3eua0brpna+mzHtXfQ9Q
mZgm5aQdzn43tBy52gTTX/h8rfX9DOcrIYRxKVUBIPT12qkg0CzGCJmJdRL0Ky3a2qwzu6NvhInJ
XOVlPt3DrTK70vGCAVrV4JbfEqOhd2lDRWppP57OLWfWf/blhehHwVJ04E49qsRdKE3FbZST4E2N
QI1uyC+AGy6UOmJ19ODVkyvI7UOc0Nx7hoN65PU1fHKNcLCEpyPrAQUzNbsL0NGxZaQD6lef0E87
zJ6FMkPd+DG/UT0DSmqJdBPWwZVfq0cRYsoHgel3CY+KIM/c3L52VSYyFeN9lSeEvzEFvxjyRvbs
i1sCDH6KLS/ps/6RgxrCWB0l1mbf2YyQ+DRF3/9Ol8dEa/6iqjzUM3oTQrdowKTbM1/ta3tCvbqN
fhGBSZcrdSsm9URjThwca8ZRyd1vtQHsRl3hHQpsTDLu5/9Iqc2MUb/cxLNZjq9CcH6xx8kMr2dO
bHsc8eEphoBknSvhB8KvZgSE6lHk6hn5SCiCDPOzKCqEPm3E2dthMzQw9yNGFVoOGfHCm0Wfjlnr
CeSqxhFZFCF17gjRAofKafbOmcnYlew6N3NXOlPEyAtSzrzXrljHcVCuAu3yYevR9jIjeOUvscEg
FZO5FULts/dLbil7JuVOqcPdXF1xRkqA/79u2eaW3nco2pRHboqLWZU2/A3cZQ0H+JmvYWXWI3Pd
N9zrQnzBdlYov0nbksvR6OANKkEiIe6ukwOS3icRvn6OCshYlG+4MDdX2Ql3W2Erm+y2uqjqK0wP
WpusOpF5PxoG4/gyyijJJxqRZbrlpkDZtJIG7L0Bmlf4k3v/lZVdOVWG1s3npv7oh4t0T8BCakXY
XymBDb7HkzMi1CaYoN97AJ3mFkUZPDxILM+yqz7LoULj/y9uuZAu/5voepjqHrmbcS30eyfGtRG8
E6FD2nlnpNF7N2auayfEMnG01zFNJsT2euAOGkSxxJM00zuGTSndPgTKAgSU/YLMnqeYHa29wnIo
d6ZUWTN3p5cZXQcZIp7z5MAKBZsXrSweBLLpd1BcBW8AE80Lih8DZ+zEy3QUP/bJ8RjYq1ZpZg4+
pCGM8dYwWpdI3OERYMBfGNvx6w+wg6kWesJjYBkRK51V9E8kv47TbddhifrBPEuANzNTykpx59mj
HkJRqM+RceDDOhNkQc4XNjZ/JXTjXPasinid+++yOly3wVJNKK6rHH0HiEVuQJ3Yw8MPEjhIK5qo
9ysirU+3esPqz+wdkQXqgOC43rH80XhoOCac5GhmWI2HWwBwTQpvgHJtUX42aGZdr3+HahA6qGnH
jqquiYg48GpHSGq3tjwgpczewF/INQ8bp+KKzoJ215HSDPwo61vgGp5zIUipUc2dVsRljiiyXS7P
yjI19MFUozxt77gXVkTXyAORkMgjKvOn9cC9MJK3CxF10dHFLwM5hncDKOBTZtvLEobmVbO8V0nI
sHuIAiRQ82QFe3WrTsFNOeuhfpvrjsGQQ39bgTApFhD21PPP3OeX36Q1I79dnRNZKpu1jD9riBJk
un4MdivDMeGEjn2j4OHnJOlVZOE2R4h7WKWGfu6IIb2GzTDadolsmyQE1KMScivq79+1EGHgdXmn
xQ/8qy4X3m+DKw1BIzFckejYF15SIWX68hcsRGlIl+KySL5S7UkQ/hU2pfQWo6xz6zqLFXviTvzx
Taa/NIbLUFs3e71D88R8USKuIpNNJqwHP/XeQHBUKujDBQ2Ra32Fxc0EkIeaKg0ICsd4vSTv52Fg
tmbF0er1CzVb+Gi+IJr5ZLXmCAov2e8pXJVzt97Kj566tC4d5eoacNHgnsKDz7wUvWzf5lTbFuDS
OIfi0jAC7HpoEVisZ9OIROcDBSGZvfhaQNwSDKyD8+2mlWMZP9o9gAz1bGRk6XJtFJviNaohh8yt
CpjlTFylVhbva82Zgr54eEwULd8sxTDXQ7IGDUoohJ+IFTNbEspbTOgk4wipgifShbnIN/xnVQ8N
V4VXBqGELUjsZA9eV5nAmKE2y/yEQlRNAfnuOjyr7gN7FDPstIBCG2ev1s16jdw0p65kj26Ri0Dp
UH+ebi3rTW0AMUevPURPr6s9hsglzJVWGb8Vr7p7l0Bw3aioaH9hVfXnUsQpBMR83NKoafiZX4oI
qwrXWkBEoolHurI0sKf+BLotP1OQEdY9iJJqWb7YTRwbCoA+X6PND7Gy+e2/DSpejIEea2hFto6Z
TKg/2WHDAQoItJF59n9EoHzvytUpATSSL6O6d0PG01vZr0sU5OID2GW0dulm/YF6a2agngZcADst
cU7OhwVrm44paxdQ+BeT9TCKmlB4M7oEIriBm6G5tPcKsGoCF3ABWsOaH8pfMFBnbh3c3n/D7taU
nVcaWcz/EzZOOwm1rJXzLg499ZklyOnROfaMiim3gLcZXktTCd3ZshQ8ZcgTig1MTOqpp1UwYIDQ
5kBnFuMQowhM2H1Ca6q3SSb2rQ5HGeu4Wi7X6dmuWDcgFZWBHV9hO2dsZvHQsfdlvx4MzV5OFee6
tf9xn1MkVI9UKOZa71fmpnij6/IHWbGxqoVZyyNGI9HkJ24LvR05n/gvoRuK3vPmT2KqaRDdRGU2
gH5Gq3EZvw5MBG9JHrq1ixZxiOuE5vfN8Pm0TTqf721GPGM26DtUh3rmdLpqbPURMzNtt+sT3jng
pMkWC9e30W40ZWPgdHcAOpSgbf+9hCnQ0gwEA1JK6dVpdYysysdaourpQT1+bUzZKdPKvEiWCo7+
bUYUny89TgGY2Baq6Zm/YeBGZFzKemVfUavo3jYrdPuXQPWirZjrEIgSV3rgm5loC4dPfXkMoiAP
yCIo9Y3qLdWPHH37P4qhZ/qxM41nUqxbXUn8j6K3eZSfZ42sae2m7Xe9Tjrf6FT7aIPgn2n0FeNd
VQvP2U7AcHumQbMUTbFRMUMCVhepylfWcmdJUL0o6UgGaBvIu4wI+fA/zQ8q0KND8HNZGhDIz27w
UisRnkWOFjCCxjtakIGdyai21aclYSZ3BlGl0vN56O9rGovDxRF6GTlra+IqXOlaWqlfdjHKeOoS
yvp5DQAMj7XGs4ZphqYQR3yCckTInl5IbRaNqbXXm3GKLrl4EDY8naHTGAX0sYlqir+cisr774Iz
S6UogRHO2Q5+1oJ0YGVuFAOHkb4GL8EyCq2GVATWQv8GdllkRVwCh/yjCffz/fAxGgwHoqSgju+P
ix1/0hGuXeLRxHDBOt3CVEllv4QaGjvbdDj8kSL0bo1bFLi13jt/7bm77BGLU7Btwko9CubtXHTP
w590MA3NZEZeyQ3pEHmKXzdiErsydvDihVxnEDPphxzs91m+06BUYzQNmB51Jv3YlOkp6qrjJH5K
zx9zBCnPKSUbCoQ5HS8vwMDQAa0IGeF6BsQT/LBwrTazCoO14Ao8wFK+aVeR0o4JAvRMp5937GLQ
GwRTvSAz/ey39P6coqGdYn7GUYy53qMJS2FnZ4uUBo0b4hO6lQ3icXjMfbZq57cZxXPlbtJj9ZLZ
hiYDh3W0WPnFm63qNF5PG2tRutO2yvbvFcWlqZ8fFfxNoPLo7fQxSP1i5wMd2so/9U/N8qJhZp0t
gUbeqYyBBzB1VPkwqKl3POmz7gDKDUeOhsBX8avz0eUlFq4MVG9jvmwhdiNMRD+HwQyudvlxY9Ev
h9H3MThwypKesGWgfzzRjFz+RcLRF8zXGZtdexdUCKMGUcelHyeP0NmtwSqZUbGRPs6kL2IXVJzC
QbDGX/mOXAiUFfLwEHhYvXfwoVcuSJE3/kBDofVf+YXj3HK60GSKXUcNSE24/1meTQs05OIlg96Y
TfwN3eS9bHOEaVDzcOHi2KADAbRyFNSZpldOiAeojBocCLHfiQaTbvXTMMsBzhXhCSWQ3oZMsqXQ
ykvBxieAvur5l8DIPAO4Znce7a0AJisVpgYhfCFd67AvinIjefGE+QqmjQmTsZocZV6D+bkJx+x8
GSF2sEFDMsBSKBg6ZvbVvxmnXraxJB3K0Y0iN4eJmFyr6qhWXpoHWwz+k3ItiJHywuVk7R7WdVuW
DEDAxu1q8aw2jjxP9PNS8TB3C9TxYrBTwhTpDLuregZoUiUD0E9rM0kFo/MTQIewMiIseGbqhPcq
1GnzK0/8qi7seRv0dF3Pp58ZvRpsuLuqaof4bPnQ361KjAWbND2oCaVorDxFs4HIuVWcMsmK/SIF
Eal7wtFBm/1UKEnNEMP+CCSrFnMM1nfBXyG7rqtvZLIcg4HoVtp1e796BmCCC2PQ7MeZMSpAabQH
jFA3Em52uW04aVVDCW7QCYSvevXhlAuDLLPcr3yE5ADyEFcKqEB8xLgV1KeJUfhJ/zzXL0bqL4Bh
TRKfmZxlbWMIQOAJhWFPM6QchM1k7Wf/EC23VCgi068YGa/UVzZY57CnzyQUHgDIZW+x38XL7/Fu
C2Wd/ZiLE2jLu7ZiykzF/pdE1J+emY7tVIA/oafXH2TYZupd3dpOiKdcyibulBMyaesUZFGz3OBt
XRfk5/1AC4Zeu0EmCGzX7KVLRuQWlaI1KEpbL2bw33uR3V6Nrzf7Lpn9BnC1KtkqqBqN3XGtyBUL
KlwsJ6TNl3bb5/sdlvvTq8ILRzhs5DCebIc4jiUVdbhny4liT85xCpca4dsIPELA9d5vmdItHG8w
OCk8fbWQwOLxVVtW9LYBi0xlnJhqe4QkilOjw4SrvqW3FjgH+OO9UIDzUlr/4JM/Vu3CbtcEsQt8
QWrGtEd6p1nX3dpjKAoJEt9OMS/tCKDh2UZH3ylncQkivvCiOph3a6pNwxSRggK2LJhGPsRkQ72P
J++fXeyK0bv6TpdNHrGgrZE+/hKRlU4a4PAhdttg924xTGEWFaMhxLCND9N1U8g/B+ouO2vXTi2G
YlbKfLdKbuV8hyKDn21H/YIlrN4haeuoDAnVEAje0qd0jZKmeh0uOyiDZeYIl4KC7odxBXIjJde+
4qcXj8fYBzCFK12q+my+uy11gzj64vF3siwUkeNLxNUGvJTCNTiQ6Q1NHfVPsa3gee/qwBlnIGhy
cCFeti3CNVP4DTw6cmFa/uVnV7I0vJ0oHUzp0jxaJvoVHZJlJkeVi9tDh9q6QQ+IErg87yZxYeJo
HYR4ao0MpAJeqO9KHHLSFuqQIOIXLyuuAcUy/ETiRaYwobZY8gWP6oWjxoO9AaVHpu8JNEaXe2B3
0i/ZHoust9PO0SCAS/sQswvPUDItMYiWQlKB+pzCgo+05gqZQ9BRHaEP34XYx2UcFKWiVrQBpokH
5iCbyPUYqNW3gIEN/01FeerSwuXHr9WkRxM7Wk8DsCm6jrU2TqARRi1MtpSqQvsa7MqsvedCb9rz
tDE2HlzRUZgsLwkrYzut6j4eiYcvf91two0MIMYqUQE9ttB9azJ9Of6Ts1CuXV8QwAL4c5Bal8nq
zQBJjQ95lAarCIaP/hQeG2/yM7c0y4R2rNqQgOdp9EcN2ohq07SiZajyQbbZcud4OUAErPg+WGxX
NRnV66LlLU/1Jnru0tDM+AFKs16vHsRm8yGDY9PoKeKCgpn/tfQVyVbKZNWgzyJvnbSFWAax6vEt
uEnHF5UP9ACgG5aASUb3K+f0q1P/c6/+Az3cT9dlSH78PWxtZ95eYrIMjQa121oK7LvI8MP895f3
tIZV2q7Wo/BUEE95AR0Q0lc3zY1tQoiorpMCgec7tzx0mcmMTd/rYJVP8aXBSG1ht3BJ3QYxrxAE
SmbF8nGPIN2Rrc0uWfsNTvzahHs8zPlNnnL0gnElAxm4nPqIpfZ4lEKodSwvJDpSOTwyq36HYAJo
GbY8gnKx+7KRa9vZmnmdgKxNRblerflOkxXessAiebeJ7MmTqeXcXY0eeTEtFK0V64DSiyZbzPEr
9ext0y8GMWFLq9cPQFzUo/qYmaTWAr6BFIiplXn7yiOFPZhNq3nr2y9/jj8fhVxEzb9EotqERS4Q
3IsHSE+xz2M9Frs0gV2Y8S7j2KZ+epyoSbx6fdkJP0gnC3qYHWX/t2lac1QCnH+b+kQNW+WjU9zN
eBDDaX/VOrKwyASfMdw17Ah4N+XJOwyGizwhHWh5hXMMWx3t9spJJZGFwFbJYFTRdg1Z1f1Tbcc8
AAjv/cE9acOF34x0z9oqFFKroWlMpLBDiSFAFywc2abEg4TeKjzytob60jKLe0+lP5Q31X8KZL2E
3wCkwi8wQGQjhoxxHbjGV0tgNGV2hzqTOLEBEuFFaKQVMwR1/BTQE/HYaF1h4ixkVCK73v1B3/oX
KycR6imM7+kdJvcUlMMPx84QNScNjncfGWRgLuPCI1/3nM4XImO2WsUV0p9ZPvHxIiejoM4b6U7a
2wMpnKnjMgWHpM+0jPYcGFHkckibGBNJTUw1sLrNlE2tDhGAXjUr+1Yp4UcQLlrs566XjQfGNsDf
gEWLR0SIXyFcHxgnTudVDHDYKzs2bKQQICIFo+DTb1gkpl4DYLVwA/X5RSXoNKdoyEJNzbA85c3w
LB4zjBZKf2J8Pj2IUXVdUmYGIclLT2Z5hlfgH5F27qxwXOiWggbSLRJaIllu21Ra/bLqmZZWtiss
j9ZKlKxu4vO9iz147rXzOoZwBjx8LPXQMreGWgCe3xitNYwJVyTizacCFAYgH/9y4BVwPkC4T32R
SuQrrD7MrXRtsvJqo+EK2lsm7AnHAa2fAXmvD3N7sbd1RfxkMjs+mv38nLmaM5oIieZ2f07MDJaj
aoQmtrXXdjxu/yj7Wxf7FM6WLrtD0z8H0h7OVg7Si+wlmpbd1qKZ7+GZGqmy42jwmBl4AGh41FGl
UBLqbTOzkn+chFpe5IKggBzqDYXn+79oAhRAb4PX7SDdsW0K6bY7ApFptmCsy6JWEU3zfJJcrh7K
Q4axFUezC0oy8GkuNrmqRw0XPJ7mUI8v/G7jVxXAXo6qvFIGj59HbIgyJtxOM5IYObD3Z2p8r34/
WkPBINwnvq+SXDva1qkkKgDKe3RCqsPP6raVJxao8k0Lg08yLe0b99JWTIYu8KWy/SMizRi3mAiw
BWYzCFqAbEF6QmY0H+Sql3SrDUdKSNRpCLCneynMx7OZ8OGFPspeDTlzSW/PqxHK7QR49jrp5a2p
fdzpddifc54KfXjlw+XFFgR2P8J06JZQXzquzkwXQAwkS5LoE/5D7w+RPMzFe3XdiuDb4O1s93oO
Z2yJQqHyJpk0lCd2uC4XDcsDb5J4iEFEnD02QyHGkr5dLG8KpD8oy7Lq42kPfT4lZOxvvmVpgFxX
S23nJnlt9MDoMgJ1K0Nvu5C0WRFrWEdrnwVUlmmvByzrJVYbNxlAKiP0a1TNJujEwsNtXouuVdBn
0ySD3FsB4odu4ZttOhveXZ+odZIxIDKMdxhEKaM+MKHsmPWcszNYOQMqTnDL6p070akUKjObSOvQ
rfKR/cpWqRIdsZiU2gLn5T7XW5WBJuFwn87t6DSxdUj4yXieTLRBEEGVcps9YL+Lv8Rr8ETwL7jm
iNLNtjQTTcFoMAWvzFQ6Z57YuHwb0iy6Afgp1spEpPCM1sKagvVvp9hQcDBgS8QP07G8LFw9YmxI
TOOtCIdWIndRZejukx9rAv5Y1wHdGcJ9vq1w34lcf+WHsyTqjsd+CMNLNH4bqSQvn5hOD7xHEemS
eaiQixuXzheKuC3lNC0R33nm2l5FldMbjQG4Y01jr7YSitOK+jODxTaUGqniEQL0WNEAx2nuHxfG
zHF0f+xJ4RAY2oThtvNqnAq49YF6/L2ZPySK2645xenmDYZkld0JlAqCcldiyb18Remuq0t7yuEk
/5+oXq1EmYPHXXlalNLWgsJ1gCKJsrEu0neX0pZmIs3oTAR6kRADLDnYksh4ZrGSGnr3b5QthI3X
ueSzAc4t8Wh5mSZj8R9V3E22cwksube7YSbpnymPni6tctoOqDdSnHVFFW46JkVNErvYR7CfleJR
PJSZB0BJ/0L3GbW1KPyoYlMlMxz/4Au8MbQ+D1RIN+IRLj0VHHU2AYZsKUrpjJcdqmgPIhXjqhrY
yArAm9C+0VUsvd4bKPa66MytyU0FrB23TRpHWf0LrIiMGWKtOrPPBgD8U9n6E+vdt69b+vKJTshl
XiJ8j/d/c3gRa8zxMvzN2Y3ZKgkoZd0vhOGN1EmByIfJ3LqpMxZgboG1NaQb1vdcagBAcgGqhGrA
1whhpQYxSY+ekSCElHXbBZZCkDq0VCiDMYVyL+9z91iu9gTGtKRwF9cmGqpfwikLERljLGnPpVBM
dhdpF7mIDpg6FSbxNvF6IOsnUvcywjxduYC85taK4ZoUUNEC4OwWRg3zU36gtVrNP0Ke2B1Eb+UX
qQRrdhaMbERdclIQ6Gf+FVzBPojbnaV6C6lUjA1BMZMaaNbSebznvtA6ojxuT6xPvltfYAASgDpA
KG0a9yq2DE1G+9bxapWPmxcluu+rbCXLFJLs+7mFrwA5gHUjElHJdND0NTSUNJl88b5rW5CPWIGE
t9TPN3dg3ckJCdXApqL2CO/+9WyQZ0mLUCpsuaM5J6zpesyo9knJTE9/P163BjP7FKx5jL8YSWD5
/zaiW3IftdI8p3NcI9vhoFApYuQ8177nWIKpuM3wWc9sf1TcDNPE1VrwJ0bQn6WaJ+45cphiy54N
nMKqAwWY9md3p2oRpJixqQp+Rh2b4mBLxi3o6jrwBBkUcGvCALhHQ0gDgMmJIl7Y4m8PUCJRLdLm
agWXZYA9S5N5ToYMhjUUfiiyAbiT0kD3TSrM1/JgIIiho8f/7kTMxOdUJjrhL02cFN57JfoX7xvg
mio/eTlgf1B4whQM+fzvDKsSF1DhKHFBKQAUsVprKdEUQmn/iHoeQjVRx85yzwkiEc2LgSIQNFYi
Jqu+t/W71yvfLrCm6i1pbH0kCM14Zvdu6bE/JZopgeWSGsFA+fGxFj3HSr6jqxWOA/3qUM9X5CUX
YmdTg7kgjQuCZC30wROMYAdky6YgV4JRgZIvLpUsRHesqcsUEteumQM8eBHs8AiJk95F0AljKKUd
7bYL6f1v0Ayg8f+i7SwvidZ++afrNJKwKqu9VYUqTeX0b6VVU/IFRpMuO3BTM3FJz6PllSJuUJa3
QHF/eBZVSN8uxQceaWOxKeUNxmV+Yq67dGctk5OnhU+JnCorsmcItCWvbQGuuV+zaJ/sWiPx7Epw
bjeB8n60yFNuK2m/Fo1RvWi+O5pc1Ae6U45UTMD9sUZ4vDFUKH8ynMtzz3eAwDBhdcUjvFzB0M/6
tGPQQtUdjUjXnH22gh1zlaZxPa2SmO+Vjq4OEDPDi36+ZuFoPLWKgaNwIg8wxjBaZ2Nf/FPzGRR4
xPFlEveike+VIJiuE2jYY8vuLmIsPYCP8I/LO289oIRslGO5WlvAotbx8gN7Jr4K7x/5YfCZU9GD
+K0EH8SAKNi7gVipgaFnmeVjHOpKHD6HWnnohq8Y5qryKFEz2hvY5mihbRJgN/8uGe2aUw/hOr3y
kRktgbQ/xTd+wjhQj3z9eoYMvkFtAIWBsJxaoyP8HvQ3JIzfWRd4oY3VycDfVAygmi+5GfIMkuK/
3bWYivERIM1pfcrW92VPWFFdZTX3HMvGZ6BOZBq1VND5oijukbBaKB1jrbBUb4K1uYfU7Gr8p6la
zEkIiObUrIwQpJ+V05qrzyWEQdtx2lpq/7uuFtEONM7u1XnnFM8UH1j81lTxe7EI9TWKAwdIubT2
2xP7Q2MuUQKtpkJ8Ar2ufbNiUN5YqlBd7oVhZ9rYqj2gHnDMrPkJPZklWFLwBBjBr5UibZ1fNPn0
/S9BsUJ/Qiuwun1lKEA8RDSp6FVlBobEwUsXuDeuuhG9OtDwcpWaeDWzn81fKdhjubDGRaVETteK
7f+VvHYLFbui634gZBHKgDyjyOM6sqoqw7WFj1wwZ2ghnAOY/wzqa3MJdTYxHu0AUOZI/S9b2sA4
uvd8P/dTDTlxBIExW/BBRVpcbHC2GS25Weg34gKKXqhfwMy4a5o7JyzH3CGMPGlS0nya5bwBWLxo
7JE0sU8vvFpQuOUi+CKCFMOJAQ/tP6FQOzDROGFHChwd1DNr5QKJqFIK5zi3p2MRn4NkACd6HGyF
bEpfjq8eba+ZcioIMxS3llmD11kZaj/ClLTXO4Dc9vhkiVxeRN8CX8mzUmKrrA3jIYw6PXOiNQQE
rqmnOPTTiVN6eQ+3tKtZe/eujIYdM+IbYzdWG3qyGFMPRWBKDoHW6w1OYM0fozdyceZDA7pBcmxi
2H0pxlxXNWT/xqw6grNSrhVcGpVnRQG6ukoW8cz8dIjJcp5d/z/y+n5/kWG33iva2cKAFMWYYUmv
hZRzESXYJwbUL0ffk4u+ktmM4XHEAcoOmOzccRxSjitYvlMnf2dAD8czVIRkZjZg3mfDOx9251hO
QVE3D90PiZow5Woj/nziO8uyOJqnKQ53AL0pIDCsp/+Ydq2XMRkip2Jve7JkH7y/Gcya5WZ8MVcF
DZnQgzqpC2nYzXaEqI9lNnRUN1TTC/aH3XaeR9hIehu6W31Tpq/Jn3THiJidYKNxsn/KZW6ov5sc
Pfd6JiRzBEbws3BjhBCqkIxEPGtoWpDth9DLc1WUDjOLEzhxUP9HiLEDdqIsjMH1kJf228Ae6Bk4
+i+RifKN4QJec9aCBLJwvRL3f4V97XVU9vIHxEZwow0V6gPXc5sc8oq0bDiQAmWm9jQKp2XRIxcO
7fH+WUZlBA4PSS5KSeLe45dsaf5/1QPFFOEPr4kN/xUuHuTh7ull1ZE8r4B+m2vm16I7AfTZo3V1
UHeAZW+CpSOJxCoQSINzYMUl8y0TBfebFjN+1jkDCJoOxsujNx8TLkEezqZW7oPzOJqXzzkS3rB8
+oWJvokXYc8LDlK3NlG2tCOT3MnnY5aaFN0VtvXGGnD5wLXAtn1elDVAd+Tej/uwtVF1mz88oyS2
7sityVM/8rGoFzqfqxvEqhRSM2zZGuw/GYOWsIH09uwz22nKXACcnmTlORtBeJVB5RVs6eQ9oG/e
D4HGO7ujM5O02uiPEXbXJTmbnBn4EqNVbryDNpe5dzBwFdrd+FL8wRHJ85JbY10N7X+VpKsSICun
YHyUxwn7TIdYaOVRuLHwYF27549zDEg4HbMW/s9x5pU859+W0rynWo3w1UWoGToDnhvVGyRE2ftU
vd94UY6hF0hD1pd9/E0XwGmaXfCDZRYZQ9l61zhKQk//iVv9aBE0yG1hrp/rFpSUeK4UxhEGVL60
aEDuVmFggG4AYCMJNu3gtx7UEYx8MdXF7oPgxQsuPrWF+hpTZlp9aYWG7opB7bV2meaUJiiRlqWX
4LMIujQ7gsv+ILTNr4I3W1qWnT8sZOeU4AVKkMAhkAZNRPOv4tdMu4RTe6Z4aINPEmxNQojCpc16
Z7NTHp/RkxAQCgaKuZaest31762hBoXCCljDw5blmrMCyab3JRvQX88DshrGBlpWbFh9+ThjSd/H
RQE5rHeimfEONWvL5V5d6vtr/EfNWeSoZNXQ8qTVKOotVzmoTN5tz3tfJU8HZjl/aDYBemHS8vrQ
q8P8i41qiBZynr4XQr7R7noVfmkpsCPTbgi2lUG6TSkJjqHtUeWGIajMvTTHleFiqExQoyQevrXD
HiR1I7Ayz/sRO6sGI51mZYz0dz/mMGbYIVtiLh9HtbsHN2VROufu/1eH6QcHpV6/tAb4cQvBt+Fs
A8CAeQwGGac+cPQWzCfhjxXhfD5fBc9nonZN1c5RTnjJT4j6rB6fXfb+qzKXdxdJHy4X405FwizN
ayn5a+wl2oGsMk9JpdISMflKcCR++Dhs+t07hHm7//1XzE+pfFveJHTss5zEN3onWvE64dUYgWE2
T3u+17Ps+3YiyjIWjotD/5tZm1yLJ4c6LdZ2aR+NPZO2HYro10LO/KCUROQDdaECLpEOXOxA4hRa
L4QjtZ/xLRZiyjouglLaMPWqjUMzY3oUdoZZcfDrv009kM6MpqJiyi4OLFj8zq78BsrFPhXXZJz5
xDAbzlfmKsEOlhBPQRSist7XAFZM2H1V0d63DUF82VrVoLpnuo3YaihdqnOMeDtpqGtlTspMFAc7
dsTf0PLyQoUDGWKf7gUK1+Nf1iqAMXP2FhTGLx//vtXyaZAdgdlYmninQuQa7HP+cYxB3ddzm5vb
p+GyfCcMz5HE0PjXHda0hVRsmn3EFd5/n0K2qoK/3Vw/hqIPAQ97srwiirNTifqckSFJDme+IDVx
67S/95J211Z7XyqTnEN8YTqFCzfjQWZxUo4ps2PyOaoin+X6LtOSAi9dXxzDapwODHCDIR7N7Dpn
+S1sFGkEkF9rcTF0Woc4AMipJEyD+PAVjfdQxZcy7PCG9IXqAeCOAqQ7knjMjPZf4xJjhsPlTOcC
faBG/7k4cnUwlqPtme6SmlkdYYiIO7xN9eTB7YV1UGsZyEbwztHh4TpTIlxZpl5zEgyyzEnSOMOx
x5MbFsAkoHSC6j3vFjj0MUUPXepOX0ZdWpRR63uhbMoAkxgPcoypb6qErVXswzsKxwgkZXCEkNwm
Itj2YpMbJnS6I9AO1fOw3Bn0EbecFvu4dJQeF7mab2kkIlsLqbAT0SATRyFyiLF/27tjhLPjauXE
jeF0qSIy4P5HC1+KIcfljQDXdkXWju4+mHiZmQriYIHpGBAzmGWjV3Ypa2hJog7b2YYalbecoUS/
JcGNTJQXMVoGh0qOvaBfNX+8nTvDbnBrVkkGIXsFN7zxUt0COml4zPstiO+V8WMa9Ua8uRbkMzIu
9D3Koqeimbpe0UBol6TQ/dFFvL+VWyh5TxYybJTxPySsRJ0q2JtRJjdLUhwHglQFLsMFiiw5E/TQ
wuaslQAIhNaLYgV7yjwUV5wVCqLGEF068GtWrNRoEI6BiFVg5LHWMmnm1erBt8/1AkjA3wq2Gehn
QDoYvDmrd7QxqY5W2YLbi2AOnH1+JX+aC+VlexBCOORo6cqXFVreRccM+GOYPto8ZyvCg9Ishhem
xpKZhajgx8/N8qDCp8dKDMtAlaUvsRf9UP3LIMmT2rflhZ525SzuiaUS7hb8D29ED/0nbYMqjG5D
Eg+bwUcD6bNK9r0spMSvuhOy924WKSTzcB3/VWw+P1Z5wlPG7S3FxUrjFBU3C9CjbQTNIp37s7wn
HzdC8/AtWQf31qjaJfgYV2J2xvp0Tf5Sj3yQnjuAJY8M1RTsRsxLnarbBEe/vURix4HNwTdPdcQk
YWtQlY2C//aSNnu2Evn92nFiRdGfWpZW4zMMVXvdMbJ2Rf5gBRrXf/m8WLv91mtamSRV4QyVE/Ak
zji/PyzyaXEBlw1MXve/IX/g4tJi9+41FC6bcD3drKHfUf1lnW+T42sXQ4b6Fh/UuhKpKW+BcKDk
lVrR3gtO7qk9uhdMOWuq5ZeSgI7FZMstK9q6PQlV/zYCVXBfn2N+k2KdPkN8foOPVnr7vF7E9mq1
DD4//iwKTBaUaCtDBl6Efns9sQ4zu2x5ef17KfQDRqIuhP7hkQopPyIioNQpnLGWneky9z+OgMiE
b0w+TufHv2MAUvm8eUnrqnDAcrbJsGie4+cXJi/CvaXlvMDSWAqPoMgimd7EP91+MYMBzSS/FaHU
bga7yvw2beaEGWURDIcFMwPnbcKXpsEXjl7qDRqcRm/3FigH/yqdgEGB8mHahysdfhVSG6CnaI+L
dVy7Le/49LA6MtJVAVpT9G8EHLNmuCvZgikeNwI82InfgAed7X8ZeNk0wSfUjBno6skG8ufv1/zQ
67mAdlmucWar+1cwDxYjTdUp8bTriOofoBoGMgvxalY+diC/3WSXcRMsjvZjgk5xmyL1kUPuDEwE
znPAfms1M1NLJouhtCZZvMjy5WwNSQNclFWbrDjZrgrxvyYot9TiJmDHlNhnHPgEdKadtDYuhlE1
qHJcGs5o1GT+b/3c5B4lYlPx37HelpwvixT+9pTM+tPA4SLLbDygCmDeDCvBO0EmENpS8qLy+u9/
Z1uNkRoEzEWARjk+zvoaCaFT+pTfY9VYYE3feuiUh1OG1uTRpDgwui3V5iIoVJy6TIFDdG2JUHBQ
yN6uLzaIRmSMrODKP8Ji8nPOQmHhCwrTVUX6FgKjxRxefuDprtw+NdXSbCqxNWgV7Vdqcy0XL0Mq
NNvET4dMc5olzU25gGsZSgM7k+lymCqsP4VB1qlQQxcmCyrmpvkcRQgLpFgMfbiyoFABwEIKooO2
tDUoIdx6tFujVNqio/7kr9h7DLuv3lbP7FGtkM97wVoMQvHBCBi+2H6UMivId5z9KpYspqQoALNp
lkNnYyqf9PDYUS6N90ICzf/yhAqWYtTgLtCdFiszZ/oyN4kgyavB+CphsRi7yrE64OmmPOMEqQtl
gfQVh1STLVfXsPasoSEjhtLN+aRR2kiOwI7cksKNUDAGe1Vv6AgDGmfxc3A0M5DwEykNLZN3k31J
1wEV8ucNsNPwALBD4TAuwmsE8vL4QcduZiam+7D9jaPxW2eJxnvhaotdBVGr5RaiMTkhZxCeOwT6
DPP2evxCADc6OsKuwgR0yM7zjcD2t0MnOCvMhNjGDwI04qLv8Gpb0/PIWCCm3zzNIgZlYuEVNDFz
AaIHFs7ZHe7QNRupxDRN7pxRxR8VQ+EVyZmCvtEIxlOmP1uNn3M/Tu/VzOc+RO8pHpIgsxW27XLn
s/rU3PwjCh3ui8hrWjgDV2orq55fqPXKx8N4ba0J1208YjdO2fRDwoHjHwxdnkvf+f++4mRp54eW
ZOzAur/7R8j313Ojt+wGr2XAolUnm6mDdboTVRH1ZqQcHYovkI/acit46ZH1t9uMedRF6qy6Vmvv
YCh+zHpxIpUrc9qXyL0f7qsbsFXBwGQbJlWsI+qcnwDjaxas2FzaOavD7z02ex9ERsVO08rWngE5
5aRX0yIAbtQ0ql/QIlzM2viqUfxkKQX6ykf++2pNcmpBN4fic5CcVLHkLNhxags/uyPhozU7V0Cw
9fPR6qA3Tzkrc98HQNBey7soHWOiEJxvchnMtugymJJRLmYUCEFJnXyJsjUq/0WWUfRGym9AdDOa
tO/Lc2o6Z14Se0BR6b3jxct3my5C0NdjVy4ATb+Ol412MzNhAwh3osXnjKQXsL1vXiq3deWU6+Kl
Pgj+ZypyqzsNQof7JTGdGErSeAQiwXJeNRBm8XlGDx8t1RR5yN4o+zlhIDUo8eg7AqemECZLgn3o
pzqoDZ2OXx8PRUo8R2gH9WsYjYt3OFjwKrXOIlxx+Wn//RhoBNCw+8IzzoLzER42nObRU6uelyg1
gGsRJMunRCHvYbl+vZ4CWTLQjImbL9b4KoK8qLHex6Ssm6muThqzM2p2UccjPCxwJmyPzyQZCsW3
lHI3TMjreKKztk9mJ7ZQiZ9xGN5/SNBzoCarMzduCimWXtJ6XLLUlKQe3kFcurpoAbh3HdIweCYm
+GmfXVaqvGj3aV+NbKVPzfiozqpYtLnuw8tBA51Y3N10hlZpdiINuZCMOoCqGhCUOXlbUa4Mu8Fj
kskcTOlRBDMSXtHvbSnbUv7zZvRAMCAa1p0aJJiGJ7Xb4t9UlAXMT7F0RgHVxleb+jbnXRW9aqg5
ZKycAWf5oFyUkriPDtd2DMV6Ky4YO8sAl9BLEsEBBnAm/vek4Kz+9er1Z9yn+PgbZXyG3gKAB/e2
/sGknfc+fNdPddHKcdaUQhd9ie5E6s9sOY6eTKiXYIgXn51hcweCF+LAztW1rA2zXz6eavkb2c8T
biv7e5RfFuS2Br3jyqi1kQiUoMv1YNmN+DjavxmbiQ+1qHlqEzaf3zhi41x4jAXO2yLIxQCXp31C
yWW3NXkUdoX22NJXJQ1FX/oDEt1J5GKLHQOrdx31ReHFDnaxLtS8Ebx/CWrRDGO7XFXhznaha1EA
XJPoP+FoIzIgz0OOUTQl0YgGXrEldtw42FSUVEd44X5eox/CejKgbo+l6W3apHpb+Y5ocmukXiQm
dDxR5K92XMc5ov4llnCQqOwiznYiu+45tKvbEgKA/PP8x3Yl8qSd7d5i9ViwNJb/fGh33Couyc0u
v85AIRZ1VUfINocRtUPxez/xGqfwuaYtkbXUjzUPOdkNb4QPjX8fs8M90ZZYTkW6T2KULxooZTZZ
9h5nzIFokWXvo16W8DiwVRpFV5M6OQW8+I2GRi4phU4YaeA/WHJ3DhMQ186Xrq9dx/kRAHcfq63r
w2m3hoZHM7lLW6B+MpvWu/VLFKtpewvQUmVqCnmMMNRuCbWsqfSebqh4csV9lC9n2NNPlHWZwb8O
XUA/zXzol08BrpjmkElQefcUhKhcAE0QXN/b5IPWzfb9O0Q1fTLaloN7iLCP9WpsOXo/DKsYmBVt
cHuBeLSq0Z9HP5OYteT+wLwQwN/iZq0XGkUnzqXtQgARo9GlnBSFQsNE3ecBu2caGZPupJafiQS7
P05az9V0C2BuIeS1giH6AX/+98mPTQuDBVhsbS44AfoKcAZ/nPSh6kI+NRITbDTpSwpAWhSNiwpH
JBoF2JRS1S1fuKxdAOSLWRpOON3D2P160VDnieqK4pPYLqlL5PuR465P9dkdRfCdP73p6YKC7Yak
1ijT2sYZaT4dLlx3ws7uq911gYJACjgPWqGuuN5eWd9WMtcGXNtArRZp0kc3kNWAxQCBKDiR/YWq
L+EYzo3tSLr6M9HnEZB73UDUd2Z0kvjx6xmyFpQbt26F0l5Ilyr/P7KOgTQZ/5ZfKt4sK9DYjnbY
UxPk54bb4fE13Hy7EBwUJGaVygF42szvnvl84vaA5p7DZpz5d9afNPrBI7i3vT15eyK08yLrVxOk
mjNEiidf9aEPuME6nIDoXQFg9nexvbRcuwqu3dhq35wcJTTnoMv1dgkarU87A4ixYr0TGKfrriCe
sgiVIgJNRHJ5ueVqw47mUkRVCCgpDRcR5DYWnIsoAn6TYdxkL5dSppUGqKlElML7TnHqmbiiF7C2
4QKf4IFbVYFZSDUFEbeY4RAVZ+QswZ0V4jdQJqeMwQEFCmJUH9AZgjue6AuZ5AElzkK43JOk4JxO
0mYTaaO65SMV7FxI5yRtmaKleg73PWzH2OTgmWsRpAMKeZ7mQWsvDJu7bpvbwY66C2sVm1+zhP7g
U9uc7VHoj7ZMZwIUzDzIWAi4vj0fL6irDAx2M4+YfAI6vo7kDlsGBCxiREueXykVmKIWrpR9egOc
+fTRppDmALTV1DbVheO+t8zF8Crn0/oLD6fTyT269EZHDu9hLooPLR4WIQytqG5hvfu6II0T40PW
FtD0sXYpPzU3UMAMbA/SHo9VtKrf59JKbvnUWYWmz8WzFXb/gVCodqYZD6mg737jJdgI7MicY/mb
8LLNdsg1B0L6+TLoD9vbkDWWRbS14lrU2xF2LpJCTJysFgkRaHN3STZzFvn+zGf6+A0l+HB9ZJCD
5lNbm9N7GSVjm01DLW0Hilx8YTPEkMGHnPBaq6ALlPYLs3FTSxwdHwiVnVHh4YqecoQ72zyPj0Uj
NVG0cISawR1OSZW/7qEZQ53STZbVHNdmNpcx5BrjB/RGhahMeXC8G+QYAsKzsEVKChXTkD1++9Ny
Sj+WAnTTX2icCVka1cv2PRJxnEww1lSq1KBvEmYL5S0r/27hMnHaT3N1zpu2NOx88uMQC0FYqh0Q
q5Z8sedRZ+Drv0pJpxAyIXiPaowDnzSNkHXCn06/A59US13RAu+1uQFcuGb2vpHZMod7QWgwvaPh
DdmY9Z0tpqm5WDz10O1TIjCvLqrYyNoBSX1dQbXRRNiI2rNNziBHuq21lWnAAiauEVa2ykZoGFri
2F70jsR6RU7QEYrlAir7k0tidWu334iPW6yLTsUhGDgJo1nawWbNDnHPHIZAYi8XqceMTtFkpBf/
XwHkWTLXUsEsZfIy4j5xCMBn+rwkVj7RucCO73OkcH0qDqzIH2Kx6vRbyoNT5OI6z8AM3r1P5zJS
FH1AxcHChfjU2rTHx2SN8FoLxpNx5CdnyETMeHaA7dl/yOnLTiQZ2/2KPyJo2HeiyDzcu396CXNk
THuUgSRICLr+7gkPnrR4PoFRfI0ChFcYT5E5D54biXbLiEBwyYX4yKUs3ErlYl5RWIWZqf0sEp2q
dfd2tDX2Harayag/1/TH2545p7i9M4FHigkiYeirDPR2cyqY3OE9tU4SWmQAAi/Lka52XSgE0EgQ
Wg8gnBNiyUzowmY6twGARxlj7cLRN0+VyQrleihj6dpVkMHeuW0S14Gw+WCnyX4VlN19Mll51i5w
5Oxcm+4hlv3IVUNRjl1irhvvyRKmrhWmuG7UJn+il3EXt8ezEhLGMdNP5DciPL5CiFxvE7kfE+gN
5U0Tn8l//Rp5GDsiFj79tW8vdhWVizTjeHv/kdvkX/YtGHHwrfzp+bqbUq8M4J0RPghvVXvlc2SU
EgP1EhtuXAiR7VCxqNG6rMwc8R0Hrw1nEQvqR6axHP4ORdBM1fIkD7VcXL0TiTM+MczYxc6tVfCs
LkCOzCCpDnXO6wNVylXf01nWdAXIS2aY1XUd+mMArZkoqW0SQT+hPNhzhAQwluipyNi+VX+UWl9B
zy/hwQ8t4Lw8hd1pxbmLdicBoJyHKPIaNe9nz1LDFvKLQrQfSkAo0DnJmVT3oAR6x28aDCVnP170
1zMJKS69dkE7julB4CRL2XSB8sJ0csO98rjlUEZfXE1eQ+tD7hU5RH+/bUl2Zahg+q57f/M5/39+
nZPAO7skvHCcHfbODKCYA1D/6poExhHHSYsGweRveeijgUzfabPVbv4JWE3GbQB+21he+yQ/TJjv
+TiAUvHnzAnmdczf5v+9uFkiOsrHD3Wzko7BfHQl0WF6XRGc0fysntCy8ZOJo2fF+6abSbDSfbPI
jrJQJklASZhogcd+dnaut2k3cFkVEuhGdKROijs2DfDUiXUwHsnS23784ejkIXirOsmr16kz0xd/
NVdar/sSOl+XhJ3i6DhOAjLutePTyOhywG71NcR84N9qP9M+TjWE6YbTXu483+XwuI0giWgMHXNu
VIWKSeO9DzZxZDdHPORB2xiIJ8L0my695hulNd0q8x4zl3Fe4jYkWyjMoQE1F39JmeGQ4mIayghq
YTKJqF8EnxH8J1MWsQ/4jXQRjaJdGNVBFzm6thMF2iVME9MzEcpezIFXlmMV+kR0OYxGzmTqgqWZ
Ne7g/rjzEcf4K0/ogLs8mWqqzPNF8WTcO6euimDOklSFvu3KRH8WOp2tLiWfTldJ9FVxA1oAIVHh
FGWeV4R0r+KrfH5sFt5dIGWnueJkWkG8jGVhVq5kqY0DOcssqiU+OUf0CQ1MsJGfTqF6W9W++wH4
DaTB8QJiyZRJJ5cg5HGtonfKHa8KgoVGhH/IVvEoe3KWNypJ9YGdL30BLtaY6eL4SxK2UatHr/ke
AcBBRCBcpn56huPlFJKeTK+w96z6VgmlG42zyqMDkR8SPRK4Nkkpm9h3cERLD5DlwKhkFkRK6Abf
ixeaKNDCn3gADOUo68K0BVeOAH6KDDbYd3n0ej/u8h3DYU2ROguzJEA7hNCxG5Yt11e9HgkFsuoG
4TVJekj5jT6qJDVW3Jm1+CqDfLnlQ0682HAB7z7V0nJigZYn1a/GhN9cS5wYOge7s9Z1X+NOriVp
MLS7pov6cpqRSllbB4K8Rz+7uuWAf4AttQRPj9xtdlrsi/5zll07YCKZSbADdVUxiKwWV4UHpjF9
8BNJYlEdIiBVEe2qxg8J9XNyBhidK+OJ9SMYFrafch4mPJ1k+eTPzuOlXAVneR4MRFd3veMZv5EO
czOpwZRaNqacNxzxkMFGCCWYWFrf+xbk+Cv7UY6IQeNZT9+YG/LLVvdDa8hjxIJMYw+BraCMHGC/
v1tFYd6WVk5zq/1BGbh0vsNzul9/GjOymAPZEdgXLiBv9zDK6JtghJuXHpHY3jTLXKHQRgoSVOMG
1wpxvFNnSWRx4Gh+MMNVROR1PORqddES+S11rKXZMKXNC8A9fceSen9k1QlzCKhQba69nwXQpFhi
Zk1N2a5olSBfELvlT+cGY5wRq0ZnNfBmPgv1LyfpBCh4eOI9xy6HwN5yru5a5UWVm9+BChKdRHcT
xNKJMYlrJAr/DxxTgJVc/16jybXcjATBsmOmmxGDU6AbfPTOhKuWzDcOB2iD5vFk44/9/XZcMvut
RWc1ciTHqsqa7nmAS/ujMB9ob6dz/nTHGnKJtXmtpBEXhxld9UCjb5f/bMl9UmYjKUgINWMMPzR3
uDx+/NxHj11/83g4dsgBM/7MKgaVnLMXRihnhjvysW1lfkLoq0647qqxurwaYuR+mPCfWCuLy19f
rwx97OtHLHhBu2V4xPyG2CteGCI8xcOYr+7MhZJNIKoHi4CL3CT4x/LMTCJnvEOqKSGWkSzRiIFf
2wol+uV7U/w1ePGVbMGpi7VvD+Af3SQf0XQBo5ydRpmanxb/EZtaMgdizuleAEZLrVy15eMxTujl
mhLTF+rdJfZgQUZoP1VxQeG+da1dqaMEqrIdlZfVWGXpYbycGp2POEF1Ow9UOfz5CUVGnw9Lxep6
xUJVqO+MBNvUN2SZPeYKnL+7+r32mQiU4oOamSbH8qHjTqYv6uOScNBpgYnxMkemlxaJTWoI71oq
4//a60X/Pn5AF9zVcWmbf/E+sRP4n5AmdkfiXt7Wpji51T++OR6cmu9IkVxYQ45NX6S3GevHHn5P
sBanNvWbF7PKXxYgwXvaR7NmO1WpOMeDu3XTcT/5MZramJ+SLA2yju5Twm8M/SQ/PokWSYmaRc/J
MuoTHQKNXRGlN7GuJbGk4+BU2Qt+TUOrSBQAhFtaTatP2xi3ntoI6waDm62oca/7UXfDReyHezIT
RnH4A+urzLxx4oNwFk4uqVJBlRNwxmKkgipXouwGqpxAARPYkl2mj9wl4L6icT2EveDCPOXJLOc7
eRpGoiNoTWEOg5htIdYmW80Jpw4oh4mMRCUqAHoc755rXq1xL1bncTKX/IylRR91PeeFkC3/6koL
DfGXEj9cCiTOM5ynGbV4JbUaybSL+3KA/mmnxaSPOa06J4WY3W40yrMjHFYyr1FyFdgc7OSYOkeq
w3iASBU4qisIfEFMJg4VCA0+n2o6tHMlu9KXKSJsa9h+JHwFlnNxv6TiWEsknvy6vGB8j/wPBLXE
Ff+sEt4FvmzBJu0S941LW373qWk+ZlMRBTBfZSKRTYnR+NyFkePdUaDl1SN+vMDytnls6+cnzUT6
unkGEY+5FD3Oj715/SdXWME654IlSQa/Ts74ruzXYwMow2GgdeX85Ra00ApRwtekggvCx3U6zrjI
wYZlrFIPw5QjGuHOn2iTgEP6ahqBsQf6ptJotJklpSXI9PEwqC0R0wYQMRztGPhct++wIHuXMAAr
g2PDfrXdHoe+uHMhparGLJA8yXu6Uy32+J5OxnQYrdi+jD6POVavnFb2jh/ZWoocy9U+eSQAkjYt
M6ey8U/TnV/fa80LoHvFX6K7rzeoeuaE3eQ3w8W+0ZovEfH/5xRLapOWSFJe4/YBHdx6dzSvqOvC
Mv0jmqT5a1lOZZQCF3zBJpLCOMNW+h5XWKQHPpfzDGcSGuV1P9M/3PnzqcjLjOVOLmARJKr4HFVC
/2k0fha4A5o70ma+GKLolQPMqujLKh59+feMXg0h+M6selKE+jEM/PFMVBWZyUHrRAlYh46xHg1y
w0l0hzqW20Ex98YAlW/9z0nEnqZFrullzjeeGIcyJF4RXYXghlZw8Mlx81ZLVkDQsbyA9QVTlTpT
/XhZHIffiLNOzZSWRurcQROiMUknLrEoqkMXWmycqkSNC9z+6BPomy3BeNSypZeEkyA6lp6tdJK+
xzORnrAyG6wEjzlCY+NTBIqA1iIYDWGlNULWYUI8utPg3KZZpdlQsQuOo4jVWCYh+B++PxNiaBVa
IaP79LT/yQc4M49aCMRsv274Q1VHRxm20ZCu7mR7BAl30UXhyi9zfOhZInL/1fxGsb2pUXPpoUwZ
vPREtiyrP9NWP+uJnsn7frqYCX6cb0nrQRc6FtfYhk3ijfKCKnSKkanjMUoZLAxjYiY6qhULer2u
od7UTw9l4mHWbvktOq6cSV4mRkCnUv9hk1ai5Ktn9+LI0ag7Rl+Wq3pB7PJtJGIv1JDpeIl738XX
6ynzy8bwXIrB1DYYyryRUl+4g1h0JXjbf50rMuZDaZ7yJyDq0xA974qNj4/LNXqVyqQRKTlCRTmb
yJ4+lfOi0aLrCJqyXj2Sk2eeNtUyh1DLJztdKjpKFqmQYkAINeBAB6/pcjSbnYbmwCutG9fv20jI
b82C+S6zwi71ThuP46jKAlKQHK5B3+QhPynLqCm/QB9qqxXD04a2rk2eZjbRDYOABFpN68k1S0+c
h6yXytEEUd89Ynq2dnFbIP3vuAV9Ad7M0jT92MrI2yQd9bnKp15ndJTmw1uzwdVbwZYjpEOsU9+Z
muBib/v/3edPJQBy5wiaH+b9jm37m/E9yxDHggJ6CUAq1mNRWs8BRNQnM2LAm6edlGj1THxYiYPt
RMGoRsfuhiBfT11OhtAXDqHuWukwj3trXGXef3IS7niNSWMRlgc84S3ewdZjJZ1wFIlvdA5tjgst
BO4D8BJYT1mqKruivFyjg7M6ElE0PUuPsLXHmvMZC0PqcHG6aZtyiRXRkPjwxo5mwJI6b6+Z7IDH
q0XPVAjefbueJ0fhIZ2hyT+Da8ImjUu8qc8/U0+YLApUlKZ1jYtcxx+8WJ5Cim81s+5Lj2vesf1Z
PhieosXy6Oi/tzWXywMR1BNN5wJ6ZJIsLCaNay5bPrS/9E951vPvVV0EL7ssSRXEajU6Olepgq2L
HShK6LNpAL/Cc6si1lSjvKJZNjR84AJbmH/HPkTZJysgdk150WDqcAHyzEJ74Df9IMQI2Do6mZL/
50XIX9V2FEkq9iRE9K6l9a0sIXw8N16fMbi9MSqceQiawF0F77QC17udK2fSkKhasV4wFYGa21Uo
d7kDFtJeiUfbaF3myO73kd135/Q2ttYWm9Z1SZbit9dE22JIZtHKGPGt022dbwiLHKlPMBwAI+73
2LehSgPoyyhvakpEI/HXoBYi20gB7Kzyn4RIPYeD5Qgj1qTR0ego8y842qcPLwXX5naKDlOsTCbt
jH+FIkjqvXs5596kp0XX9lB1n/L06CmQ7Epm7ccagpy3f4EyazMFiOgQCApdYHcGTvDEAfk7KGw3
v9Z1exNZ/B6W+k/Vdlhd4CS7nP1XgnLHVcIulPZPdcF+RnmM8vTctoDWlRzGwh0BG7jkLksej7P6
ejwJCwYUuuBiVB61tyqoaTKX4uHvVILxSLTpyOa8PWaRfmsBMUIrHBQE65DvAud/24TxpOATjVnm
6kojA5uhILlSOBm8PT3h5qbJ14ItVVNvZUym9aVMbZMYSYS4me0j0k711HjqYOxqnlip8eJngR2B
gT7jdq47cGcN3ExdkvG2kQGlMRY46AFvBG8jCSlCng4KAbLwiEkMdF3PXq22KP2eYMbIf1vXv94X
IHqR+EAj0+CTC+h9GOJuvylC90snlsTsxeVF60Brem4osuzXgd/oJaHnGNOKKPnykWnw4jF/qx66
w1oyB+mtskgjyKM81suCx3U7JVvcpKjKB1p8nwHQmL9UQE0XTr4oVqK9+3MB4d+QUayw6+0U7i/n
YW5d26f8xX78v1ID5iSVFnov29uZbRpSIYxjGGI4TNEVHPMh2W82TxNUy7mzMMmxkcVm+Lhqg5M5
eVx1oQhqah//BITgwklgxjzK6wZH0jLKNVGtwIE2xUV9uj0UMsKwfFmMoJKObaVGyFmJjyNTQHTc
lj/vtFKWkJDYzC/+DK/nyfKyjncmOaksAxehnODs5i7A06nMtgCyik96MTCHLWrhNYyFp1Sw8zNY
n+yZ5r7TnyU0UJYS2pU1rwCyHzR8MzCs/Ce6CAvFBsbeaOxf16o3nWCg56GSuvdFxSb0TqQOdaqV
sHFruoZKu265UOSfwKRTXjy6joVjX41fCJb/ANJaeoCYRf99dZ8mJCMkwkLwhAfCoiRJ6am5hcRJ
lnA+BJzDZAG7hy5SAgcWkdY5wUeV8wmiLLP3vk9GmIRP9t1dXQUzVJ6AwLewe0XHyTLiD18ezsJ4
2Z8wm8xz8vBf2PcaZDyNx81xXCKPbXA0e4FIvzNR6AmSVrmddJPtHi+tsHt9NJ+BqZz3gW32mP7b
VFcj+7Kfe8V8wl64OKAp0U8JwsjUK11dQtBfCuzl8++B/glx4D/Sw3rhMk9AaQL+w7c9/kVXlwny
Lvb6b8sxDagYMWLpdmt984RyHPM9rz+/JFtIbjV/XKTJ8lO3U/BCrRiIwzZw3yZ4vRQuqfi7einD
F+uIruJ9xzMFK9/RsZS1DSLXNl6QYxYr02/H/7cEm+aOLmT1X3FPA6eFtUGzTyQE1XRPDT1TGaPm
l4PQKFdKz56x9uKpKeYEuUBY2/6/JwxXd4Gk/QUisOo2N/YQTymBoeJ6Ad207wTeaJ6qRmmyMX+k
KaxESASS8sY+KCXyJ9OVpAzkLlCL2KovECDgd48d8kE1unh4T6XyDoRjTRy73k0XDBzNTvhJH/SL
YwM6uUg3VK1LGhnp7PaptSQ0+VORY1RziQj3iEm9o+/2CYsbW7dAzmQ/hp1ZxdAWmf4jiiNtBu4C
571AgqRuKhimZU4/+yyimy0vSugqsdKNcPK+Bmb4NUSwlpsRj028Hy1qYk9wrjqXNu4dY6f4DRgI
pfUALh9oPOS86VcixtrG9M1H10vzLGPN1DvOH4p23HfzX9EjogQV2M1UTfTwBwp2zdzfNY0L0AWA
4DBmuew4nvGlPPmAFWKRb/KlqJdVwVMV2OczkwlI7eoASWqDIQGL70u/CouqlTJwRzPZyqlWbSLQ
CqqSaJUpRUzkb6J/eSH5qhVeB6irMMvB/emPTLLLEt+f9DBhKNQMKh9j7TV766CjH9PmRHO4QoD1
TqJWxeQStFAUefJAZGtCMIaIc1z5HcLLnRchNCxfNsyZvMbS7dJQ8M3vmgDIq1Cn6ZCQ6TXKbTPV
BjUqfnTbjXnxPmX4qaA/CpEiZOxpmhi7+ZXUiDPQASNzqyMWqU/Qe+srrZvUgiH4oFaGDrqjJ09N
dXM9zUtS3D2SmSsgge4xi1rkENekIHE+I2DNDfB2JnpD89hnvRL/uZd8CF9+eamRUzh+VNjoK7sO
X1esv3oA0bBx97QySBk9eXM7vdx+VrFFWeo7apkeZTBGgY5uHhiTuTX2/4CFItKO0kMFmj6bEkJT
PQczAwT2xSL6APQnv4KzTUyN7rM43ndqssfucWepgXZIeu7ocDT7CZjT/iPdlFPK8/WFQsR9vAlk
DjcNmVMgvDOoTex6xeUgRPh5clMnpsxGeXKAqRWnGQR7AliPg1TNpzYFTtHrTzrbRL8c6LPo+3H5
1NKW+l8ihWO+ISDfOYHfVRTttlK+HKCuvadR675UKPHlX3oZrhp8pMbqXHbHDopZsusozDXua+8c
jB8rLDvm5LbxaJnwUmLYRfFHvc2/pze+DcymWkommHXOqdU4dIAuPrwnAz2XP/ol1tQATumN/qMj
BPmPbh0hC4WW0mVKb5wOAnAQUpM3ZO7leLRpv+poH/wFJ0GFrlRrhcYpt1ZFKY04EgLZu/8f4aOA
gbxNLoJf4QEtf3vl33NhHfSQx4thzAw7GhnkWHRRu2/mgypKeDdU9jaMfahy+bYdeYtcR5qKP7on
L6owr9ycEWqCDOLcVtO8GuYJrNFd0wj9U5WbyFxqIZrnSeRIasKUoy9N4d/KLnRhaipqX1AWatQL
fWPOhvQ4lplqLBbwTJoPGETGBDPkEUHbOddC2mIj3aCXfhp0Wpdjh46vJbmdrauCmvYczUC2tKvZ
I1GsPuHuH05PisgvPDBvJ2N3WkkhP5xYRqFPO3k6XxEhBNRjTCBH2t+A3AOccjvtBFar+Co5fekj
ijOvkct4PwfKzMIrXEKWWH9vGb8XO8MOmzUcd4scF/muKNTQTh6+rPhNCyl2MYztCOY9Da3BRZMy
eMMcuO89XssYjaSNNgorLKhV88pwOq+QrDufuaNTVoMe2WtQabEIfnwfgdorSMIrWm1UGmKaR9IY
hFAMhqKnrif6/QHjetdXX5TUnQ93as9S7CPWFusZeEiKp5BmpOvLrbDDTHjI5YXWGHHZebmQyUP9
yOsw5a9ShPSsVDoaTtoKmVIOsrVnvc2ZOMGpRwaXUIcBg0el6YSq4L1UPAuygXAN+FqTtyfRccMq
jv59q8EraGveQUNyNL56hXkOvzU4VF9fxo96EjxsBxUZNKaoTzGS2nS5EUp+Dlxz9irWPJr558Ix
AUDLQzIl7RoA1w9NqzEcT0zo9LMWHASjSeZnr/htWuquT9G7rVw7+NUj3LNEBTeTk6duPbV8Ju/c
2devh0XE/GY8N1livAex4GNUdBPQ9LFprgO7muU6aD4k5HYYCpyqL5IR+PviRh25+lH1TpNa2f64
Rfe2MYhkmALHRFKM+9WAvkIDb6NsIb4y7W5P2X8wEImIZzkx607fFsboaDP11TW04tUrznR74EhC
wRSFtODmo/3seZGFMqKWS401hjnVRKADk4ikwAJdDGkHjmFfifmI6VO5Q0buPQ5ewlKmQKDnlrLx
CfaHY9B8LQUcd+y12DhxgCNQkBq5cgH/MNOy5u5iXuJ6si1Bx23j04EKFxDufQbzYHh4oQRMW8k/
p0hD2+MfwQ03FOnF/iTEZeHX3Q/Mzzfxq6e+d/wGBO/zBfkcntw1boWZSOYbXosEbQOTdhLUVVPV
ZrTYqudfHprddzFfVttRWC0uEq94ahbsA76YDQb3oTzkXIjL1qJOh47Zqrxxw3uKRxWjIZsB7YIg
3/sgEL1Fhzc9MvgwaM0wrsbpJe0yn4/K4kIACtmlD2xnZLthB9QUvucre7lR0h4YHY0agw3SMAai
9arJECs/kFhkFl23kVffF0cqsIIucAcQOkAX6nQq6Kzo2hRyUX63n7eKJhyLL4XmfsrViYo3BHTt
53Xx8D1wj+olLS+tJsCX6MVwoo3+nQ/taAusgEQlUtuGWvhSJVrivyoxXzIXbwI+ATttVFF0ukNp
pyIG6C7vXNGqAsn+Jd38w8Acx01tblPHF4MaXazSnoN2lzjvwaL8W0Hv3mcGUnzUqSnebdOOqN0d
iDiR9WpjeA8453Qd1JFlpcDi1tX/84Ww2b7978OhuhvtaXlvTPZQSClQeMMCINX4Yet5Hk8LcxiO
KLOcBMj9yArk1vgQMbr1vfmwJLtPChQl5r1TrjGjRDUCLor/4s3nD8JD9J30I00NauOqN9l/1V2k
JHGjUImtrI7xoJaU3Rg2aukepU/kT5rr2YIkbJwecCnGX9SiQ9EZOSJaT/h64ae9thhHrqlKCmnz
jMFQqr7KylmCnAs7M+pbjGoZLbYPLK5UvQ5zNX0btphvJDAwXcRi6Qo+WW/fw4N6wCxoKBBu8Pso
uEnZuEpCrfll99pRJmej5fA3LstCFZIOnMThAznJ+Zh9+HK9jI3rq6Yhq38632w2HM/YS9y7uB15
BFpFmeLMbMPNbHwaWfgC4rX99Za+uVrFJWHq23E3fydSamzeJsKZW1OLrIgb+RPGUlC6PjWUdn6a
L2UuMCfkDn/kp4ksOD6Pl3UXmpskgcmRpZLa6TclkikEjqDyPUbrumDv7rrUUjurCtcSvOr5zesv
sojvg74qM0yclTo/r7+ah1s0bm2V4unbuKItkWBJ9Dgsc4sY4iODU9464i3lWu7zYLNfl01VRHoq
S9CmdhvBPRvSNmLdHkgfxYpQ+FNbE8PUAAoiONKFQFWrEDuX+p10m5FVzdY8JstNVQiy0wEL8gUE
SjWPrz8VgDjr6TWC89YThNoLv8sPrGOBjwXK8NfukcZ+IANWwXecN2hfjhvKX7LI8p1abe6FkTN1
2IGtHsoO7GpyBvxCVeq3KYCTr6KAgBWJfq/dGZ1Pj9jT8r1LYMuOM/Vs9C/tgNgPEzZIJR1tlB1r
32piKvw+FZFP7x+n25x0hD2rko6ezCGhl1te7/oUg23Nn+V19++65auU7oWXG4B/XIJUqMAaUECR
Jp9xuCw+abWLlO+JyWC54WxTC/mK1I/IdIZTjCdt/1KjT7n6oopcr31DFJOBtGhhkgdYJ+2mhDVO
1HpNX4SOzs+wtrR8+ec9he5D4yyDtKJ1DHfvlRCBeSyEJh4eJkH4tUR4/c6zjQ+piMuLaN99EVML
le9wYv4fgRj+snVifOj1Wl02GJODhPe0BQzPh9M9y7GLFAaZ+baoDMCS6y41XOsmaSOaAkA0lCF1
4bL5K3EfJ5o5hYttMlIo3OBDQF6k3qWlxZkJVQQSwx+ZwDQSohw2Tw9K0xp2jrQ/yMJI1229pA/n
9b7dQ4eyjW+qIiW/yjHbuCCVJOHthkEb/7AprU5AxtDUARC2gHBpx1FH1uSqzkGLw75aGD79sBe5
XIcD7A/m4P9j5qxYJGmmyOKkX5iIbeYO1g+7qhTzZc/VANQ7R6MPPw3AsvowEFwsjiYSjjee/VZT
Dr/0TaiNBxujNnpAqGKSe+17BoKGsWJsDIGI6DWXRJ2tC2HSp1xWZQmkftfDnWVz7MBRJM6IpheW
llN5t8MZ2oLAf9w/ROrIKOOeHYO2y5jot5VNOsoAmOI9igdejGh8YuQruPFpaiM08hnTSFvTCyor
J5YzzS0jmwJXzpKIt8RZtazXDtp4KJ0++Bw4jXTRudxly6vL4kXWsaUWJT7h44GjXSTdkdnDjnGC
n9MR2+Qb8UvCQYFvOBcPGabgBUrxlYTSfmajMCFeuRXASJkAJLfaPeRQzkl4aSvONqwbwDq4EdjC
JryGQoZ+CFZtMY3tQgQLRMz03MSoLIW5e//FK2qxJ6owk0NXLiSoQgqF0qIrjFSRh83DPRL6IjNa
K7KvYdt1sv+9qp+PA/EyzEJX0qiWaPfkUiwHzCb2IpNAvP9Mwr5tkjU7s3Fg81GGxUnyotaJwrgl
s1kGNJubpRclNcLl4kdSc5zzQjYWIyQrd5zB1d3Q7ks+HijmjTqZOE0wSQ/rV9+3mD5xr+hzO4WD
49Dk/ryMhw0hEb9qq1gqDKLFQdJSVQyK3zJzwJl6Qso/2n8dDE5EnZbOO4Mo03Fv1XQxdVY7SWTb
zNTLDTgLN9CWdof/57KHGJGOhgB8xmVJxGNKzKrHkc+udILIpgcBkgQxl2L/tmGaDb10EC53oSn6
bQw2GNv9leCwoIsSoqZdrrvErNmDR7mDdizNNDgdnJWtUJMt9wcWAA4dBqgvtNd++RXJ6hFi+Gcn
sn6ls+FjBo1RKflzO0J+v3k7b3MsCPuIy49FxL7zcjwc+5fNlcUN9MxHAWevUXOR+d9EupVtsh/A
CsJtg8URexrcbkpXorWpUU8QtG0Ctxl34Gc093sv1PMyE5NmgPd9oZ90dkIIDDtCfy4obUJnD0QK
3pkhnxV3TFN2aOAWBH4rysKhtyCjdBgm5JEMaUHfP208G+ONMiKGuOEsGAezI9W3/ymt4Nhivi2d
u9Cp9zGd+++u8jQF957m4tBwm23rEh38iTtF//jaxDJQbDIwB7LnTXLbYYAqKb0DDRuWvHqa6Cgg
DOaxa18KizaNzX1m7FYAKLXXZeuNbt6MoZd0Ll6qqK5R+twZsUMAftuG6PCEH/9uD+Vr/gAF4Mk0
ptzx22Z/Shh09j/9uo55FKuARamNvX1E//otMdlJ/j1v91umOz0Ip65EkuGLkes6zNqVi6PfjCUa
T045uVd/LVJGmoVVM9eWiSOa/B8ooZvWZVRzIUQDagfeqOAuwebOnAY0y3q9XPp51amJ3XnLEUlA
PaqoMBLc/uHXOFBNG/J37blqYscak05YzFUCu+ekKG2cGas/4AhyGyu0+7hxS8qsOoBDdu3fA1rf
Em6BVVD20gskJTitkv4DrEk/cNGVLaA8eOlKeCsc0dLY0JcKRFGstaX1O/AIHH5qriQFub14k6qh
acA1q0K8nXeumQZYaNC9wmdaKE+x+Rm3ORZfBySB6Jdd5M7aE3C5W9lr7QxTj9uDl2xd5hgdLJrg
RevmrdxvprUlW1uegPkd2NCLwpCuP8DTyX1zPcftCcoQCZ8b7nPxeg6cPUhQTQilTGWucv2eLkJG
l2g1JG7i5I+1UgZj2E+MeRdvpwQhc33jmpZn7TUrcTpMvR5uEdgxkTj3teM+8dYAmcM6QP2Gqg3r
Fv0zjg7QqGyhPjMfxOhEG9SYzPnDuqHhEvkJbRUwEMBN5FuTYFTF7DR7oIBA12ocNGZpXHodVKzw
B/Q1bsV3JUt8L2oWtepbJWXZLVtxVPTyTiwgSXMYPkXdoMgRIj0VZuulzY7dwyOiUxq/YwGetQQ0
OT4QL401pZXkg63SNxsVPrZEj/ElO/g75TkmuqpK8UwSIiSoP8gcxZoWFWzmAOF6aRs4iZXy9Tti
QaGmVVlO6P6wd/ROBMrDuIQDBGrUxda3+GH4KlTxDDquuCfvcSeWm5DnCuYOpiRcsdMd51wqNzey
q2vaiUuvYvTJKUvqY202fOCn0N8tjps+vyfwvQXNZR2fkDF04BsZAfJeyxyiMS8XA6h35MnaDnYt
vJ7VKpiS6kE5xLd8eGaVOK1TgyZg9YmvzjhcfkjDZQGhQ+biotvInG0fngNOGPtm04RFfEfD0yuq
J3sPTSgNhwJNlcNoaTK9sM3ommirYNvwvHu3qYyx0qb9Ecms/kjyHW6kwkr0i5JJcR+4XsjTAiFI
ASqfQyHjYvbe4tROhL746WjTaKJAyE+Kq7Zq4Iix2+aIjRMf6lbaN4/ZqjsV0o/p0ItXtsBdUixN
DFfLcQdjpnN4wT1zyvdq5Oolh7HIVEgsjcwtcI6w4pUoolT1vmmphgeE7WyZm1uOYy6B0vIQlBoF
Wl9CN0JvDkakOodHFx0VVkX1FYvdxr1eUcvwWmsRrkazi+6+r1iN15CDNRCMpSB5bjE3+8ghEfCk
bivPOSx06xDfNz8byzNFU83nLW3blFZn3qstsgNmhdxDG8jhtxtEMMZeEu51hFBsf/meLqJZQ87P
kq+i9OkDIEuKwQawLeFlb5MXJYVrmXvQo3+xndWxR3w8quZnDoJMrQGYyoW1llNR0efFH5KDQp/Z
KRAzTZv97L8L/NKSKjq0sHVMb5KtCEVCkIi7VlPitJ7w6SuOfqSLVQku99CT1XA51gRoAk5hLvFu
m0ZwAZ1sBVwpxukeNTNHSKHs6tz9JTIYScxwTjtBg7H5YeHH9cFUGgZGIi/H+kBSA2cMyagtdnna
IyZa6aHprgOfg7JX5Hy5wSJkTMhCOj1mOa16XZwSSSuOAOFVzRc53P71+jgSI8MtfBG23ivSY3Y2
5BalLb+FlMMNsEivge9NiHj68zmiPEMMD6E+I5xYs65Lol+V+pgDbKxMQLPw9dvRWnkmjSCEdIMy
6I7N2aP8NnCtKPUGCxHnLPDNI920xnCrrv3l5yQ7nrXEKyy9CmYYPckMYJho1dCwwR3wVjw4Q4i6
YmwljD+I8wQ4ZBYfKtdxxwJq4Kb32P54jaQ0eboIWdKfUlyJZoTtFSiI2HUb6pScWvqs4iw/6YFC
5afGbT+cfhuBfaR8lJUs6uaX8jzG2S2ZDiDJQhGxVieVn6FOjLWA7CTNlFZkPESK2zMDewNUZdPa
FaRYSmhLXyKF5V5G++r6LaDqAqgKJGhP2O2Lf5HWDCQkLHzPD/+wj/oU6ivGF0y0Bx1M/vOWCZCC
oc4ytgimybNBNv+JqJrq83GetVIkvc8LxQ6h26lMvbMm8HoZm8I7mr1W4loqNslIv8lRf2IcAzWJ
By1mAxEpBKh5wOboWNz7EEpLUwJFTYTPytJRA+DfWXESz73svHPE1t1yZEkazrpQKRrJnVxlKyC2
r2/bDWs+5C5M/60TLGcbw1mtpFCsXh8+++rlwUhFNOmUPOcE5p7uv1tJV7+6MG6X0iWxZy0Mw9Py
Z2SJBo33oOa0ZPweYuIQY1X3/U0EDmMXueqWyamWiw95gQ4txT7P9Si6tEYk/bJmb/lYKvmzpANh
6y1Hk5IghsHvr6lzWKA8uneYl/+TGkhlkh0Gjk26l49/oKcHqMCWB5Xv7dohpu4RX2U6DeW5CC64
PUG4jLtoct8jpok3JqfIblgQ5iG2nrAt5R30+7vToujHHk8PwhKJ52ONXrpw0sq/wHU0gKMT+73O
R8sTbQlxQeQJvCbvq3tyBOgRNfRK4X9P25ITS2dAYykGpKk9Me4Qj+nxy4tcJX0x/tf8ge/z3jXv
ZAACihexK7ETfj2fHJNoE5iRJsUggc3j7x/tDhi/FOHRuxh1SGyvf32A7RDBqxU9YoO2WmKYoNzh
K9TE5IcwTFQqAMWtshNEwqnXhomgMYrJT7SxaMD6p7lhDERycNPv9CMWs4jSIo4rvUUtQ8Q+LuB0
c/fWVgdcdMFeA5s3YUrvRKiNNGIS+V0kntrR8XpM4/Z3nKVEZp6/KOoxma8kECR+/Vct26Hiu4Zb
j6Fqv0mVBZekEuEcymNodSz59YnLDvcG5jSxeQWcW74D9i0Psk9+RE3TZN1YuZ1Z968kg+hd/Mu9
4JXBvtMEvOd4Ly6/jkzTgdFhj29rk3sXh+m1gCHaPOxU6rBQwmgJVnECxDOCIOR89AfeCW+7C9gE
1ENm1eBYgA1XX30fpMBu4yIDVBPcWDG8J2Z3fKOWCTM1PaQhiTsn2oaZlFgg3XiViZRcXW2YbXrs
vXw9MqSwWywwKZVRKwSc1xGColiFDcRTRj15eFMZ4BK7Kvo13+bhvOr0ogH/7fSOyaDpdFMzv5Y+
KVCSdtKpahA/fxMYXeImBiTB3JkGhoOluaLC+fRwUIdfSup98YgYY8HrlJDYAesm1ZMk51Q4/JkR
If6kAUa7F/bP+EUk+k/jZSG7RcA94M3a3t7UgozgW1hPm9dPNwGw1oYpSGy96K+hyiG2S7N3KWbi
T1RG1f8QreqIQwZhuNZywo5NwLlLWHNemFqFbbgI68eYnYFXQvWSJRu73eO40Pkys2gf2h5vGhvD
1Y6CUzYzLWihPEMh5vtmgwfky42bUrWgL0JJAcKDcw3QVEeTgCmtBqBJ4ITMlRvv7I+tFWRtpTKV
DtF9lQzhdh7cb71jgV5/qSAqQMhcMAW3Zjf918StI2FFFVexyfqtLCjzjirBbFip1EBUIXG/yZBe
pRbaNXNPUCeXjRcDFIJ31oOa7wLn/pBecqeOoY6DJZ6V/YvRqzpfaJY8vtuGJ2+dU/EcOmux0eD6
n20VMqp2wkIvFgCTc4LrMwYadyFylM0jpfYB8Eq3+bFizB2geFw56jl9GQ0Z4uVk7V4iU3M/yBHH
Eor6YLGpJ3cIKYZXiNqrIsS88vv4BGf4TSodXVndLY3RwTwzzcwADXLC41OPJLE6K+sy0nfH4xyn
GFO+SldbUsjlw40qmOmTYB6pE6lDRUkVPi/KfIYhYgRMM/IXFg1eUpg/R1hGVR2NgEp9fQ9Y2V+2
U6h6akeUqzdZAXIEriadGO2VQZLDQaZMBJx1rEBxHLfil4v5ec00I52I73fX2wkEO+b0NHRRZxDL
EpiWryoVqgiBc/x3fxKzLfzoVzw4264ZKJgOh/bzyWdECf+4r3A0qcI7OVSDd7c4CzDyUo9ZlDta
JwD/sKsSmg80e+PQL/PWsINFzfJdBOdmjL3z4QjzBxjJv173Ovme+gT/rbYgFPajZhTzqmjPeWo+
hV40JY8Ly5LMpJebb3ijofj1u3FRsqUEPELT1xXR6puGcik+hAM4OcFG6Jwxe7oCbZhdZckwaCYp
2AWQztn/ObgFqJYxLApwBYxtLqkKbOAjAId4k26+hTi+r1jFzsxQsph7T7w2KSDdYLw338nbnmfV
7hxHwcNSfockzQdQQzgghRrLGeU6x/Q8JUraeKlA5GrCw/8gMwJVQpWHmimL/4zVDuUikiywhhfG
W+amrJ6ptDA7IUr3clJFDG1+NmIfAvTj+qUGKzoRaocXDE9yMb/PRguRIWo+zVea6HdRiH6BSmX7
YNUxUBryS+WbgmZ0Gwk63BFZ0iU8wCHzoHv5QKjiqmRKfYmQvLS4slBqhfj7vWlbuChKPv/mdNE7
Sq6IUBIZ6CswppMBNrMDrYfVm21r0MMf6rYYJcDIQoW0AYV9r66456fDAr8xghMqO5gtrpRRx1DO
wrNQ2R0166zJ/a2+lzBv28pzpeRygbDPCiHhNSoyfA7HsoOh6rlx3eDLkO5stGN5xgnYabeiX/Dh
bCdULamq9ITIZXBdq0Xu6I1YSaeuxiTI6aPUKPLZZvfFjytMV9sKOWzYT9ZlCKK1URa0fWYqDg+a
cskVBMSFzdrEy+ZYjFLs0UWOcaX0pHpmzUh38YUMKToH4czbFJ0QiEJBnlagGgloFWa8qgc7AEel
67yfOLJog7oMr27jmydyUWzoNVrFvDq42e5qpTSwjg6ri+xe2ijJ+glcv7sTBe8k5pPM87mEqoCA
1PnARSo4QAq9CGTG1KT53Bt383zcnuOznO904JEs9WlVwC7NQy2xkyP7/zhrr3uV+ZDe/wB+RAcX
ydAYEU7DsMLjVMr/lq/iZcdXDf9q9NVirzmc1FOPR76p0v/B0Z3bS8J6BNCPdkBL/2lFE9/cz9oc
qB3z8jvLnqI2Wndy0wXhWtJCBYRXR+Z60ta4SMepTOLXSJSKfI2ZynbZcUEnXDcbZ34gX5tAB++h
QNE5jMsSKtj82Sh7Qgd8xuBhzQPPz4I6LHF+cpacAPLxBF3Z4cuRQK6q6FSS1aX6oryfL7fRl7I6
OTBN9lmHMPG2t+N8EXtNf5bZ10wfZXEK9HWco53qLVcPfzj7ZSaHeZU0J3OGi09S7HULU138gY4A
0kgvNArB1FOySjrR3V0XuMNIttplfTW+FIDB1fF2MaIoWbz0PHV07zT2IoxwLD9TlhEV2TSUCjCH
BfeGMEg3SmlaFlpqnK+ah30ttY78THtCDxCKzLWxLGPh/wm6UsfiOEfk3u0o+jQkvk/sDxRJULof
NBGNbhKgvJM+fH+B7M6fR6mCuxCy6HSFJdrT96WH3pzqv7gxUDy0AoE/2LELwsdcwJ1YxenkvVhO
+ClGRQudTgPN8zRydbmHms0D1M34p9ioCZbP91VWDZzV2ZYIYtuFBqJbLRw20ignHqyuTSiCu9oq
fcoBepFvChyrm4jfFylA2kb/92dqOe+kzfY76OX42VaUwjsQjrnI4EAX+UhOOnYc6PrdBn2DfngX
HwUQN8FoUYPC/oFwHFJEU8GRtalCuKKhDqUcyzpFwiQwRpYKzQh7lKQzqWjP5Gaoz8dvTUZYgPgN
RwzX/UD+jJyznSdhavVeB5Gu98b28eURLiAo9Ns7dB/XIzfHHP/G0rimb5nZtCiM+2BQts3Nz1vt
IByJpIkhiSbImB48WMW/lB3D8IW9PX+wjyFBhPqBNdvLMHA4donfBBj7GVRCNZsFF8psdQSfw310
BG2dAfxqjbLHYFIGGtjn50jXqyc1EufwKbWrlrXD3axTxZbEBZ7u+2ivzgkiYBH3E16tnmVmNCpa
oCUbeCm+lYOuSJ28plNtnFWzXylM2Y0FjTfW7WojTZMYVOF0lVyuy6DQ9mITr4ReGQ/yaNCQ3Jvi
6hT6JAzLhKVVzcNwu/aSc1hwNsJfmcWc5IkePPm2uSQ0XQiErwTx6R8lrZAbjBmYDE71iHVaAn1y
W82W2gzcRZvkUmXLgA8uTHa2ts4bjH+b08mrtmHsfBYQog+sJkicVQLW63Ch8GLVf/bNvsCbeImJ
QFbJT0m8KU2WIuM7NHrxQ1IL95RRjAIBAXsxTfM7w4P6lj3PFswBfFhoeBY/WPiGVu/4crwblj3r
sea9UvwaBZf9mnTQOO9J/ayizSBbxuoG8Dn+mtHzAue6HmViR7/1D+0vCXcx+8P2p5NojgyKJgcy
6JSdJdcBAASUux6AvcfeoXn42tjU8uhmzpMBygjYKJArkCHa9Z4GP0w6a0rtsVNDj08PqJwkZABM
enUz09i/dCB8qT446bbpsCHIjke1Jrvg2DWsDb6tHHyedm/1+7nb9wSgjhhqNo2j1KGdBr1+C5F2
TZU9jQX6T2dPjHnfuLrmZjZjNFuYe8xcfUGF01NICOrgl8KuxxyHwlZA7fBKsQ8lt6JDHKh/b0Vq
+3c8SbwK+37RRq3vNrPJbmqjyvufayAJDHaMshqiaYhwhwW/Yk9ShtUyuTR8MQqWK2i3oOVe0YOi
Us2KFOow/QbuURjcFbx9bY4Ymphdh1y6+4oFsHiu+S599ovRkKaJisiDC5j6QMhMxmAVgFGzeX0w
z1EBNBumyoiCTWhzdNbRs0l37sTi7DpK2nYAUbFkPnp8EveQha2cDns2L1zwHQbbafYJukrLPcz0
+H9AOdr7c1ngCpbGSPYwPvBkRz2cMXfORQ4SVj3ylNR+NI21FDzrxsnV2KHH6cOibdtOEUBiq/Bz
EWRh0mVDzXgiX0VEZHqCi85uhrEz12QOWdonuTpVT453QX2WakCUJwMt5zeRq8+AuS3zDrrr2MTD
eiQqZjPeFJLGwuuEqxDQly1VfW//IzhPiSRvvPDOEdSyLeMeYHC1rMWtWp5m8aAVpSCRvrTI87Kb
WP5JHPDG4fEk2i63VmWME/t85tgQrHw3I4zLC3xhu4gYAxIIi58TsW/LLIrtDAxufvtGqT/aOKDs
i23kNTssn8IZ/VXKUQVKKUOhzFllNLP6LlNjRf51bPpPkdrMFDZRRUdXLJyDOzIP/HNs8onObSna
RgdrgIRQCYlG9a8HnJ+Tw9HHrLQYPs97mxqTtjh3cbl9ZNlZS8sbtifVusGjvwQmEQNqH91e/BFF
VZSnXBQF8Xf+4SCNuk4nVccGAHGQDSUcJLjFzni6/qU9pIkIOTA72/8zhLyKdxiuwXdsAc8sG5c+
um2YLVdKMQ7BvhpkhNGWQ90VKMSgYgs3rU+fIGGpiSwZoNlgTXCjrMU5LDnRIi72p9tgl56KVhef
mMSj1vAK3c6oHXc54aIcwYN+4o+R8hcbbAapB6Ai0o4ZraeuJ2kVVl+Wb+YBUGIyhuczihlHWfGL
8Ttt2w9c7Kt3D8P0y9+gups/ybGGVCav6GYqVFvQkUBQfVicIml0vvBRR1tqUxj9yfSJb6Fejg/I
6YOcHMYviE1pBsHEHv32+BILPO+T8Jf9T7a80sjqy5dWD8sV4ie46NiwvEQl+L5ZMQvccBZ05IZe
7vgHVx6CtLw9IYfee/JDY0DPvOuPXgvfgqg6B1aS6zuScm48Z+cmamCCHv3qqGqKyFYdNv1W1aAW
fSTpyG1L8AopwIM+ERbyDrVdG4Hj8c81oo4jLvdtbvNKWIdaW0BUZsx0L4R+dV0lY3NKfl11eoJL
vVv7n8c3mkwthMUiyG1fWeJcjh/Ad3PqzlANBUDTNXru6tVtomdonUTOhlJS9nwCu7UENGUiufmg
yJUFFFG7AZax5D057jI4gV6YpZJHXLT+CHyq0zb9gDa9XtTiEscZ1x1H8oe7TFux1saw/wN82VCY
Hh8+08i9JqPLJnLwH+Trjk+J9hbSRCpgOXwEbYIa46I5LjUKsd7HYmWsXSYCru+kmNwskbihS5sH
leJ+IRiSUEQ4kj9Kl1M2sp3hAFuBnNlcPlQKsZwg0Gt8Fwbnqy9wznIeWKtBluXz+T0dVCDHU4fo
EY/QsS0BY2PfUPG5dDGMAD1H8qUQaulXUXsPb5ERQ/pLmM5WJWmms3CgQ8YkDq0eRzQ3qFLHh4io
+zVzVmkvNvIkpkF/omIqPQO2KQCJzH3iaBms15NTEuL4fklHQC21zvgiaFE/K6DvYMBkog+MTJ7O
S4tQ9c8eBku5iXWyAJsXlLCKcdOTaHaRlWu5oB5SaZvubtlGscYtOLHR2IPWZuuNOGd/6gXeMiGQ
D99oh5DDUZ2sQm5IWLtj2FEhsduzjBoufSNQOmKu7imdFz4QLD1zoMOPZfrRvkGhfKWRNyr8yic+
rZRdv5NX2d73jQ/oTco05S2cHzpTagNV43QLtgo302M7nOB22a2LXyYDZ1mcruhcSRVpHBfzDr86
wXj311DeEaHDJ9pIKZh9xwIT/6r16js4Sc2DFiRwkxxm+0kihTYzZaO2alThC0B1jQ4JtwYUjkjp
yNtXWC/j2BWUVckGU5sv80Wqd8lfix+cewiiCjwCkSX/mFzHDKKa4XXsfZzKPjwGbyMrLFa9bxPE
xpS6+YQ9Se8QKmU4x3iQqX3+qnHsdxgot7Rhug1T75W3TTXAXNKewGlXoBKZim9prdHLYARoCuhI
i1vCTBOApnXCYK8VAkgtIn47M4gc6CrfduoADnG9VfQFAn8uOTu6IWyAvjEtsKUaVz/OtTyNnx+7
XCY6Bo+V0diUy/pFV42AlCinAgT1G8ectm+Ly+hF/rHBoEZvhHOg7EjnIgQf6kroY0Na4sdk4ALi
eTyvMLQxC8zb1MmsXlLFfLUqZZRYKJpGiv8aS8RYY5jfKnnCTcniJUKLTPV5LLJCVLgUAxEndEU5
byV1XRJe9NabG+zZblurbSWp6SzvLQTJFM/UMaooSuQY3PZXdVHQBAKmHNIz1FU5AnjJ9BYQLOO5
Fofszbih4uGn/S+ewuBMAmnQ+bqXhS5q1TCIF99xqLpJmXwQspzFLhOD64v+iKS91UOnLXInKxHG
Ppqdzz5f8cP2Aei7knLvyprNplm6sxY6AYIOr10jOAzk4yLbejZ7lduhke+1gWq2m58e81LA55i9
q9d9lqyoOC3w1SE4EvCxBC+XW0K2jTvIIrfNhojrb3AazI2lOOxjMDTOKTaLX66WBTyst2S0RS+8
LcZu8cw8ELyGN9QqJtZahcywVSC98Fxm/XZBWloJT6XFiKFEAjxfj264Kv5OjGJkI/LtrMEdGyNN
072mr4zSsltqETLpYQWtD3pXqMaEi+LA/RD4m4z9/p4qdnrBL2iuFHP8RCWYyzNjJGVArxJ1fKbg
5UyLzzbri8C+v+XYe5xzKzC6t2XAw8zbby9i6g7pvp66JIcD0jpVrButVeVXcEGOY9pKZmQHTgRz
1TR/EMDoiQT/bFyyt9q4nXWJb0k91lCzN9EsdwWkNfUymxal/h2XDQ1YOupYv5PxzLQWeBqt4IUq
yZkcvQFOi+xprDOLa1w+NTj4WEEXjTo5805GoVKkct2ehfzZHg8vs5xXny753SQkdBoniMXJGF4p
TXIhTxlguZYnorxJ+U3SMrNyrCRWl2TlNRZTw4sr9ePlIvfSoFeuc91Jf2gWPSgJdVVf8Zn9wZ40
/6P0ZpWoowCJNb+n/1tOreH/drvf/Cjn2Z4StJGmc43TNuygU9t7ilJgnY9SO2UcCeJ/l0hPyJrI
gBXPNnpLZMdKHbf1h9KuYF2iYqV0+lpqdogJIeobh80LyEZaarDPkL2HrnqByOCIDmuMxcz7XNY1
JEcktZQYF5KYu60OxDhVqRMNSU08+cnPcvK/vkAk8fN2e5cUtKFxJFGqH6mkKSV1WHuAz+RVoSVl
iEyIvnqnvQRhiIvq5XxfrHeb9k4yCMdAWHPnZtGUUqNtcgU8Ia7XJvVlYBS+fIlb2NAFPYF1EnmP
3lLsy/Zqp31DEyw2PZfH0p4HYMJ7SMf07hOT4ebX9IzQGQE0WvgOx2yBaJBrP0e99qmajnIDesdh
tn4lXFOr9TqCMMHNo9Bfwy36A2aQ4g9cGCEaLAAGc7ybwFQH39LmGxMYvavAxz/iA0LQENqmKHzH
mpqvtAlqommDty9XM/e7o86Uc/Ewt1ggkYGf3NBZ3PVBajSk+JVdKfHChGxvlGwWojHuQ/J7w1t0
TuIDwNbu2eyX8o/v/D/Nv2MoEWu0TpzBpYMsPoZmUiviyAcp/C3yGqCsYrovmkXcBmcB7B9VwNZu
aMiZ2a5mQ614rmGKx3kM0uqWl2+bdDnJCfxbxtQF0bqrKLdYMZZLgDen57vVDkF//KPDRekvHF1U
QD7zNZjPKu6C8tBwJz8p8HB4Ux/XAXRrmbR7AS5poJk7njDmN5OBrsn+GKJEBDErQRFDksA5vvdw
qD6pso36f8EQGrbsrlgDs0jrM2u2YSOG6SGIB9amhKq8hoOsfDg6li3dFRV5gesBAjXl7N1qjqOi
QEJkcINCRo9EurA7qzlx7ZJ11o3LecYRnNtKh4UOS06vfeQ2LlYoukLE/cOOEgrdVHRU+lvfF4Xu
z958PD06cJN8exmXLSNC/RQCj6DIGUC+enBmHT95pdV9UPlY1+UNNJhCsiZxR2vD+Lx+ED+8Pwe9
ODcO7bi03i4SVi/M4UvF3Z687RBV31T6WYrxaKAYbrD8apOtD3g0b0NH3EQJ3Q6lDPpLI2BtaSLs
Az5Zl4vSJ2FONRqvyTwkdv0DYaMSqGYEOaFkFPbtymX0d7T0s6i8uGGs7DzAiybpmLKZELJpwPyj
h56JJyuiLPlRcXvrhoTBOXH7mN/tzhoutR2xBwIBAio3tSZAjNhikhwSapI8YhHDf0XHT56KPKxz
WSfzQ5+IAAIzyFAIFuY3SM+AZvT5PJi3aDRqizpLztl0UI2t+KxZPICZLQIolBs8daNYUdeLa2Fw
+TLctVdxKYJqplX012YJkMdBKyBLe063e036WPGGnvU2CJ1n/4I6FdrLhVVbS05MdGWVzmk48tPy
TAwKMjK4cQ4nUmSsTm1F/z4iFCa6/Ncw5qjJkKrGvLRktlB8y8aPAyi76yYvGYwDDHCIZHo4dhYT
wEFFBuCZP/SI7St9Og+k8Li/Yih651kpRxPzmzCRs0L4m8FCx4j+pDv4/2gMInWw0sBp6b9TJwOR
85EYGnGIuWyqDw0FfOk3c1CznDFQwSzDoYaAXM7KPMYhxndeoSeGUX+KfaDxs8jNc2DRaZO+AJ0b
d//7PSwL14JbUZieppxt+k13NnG5J1lSPd+Lw9LDGIyQIVkksnSZuAPIChsZFNsTVSTVDgjbuP1y
OqsbKgwqDFBWXkOY+par22VebqkT8Lb3+V6TBQ8jmZli51/omOD5nMsx45W/pvG73mN/jiqmApt9
hFyfFJRCjnfWaZ6OkERLdOTAHVk9cAGzdOnP2zlpHKNCyWNlWIYskYBHP7gp2tg3OS36pmhBu2j6
RM9tEIyGY0oW6ijvb9THweK0CbEf3mYU8/u0NWmMKrTvnEoAazeO8J0fRwMq8pzgrGIaqerkIOPQ
91eQHkd11SiUDxQlGIlcvXopHxhBIKvg5m4ZDvmCKqjvPfLm1aayVcY4LY02BIpkMFimGmNBtHY9
UAMIPnrU+ofac6EkdpkSmepDrUoiUyVWqKjzmxQX8O6Tq6WUEpCtb/uzai/1S7sTVTaOL2crdLvW
CqDzj4MWPI9FgFz5txR4AbbYuZjlCldPMLQG4TTfnxgWc7pYinwqsB9N8eyun1FRiAGwrrfHB8ST
Ar8onJs3uW7wKAbOzNpES0eiJgRPk8pLdpQ1QO2BUXUaSf5RT+7vLQ+CjU1Vhy1+GzAKFXSOtx/H
slUsZOYlInEkGHmSUa72u4aeWQ2+WIN8Apku8LRN2RmlS47V8ARjEEJcF9sFS5wIZuirGiMHmTVb
Vd4VQ7b1RmiDseea7ARt6Pxp6pXfVg3hl4qZBnjyCSccd3gnDsRVuL0j5sLXgvF/eBTcGPnjAA4S
HiZaSkuubkekJ7VG7E1ufEyMBYV6VvDkUr1bKaz2bI719r4Iiju49FejoA77zM0Ad76/eNP8q45S
Ihy1q56QTM4oS8nsIKbQZg0EEfx0ezxXfL8LCS4VTsIRoIfTRQHjbINyOOAFcg2pcfVku0ny0hVy
ZDtsFLWxeBTd+HdSWTL6znqbRxhhL4PUxVyNT8lOvLcKZBHxMHdJrySdKSjldqQ9AoZqJng06lWF
NUIXn45+t75HlFjJcDkowtqBAiEt9jK0lJUaXpLuWvBpVA1SfOtS+UnBdalI1GxkBjG2Gbza/IzQ
UZRRz9QJ4VWheL/EQYNKoek+dXNZ+1CtLTQu8RS9jiQ8NX6uogtlwW8j5uT5kq4ZnMmq3eyp278c
qQsiaEdclswhf+NwyCxc7p8JlI4zrW/nIZqBQc7t3xh5XGYEVn/v45feAUkAAME60rxYZMn0flae
yVL+4PPDIzvjbJX1ExucpeQmo2x5m/hqSsNmOxY8nVm1QaSQ6X0rewaQtPosXWRa2Fb51gSIUm4S
2BLiu7e1MLwSWy1tr7gRKjPsIO0YKb5ZW/F5OLQUqyGNpilvI2foHInv6c1lLQbCl0/BdEApT6V8
e05hy7q56eRtavZhBhFZZi7+vx1mXd1nn4pMppUUo5g00l0MMbNCayddU8xNGBCsQW2DqNiEu1YV
CCL8bZbmVNsZlYKccvLx+auvcFwAtgR3/QqyLhogOJVbW3adYLBZNLsdSxaif6J3h3wP5Ng7T2Hr
Zo1T9AnxQ/SEwO4I3Lcfl8PBuSFX+ExBRL1IIkTLIoooC+08kknHbDyFxebaM73tq0IeSLZCEL8u
hhxeWPY/l4DLz9IyN9z28ZMVRmjNRpK3AiCuWr17cVJvoV37KQhqTJCXrwpz49uR6mFbo4xDNhUC
JNjc2ZJzfut89RuvlepdXHHrPCEQqZ5YzwUKCDvf7GoFrpba1mvuzMvlxfv3qjq+HNU/XrCJAAv0
M7+xbEKNRAyzR8kxj0vK9REejA3UsP1qzmyXCbruIrVFWvg0bLZs0l6lFt91uE8Tqixr3L7+Erbj
e7FLTr9mLqSA1Bijgd+ZDQWy6Bh18aJCmSpKXNXhaJr/swyNzv8NR9XINarHUhgt/Lqd+TNuveJC
qOUKqKO6mMVDk5RW01+MmKEN+FV0djUw/maq2ijuw0SpmB08qHy/ey7miEAAtuCSrqKDsvVHyfWL
DXC3aMr6TSZBxmjMpOIl9rreOcTmiFTJgCQrbyZIGe98JSwvQ3ZMfDceeuq1qz2o58G6WwJZqigY
EYL1GUQK2i0T/xd837PFwVLsm3QRVkaGe07tWPPv6jAAknACs5QwGo615R2LQzKC+PnDZgiH193c
QlspnHmNSuwHXJ+bzJul527wx60Q7ymXSb/Jk7VVQ32abrf++HppvD1ckSts3RmND92U05ceSZu3
jyGtjNXu3LLNl0W824DmX2EWGOatMK0YeabBGXm6r2ecJpd6Mdj3prk1UvxTSBFVaUETjvEmKH1V
NweYPmT/ZAexIa24n9K/x7Y+72aeCXsbWZT4L7tsCxdd/Jbd0FYl4/n1Qb5Yh5c/nfSVbyrneQKO
gkZx8VJ91eg+gVhm5Dfxk9k8n5ceIrmyG4XStiJRIEyOssheZF176L7kUn3pWg6vijzpz9Uzn786
TfUocLUGfTtuJ8e7NXyLqz+8OuoKYC21ohcJQmqaGOnMf4dTjV1mZXFIO08SObm/kJ7IGu5tCCRZ
aWjNFgr56gir9d1C6IOzkUCoRq7gKQIR6I5+/lVLMbFrQHzWdE3pocoIpG4HMuynlQvm+zV1bKsl
ymoBXwB+t307OD7yCqlTs4lbMgTGy1NHm3hYT1QACUhp9i/Nk2K24J/cRqt76v9fuu/ILAlzT7NI
VWwjSASU/TpHCt96jUWvR98h3fpe3Q7mczf+vqKXZY3ia9BEpXBo952nCuejUPqSQZUehS4jHLT8
YNktHhL4PlNFM9ZxqImWnR5MPSOAZS349Hmb+UByD9QcLODHLu8Bwrb7IUydKGEqlbtKSg81xsOT
/OuFMQdtUD3CudPUF4tvCueW/Mv3L/W4Ne9txt1l7ma4u0e/ic7aOh2WooxwI4kvNKQz+df9RmQS
DcMNe3qHFvQ1slarwzHNHqA18aIBWuyvr8+gsgrXU9ez7PEBKd9tKhY7krxWSyGJUUfmv7J4EYrS
srYF4R8oeJ2EaF9QEq7tf7i82LJB2v8W2dCVK3273ZH/HgH81kMLZguUYhkV7Gaq93xXLMnwFhRu
6jNYBXTMESDN+nvZa+XwVRPyJl0nOvm71r++pLKbDv+lUAuuesG4J9Q4BNMqKu5ZuPI2xkEGV3Uv
XazEPYIr2SR4tIf1chdFkf777SK6ZrzHASaJ8B6YfYj16eHtbgkNBj/a+uXi1yS90BQceNmKwbLo
xV6WULGPZyZbBa5zd18YDS6l3+84srO7QFr5xuT5AZMp3joNx291ZT146pXQlmNY3CexgU/LznIW
x+jKdeXSHJO5dxh25f7+6iDKZyt+qoh6R3fiMtgWJncIqqJr2PSniCkbzCrJneExJYIUmVbheOA7
Odu+BwRiDki2EnWn4OEfr7oahD/eHmHSMVsEX1/u27JKqvosWO4IC9FSfwhIoiLgnm9nQV2CmhBZ
pd3KJ+ID8oR/5XDkaGhEwWZe5h727BUph2dwOBbHGPRtGyPlzV6TiVHnx4G/EntbDShnx0DAYJ7D
Ghd+cv9WvcbBwXx0Zq7qSC6jh7FVAjklwVuGgpoLWnEXg1BoMNAe1jLP5NSi4Z/8kev1Bl/HiaJe
d7bD3upXMJtY6OWu29FGRYnpfb5EjuIMnwoFiZ7ZPdyhqcGC24HyWMUbt1PyBNWpNafNBXX0xSMp
q/HtgIUSifKxWLdkKrRIQXhLaVGCTiA/6TivmJPR3Q+SKQRQdTnj0v/F8yReHa9ud7QqLnNjhtiY
KtIK2+o1dezSVYrOiYtIt+kN/8bKuvSCAFs+naRU+HHAv08PvALm91TLlZ55c4t9sQBo6LsvQNLi
AVgVr4x45tgxwurX8nT0bjUCIxrCTeQlrkCKrqpe4q60Qj9xlHp+40zQnNDbjkkgR+ezUlp3oPDC
KuwXeUPUH0IocG27fPzEptCP2nE7m9lew2g/jHDEWbxRff/xa/V2YryRxZa2yD02wgk3D3q4TJFX
c3GiyP18lqN9K0Jd5z7e8F76VJAb222wRF5vFfpzKGKorTkpEJCNOdh838t5LTM06W3Wx8zbRRlV
bh6bHFzf8K3K8LvG9ykeZ5WESt56R4A/4vXoHWLE8LwCEYvgeBVszv8N0EAGFCgp2l0Pwn3ki+G6
CAnqzTHDM4egy/o0WR5gPhf08HCOlC/i9ECUlfoVrm9+ra+MxHwYDP6NNyHSfIsbEq+iKqaCyWmE
JBZsV6RGpRInjquDxog1KCHfJEakw0CPnY3AyYO8sqsfdiT7PpIHfdcyG2bvi3N4eYHd0Ou4Pgcu
ydL5fAjtbWtafJ+w57uw/SdAi03u+tReZH9WQTYSgWHh+8JhWFP55n/dM9WySPpvcp5Fh2b6yu4t
lvMeNeK5w4o3nafmCFA4Jo0lBklCyibuZCqZktK86e2KF3ipVJogz55VlyhK2ppJEJz8kwfq5xNd
/+fy1OcjeD8dv3iHD8KeEHwRNsdNVBAXYyfJd2MZWWpUDeTfOsfGQ14n2b05nE/GTmod4BtJ7pQI
LFvRpFcGZ1oMcDpe6wQct28fMTjGQOgJcj1QJuRD7VSGojbGPQMGRFlgHNqpirc78WKFJNtTDUbs
6YI7mRAv+D+6dONUoeFz1fi5NBOQa2kz/2ZLirZaGbxxPVmUVx9IvIoNvEfAv/j/jT6m8gv1RqqS
YVcJxto65f86XK12/x2oUqgXjEKBU0ROjMNdl/QZljTrJTW+jwB6u9uOeRWvFYmTrQsYxlRVy8d6
X1g+YP6JgC3pcpQxCWrraNmNnSsjK091gmEiOTA+WfJzaLtQRhq93U9j65e2/CspAYjZfI8E3xbt
swFtLQnxyYoldXPO/hgBoeWoaRHrg6O3z2lTobrVzMoM94ryqMVXPBiTOa8kPLm83MROCBISuGIl
BnSP7QNeUcqWfFrWmGlvMf7NfFIb8XJuIXwb3oMbJr8i5TWyz0/ZQtnKdCkao318zjpjufopsrng
mWZjxBBt4B/e6XECw42xQ4C+Orb8kRvIQi49zj8rp5Q9cjvZjR8+Yew5FXDTHvHgcg26vE0R5mwc
QOLz/8Ho6tGd2l0R8sa0J1HtDZ0zEmLPmZwlEVc9JC7fuQ7XBwCOskQqASR2+1Z8mIpUzSqz2X06
UrjVhOiJvn09mAGdKqGp+yQ4N4G0OroEn9hIkQF53VVG5lgWtYsjc/g+/WC+ClHqtJAUrtY3sbHt
NAqLQmiQdFtoWwE9YwKitWlzXkTKke6zeh9gnSynNs00ixh8hZKKFXAulNcxaek2/rxb8Zs7hh3N
i5DqnE3nK76a/cyy40YJScgmI9KKmfdE/TwS7vl2o1VDtC2O92HmcTSF9KMfVM7PxfjNvBf+t2wh
1+PxmxrDXIyYreMr1CiRNmOZCklIZ6uczbe9ZSVx6LyS5iiOcFedUdPNuk/QMeGOuDbKTHgC7BMd
EgN921YzLlsJXTQ+0q8ZV4X2Ag81oXFMaJnhXSyw6ahMuQONt/Wi/1zxEBNvjOAeZcoPMAkKZrZf
iYs1tVHp9cjaBtMSXTkXN6WKC4KaDcoVPi8kTqJBmtfl2WxDSFCVmxiw9EzvbwCAtfgFtd0UU+HA
JjzBUGT37HNbqijdXP8qrvhDJd5TpmO6i1rNSSTO0DBbXX4lawTM3DykOT1TsZiEp+BgoVY4PjZS
H3bmjtxJTBia+7Gg0wJRDTGJ5Tpsx2WZtlYbVOdNGw/0nMaTUe3AUGs3VJWB683ZD6bqjiAswe8J
JjpjcSTrTjJuouqlpCx+iLtwCbp+dSsVrPvqackpWfvtp5Whl4jXCvku/l9TS2a2oH7bMk7hu4Ur
RtYcDKycM+GJzzWHAAbb/dAwbk5oHCW0DOnSxoRzt1LnJTUUSmuQEWEB9bwgShpxI05L7fPHXgN+
nkqLTEy9RxUNaEI3ZgacEHS//02XDWtmZ05qsAyVLm625e8x/Fu3vYYXEDAafnEpwlohgBKnxIpN
RVeR2tIHL6pU08xBUehSxAkAuhhFPMYICyOUkmk+jN9iDT0TGyCnJAK7z/q3GvTe/v4L5y6kLiLb
BziSGbdhqDnQv5tpDDvFXn18eTfGObiQ7qtaLKgXVtFcMJt8s8kfuxZnACUDAYt26m08JI6MWgDp
tPlpp+BdunZqv7y7m/74lTC26fet9tBP1/ezqd8RSSpnDWH4yiJJRuAX/Eb7TVmLk1hzKXGhxnMJ
J8MS/m3lDiYu1K1nW3eZvtyslqhCXhQD2F3bDca+WZ4TYSDMXxA2P83qdGoDD/Ud5HmDYlhjQDzZ
B99Nmqd90nDgLEZAYzcAnRPmg/vltQDH1hwZNOWOzR/AIiz5dMELDA+hCaLmv7hHdjL0F9JZoBpZ
0eY+jZT3bA+7veSGocRYzpx351sbk3yoo1e4hCdNKLydO6yNkjPykKxIgwlNp7umTgqubcBqCs67
s21ZRimmIAtivJ64j7/pEJJmeIhmyyRDJfsMsjMJwM8KYvKvyry+WtPqqTlIwowOpU6Kc0Zxe7KC
0Npvuvy4CmzzawVESH/BQ8NvomQvM5zw9l4gss6ZfoJtZWl+ilwO9mGD69gS1lZzN70D7BQyONxa
pfFY9Hqx3hIhVDpSPNO8BNWaD6ADOaSV9rO4OXHAcbffVd1uE+B7PQ3+zfvFrv1rjKwvLwRZxyFo
O+sNsAya4B1rwW9ZI6kqTDmGS6Y+/EHSrTa6nllUvOY7ZH2HQgnu5TCwFLm6uJBe6XeS1PHdjGJo
Tq3Thqb4ykEx0lUTgKz5E8JqnDifEsdi6gWnBd7ri7P8+/Buctr+WgaNBA2ET9vjWCMK8TKRlnrY
BfkBHTeaUL5MzQOMYPu4BG4FpYQwjfCsDxWyvg2oddk1EEvY0XqAhvBY3r8aBS/CrM0CBatMY3+8
8QKbs0/d1GDITiTZniuYehblrjeyOGXlRQHYHf5mCTBO2CHDs4iNMvR8nD61RxC5z4yGkVpd+l0c
RYHn1b4Qcsm02mzzq4PgVSbHU7OtRFA/s3VV+Mgiz18RddlBw8tA+iEJdUPMJzYiWPS8QTUWBjBC
m2vf2FWFm7wRKsn+AFt9pI8LVF3vOYlsRN/0ZCvlIfK3EeT/t0VxktNGiefCnqcJEmylRY4H8VB5
kJY6cEjdOVERNXklUaOtkfZehJ3AezPonZSoi7qh0feCU0s1O4eQ9V0aEfMrj7o3ZxhJnD11Iclm
NuzI56ixOua6bqnvnzbEcR6svXTAsT3cQ9VdSH8wGdtp9+BF7e2huc/pvcGb3pcGn05cjHmTdTlA
VtekOEFvRZiXu/5JO3vHTXxKHoAOUSw5767b2rTwXm/EIB4cmd/emIHb/9D2spabgRWsi4KXNIax
dovnZL+hHjDJy2rFLCHArf0zq9wumCtcJMMjBVeKHuF5KDIP1myII3f4tyk+NNG87IVnb1iBfF1Y
ZIcOshLhAOiXMNmD5t+5pZO40IfCfaHr9B6gjt2YfgFSB8vbAxUofoDCy14BXxE8j7v01zOx4JVF
G4AM/+xyNv0g9yiE369WWPnlwNGsOYGbNeqPB5aCz+zMoYc2v3zWCk/eCLKhwXe4nCAWPBjm0q9g
EgAEvcHZFA1PNFmxUerCxr5jffwjQSlOUp5i0wR7nhQnYiXMqx6fmDJbMkxkhrSufbEDu96a5MK3
JluS51J2bYVOx+zUG7GbA9NZIPIMzJ1O4JdyEYSMd58xezZNO93qcsrLCW8cug324M7VCWVcSfC5
WrWV5pPA8rWikoP7c2v8Qe+sdc3wVVdw7pY9oX5TnTp3G95RcI+2mSs8o3eIUGZR5f8ffpMQWbVj
YqscHJe/43E8vfGCM4wxjWN2avO28SsqletJlVf5bYe57R2+OoPP0XklmCPE94pNbPJ0iMS7dsE6
KSKHyKdk6FjK9V/rKCft9SDKTl9Hb5wnKjBsKkER9gxJoTe8RXBTynle1saL6D00IkIRq1/83Kxe
Mb/UxzrjD275wI8adety4IPz9MQlOy9IzJjm1IFsKe2Y5PygOIhY1y2QqvHkHao8CeXCgye28Kds
+Hmi/C0zAcaPJDi7qLa6shwWGBgPGt5W9PcKlqR0/fCPcHHKaXc3Smroliul7YEkjQqEvEe5rt0o
YyWNqSOgSyAlTxl9ZFkrfdGXvA4GiFrDzqKzuNvW7mnc38BqePEsrDLcVIk8qdbehsoL5kvf8OSf
tAB40Mf+ECe9wwkLWtVQjLtgxSELhRmwXkPUbilr2qAzkdPtEhpUipoaIRDIEx3CtFp+eJFL3uQ/
EkXutU3vpCjuj79uDI2MxgwU+dY32RQaLAJzJQPqXeeUuaNDyswi4emfLV1BhSRdjXbO0q2oMfeV
gKaLcg1EP0HcdaW2SSv5PAbzdaF59TrbHxqJ1IwXdwgpb7z+6GUkzlj1gojTfoyL8Ohw42vZupu0
alNeVYSMbyPYlkbf7MfZjnhFLr8ckTebhCq+HsnRiQCCRJy2T5pGyMWXv6Rwy7e/8iUuGEKBwfdU
LgBJsRmZMtaaHwrBXGlLvQhhzTnj68WaLj2pU6LTLRBHswn1IDoGQDZTiMZYbKKCEtxd+LSIl1B7
VsRgcf8W8bz4zu+5Wj8W3Wg7ZNP0m5MKEeAfPSkHy5lcKtawenyAsWz58O8FT5BmEgou/kpUJZDO
7xb71lcPQACHeCp2jQUraIzu/d6E0iKwTzT6RmFJjDTdwv0N0m1poe+Z8nTizXt494d2ImeE4ehT
29hYVmyOx3CEjJPl1iL+4kIkPNXsPketuQZ8HRB5NUhBCYNnH3VbWZ65SkB1x/gVMDoHeUfV138i
jCaLObIpZz0EP8yyZhBpvrZomB5azM4JqcytlI5zvzKE9lFtmvovVNM+txczxpbXzUxwwx92WbEH
fV5sIgYeaEGv7tFvNGGzqbzU6zhjXPyJUGn3ipuYngoVEIQJ7ephTRj4a1JMx5La81S66Va6oiA3
nzZS85G38DjrV9uzGZXkO2rXt9nhqQyks5AzQywZ2mYKPYTPfokbMlZm+OA5+ri70YhNerJ78sAV
IUBAHibcm0sAaKHpRM3K1q3m2UEZSyRlRAhT7TKAQ3vw9qg3+rwqhaFzGQT6dzm0cB77UIEXmUgu
jkl1sfKSoOpAtxSwQDRp14NUUKMBom/XcicshIrHwKoutjtd8kjAVEg3Wepx7fTiOZ9xjE8ap1m6
3w57sTcofR75ufoxgo6Tst+CD+vDoEYd3f7U65KYbgzXSlr3manOj9hG0LDCMIlFWnMHeOklE8EH
2syMgAWOt4s90vaTsakKbhg/SuU5N66kvtt2I+gdbIfNr5XCC5JFQ7wKzO07nxXq2oET7tBsrHrF
RPSCGRnp3FKSey21eCgDqYmHodFPy3QL0ntAra062XJ7QQ8xigWNOPrFecFR27w2iLM5PpvuiAUq
DsY5pEVR05aZgGas6IvajHTpQYsCljPNYcgWcsQvNg8SfvZcrCPyXoUSsenT3wiZcuULMnM88Prj
z2bUJWtIwi8FaCAYFPkndZNFTytL8ocBHYwIHytuQ3VhJDWAy6n65wTfdU6RjW2biNs7NsuAFVtV
mAiruInnGZLYRAX9eGPSVwyyXqL1I/EOEigDAeL+WvdcqL+p4PYfcB+XLb+LHBWF0tX7b8jV4+68
GSw+OWgIFcdiPwZ1nWKSToMTHnpaih1LFlJ54s10pOPNXHgIRpvqA1mUI7QO/nrjh340VkZiF0Xr
W4VzPJhPsp589Ut67LXTjznoKxsfC1M2lFtYZX22iToyu0m8ziasJ/pGZhG2GWUutsbuz02LKn7k
55nFYhAYPM5Och8OmkPUjMlD6RIhFFiemR6wQ4YSejVmLZlk6CcMdyGPNmDqjIDPc+r9je78u/Yf
+hW08SWzR7rYC1uduJ436LJnBGkqUzipQmljDKudAMGcICqdIbgB+GrCX5Ck02r+hOXy/P9wvSXU
hHdBR33f9LtTsiqmDlVNrG3DMKagEqYTPcSVvci1mk3oZogJfOaFRzVreEpiddY2Zn0LQ+2UAVBX
j04sYzANs3a7xpcWQW/FwRwKtxFWHIqlR8Jfy0tUsp15uKpqvWWEGpnl4y2JyqrsAufKcW4sRMHd
1+1JCcxgRuNGEUNFtHrk1JyQQBA5xZswXESW/7Wu44/mbJ+mp4rAqwJWgJkZ39NHNT3HCN20uL2F
whm6YFV6WYEr7LXcvO7/JDaCOZpKtPNx07yyAbTG53tXApLEe1faccaY0q/mmZi3qFbf/fy6PkLM
1LpI/faU8Ycjg1nRq4/sCbJhmwfIP7ry3URttkRC8sGMKvOSNkwNQYSbS2FeGWParuUGBktYQ8eg
o5gHx1Q96+5x6JAQ5o00yvAVlTX0xCkyim/X7Jtlo8dP1sPURMkSK/L2bB7szoyj2FVu7S1Yk9of
UYtGGjPxViLN4XKIgiH4nxduVo7d/xx0674iMt9trGtoSBbA8kQ/tu7FzQNrOlN7qkYdtR0/+Cqa
6nqO+fM+Gia1SDjMgEV6Z+0jT6Vi7Wgys2CpSau9oY//+6eZhKwkavy2gugKtFLv4U6oTzILIdr/
cQ7fdNOIoMlQpalwHd5RGQccisENeyIckW9eZagrL6u0uzjO9sa586FEi4yR1lOhszb6VgqEol0K
Jewmd2oaOCMBUQZ7U5f023KTMMH/WcGiuG8jUXo5FlQB9x4wAn6t/u9M59wQuk5RGO/aRmNFPQA6
5WlbxRN0F2+kXaxDKH4DVntZ+WE4JMrbNhBckX+VpvvK36vO3sU3Wr0N3wP0hHIeWL8hl7RuLxDA
xTUcQRTBSkIZucIrT1Bvul3fDz27MQYzV4xgTsfF5sY67IEDC1yWhVUBT1C7J6PgKZhyGUobF2UN
Md4AkyjRf6BxlTHk+NBjqdL7jggGfyAT564qMPLV3ynjK19JhrOCkfCr68/M7un0VFj2XSaABhYi
M8rWfJnoPuc38kxQORuN6kU873s7NwBiGcgqPAeNZ7D9nGZ3MSGl3MmfpXADGyExUwkMLiunk7+A
j09vwj42y8ufrbMvPWsVCCMdVJWl1mL0GAqfqexrkH2FNo91Y0AM7f60JiymPLGhEQ4lwE2mxgc1
tQJ1p5FyvDLw705G+FPWEOOy+kRtCdLgFIu12fO4woa2VyWhYZOFG897DkiDUTch5gaTl60H5xya
vSThwPV+yyRuuzagI25v6KF006c0F4T92SO5k3p/7ur6e7fDSpL5/VvIzbmXve3a4JCJxeoC4vU8
lFOQ1xxiVajCjLGlYYZiZy+yh8S7LwJPktenmShn4MfDHBCiAr5FkkPHSdfQee7PglEMcWJEMblj
OyHBvccZu/9vI9uj1bnEqvX+vw6F4yHMK2JdA86YHYtbijlrpF0goOmztz/fraJdV18eY9k6ejOZ
fYVM7F12pOx7paBn5e+qAManMhp1OT1GEKpD5xNqvcXNuticCpKb2uC7VE2e0vpuRDPs+IO5ZFUU
K+wAtOP34byGHPwxCGBrTH/eOzHRb08YXRyJJhVrPub0/31zUU2YU2Bzpez5h4XfWI9CQ/jruS2Q
SH1LepVcSuxTKJkxxGiaEnUW0JdlFNFDJQ0R6R8lXjTVNZCW0xKORDyzv7NYie5gEr3d9P/0UE5p
YYNONAjVts9ox1cV4n4isQHjVxbZ9a0huVvDt8k4vtthuNtNrOzA2LsAmfT2of5vGq7e39Jtfjjk
gcfYhKKqEH20bzyFQ9b9p8N/2A6c7l5Vb0T1dF6o8Wz0QQPZR/CX/zn02Fn42ZhzaLypfqH9oysJ
qpIwFGJAtb11UWJcHurBCAKeUEx0TwZFULiPbcY8M7Jj396o92M8CaAlamT/MYZ2PQksbTe1JsNt
ujqmMsQNbvx+9FYaHQUq54kTAQMUgMRGWVzfHf/vmABXUq7WywHv4lfjcoqe5vysOj7oN6Yfa8+9
F1ch0A9Rj0oxVee+/ckvAEwBSXwZP/Ft/NAwQ/pUIdiyaTcElfiT25Pq+H+cI9IzW3QLEkVKfd9Z
AGe1v7JDhiq2GjiDJ49eP1HVoQvId4zxBnfhW9B6q3wk5tUOjc6kylky620lLtbFxKKpewX295dJ
TwoLopBs2IZbpQJhceXAUPHC0aQFk8emLHL1Xd9NQ9RVNblaymMgAPpKocgJjbR93valPKltrrAB
wjcy7pSmFdgC9ScWm7ymWRGN93gVTrvYfMZ5bKkovI5V7IiOScIgue6R5LuD32qsYV4UeA+3UYrC
h2sBIEKXyTUZNKYigZZVSh7fKszUwVC5sGxWOu/ctH01UANl/fNQoAoUhUe4YQ+uIEWqkGmXfNgl
5629aPLXQSLjo8TC+gIWfId+iJnKvYay7Rd0MNQdrTWIHXzf6gPXoI2Kb2HFp5fHadY7PQ1KfI3a
DZh7vlP3KFkCqV+dx9Q25jYz8i1w4SVadzFtlOIxGo67RPXLfDOf47WDMcl5Jzusl6Do12fwkAzS
DU/kEhmvZCRd9CD/mmvngZM0QBBHQPcC8TXx/y8qbddWGF/pa3bnyrUC23XoWCOv+mKo2uFaG+zE
SO4INIjXM0NplZt8zrzGQvK4ohZ4YhlTMuCszGe1ytVIKvF1BD24g4SOiFlNMs75sd90elLe+MCM
wGChcvTgBIslq85M++4PSt4AyB73uByaS+G6hLsuyLilLDGWx4fw+HCGHz8tcyCrbyE2ltfWoocd
Fct8YoVLSOaUbZM62dXtlAtGGv42ldp8gYpX6+BvVPETzpzUvu1sxdkFOEOvUUErH3ofztfQmqcJ
KjScmcfW7DWG5yyI1WPssDjKFyIs4Cp4XvmtQhM/vbPKovhsdnpZ/GzXM4F9WDbhh6MrOo1nVdbC
6mk2mmC7NOZ7/fNJwUcHHK+itdV8fACGPx3mkK+Q5F/T3ic7JDmOpHm6ZZzBR5M9Ep5/dyKDd+tN
ng0FYdI+EoRYjo++DqTQWvB545y7C6TdPjNtAJ518K4zRz5LuO6GcHR+zFktq0+EeDQ8+/1fXfoS
PI7KuDVL2enZlNozktIawLpbNKVZVMMi6Xf2VnPp5+LTCCMgsrPsHBWhVcBgb0PAYsMyw1W/+j7W
4bXCsNQaV8N5ZjmIHyMQWR55hvUVbq+qDQlMIJEHdJvBiU99MAiSTUAlZ+2s3AOuHpFmH638MHX/
5hKTZcU+W7UoPjzhcVcbx5LgoMEZUZMNKccI2WVrkyF6nsf1ABeqtjhDGsKDnT5yk8pPEwB80Uc0
YsIPIieosl6n9TqOaGpXrP75Ak0e6/+GOFtS4EQY/0sHU9+uZKh9hkGO14VatIkD5gZVWSmKJYX/
Ma7RJL7yzW7aTqOSR6UeSBMBzvGN7ITP/4a/k6PZMlHvBaAJ/yOOi0RX2xoYqDMxApt4Df3Mc8Ml
K6IcuPpw7/fEMv9LVHF4vdqgMKCBr8saObkdbx3s+FHVcZuYIWiXy4nEQAPsZ/hAo4qwUKdzt0Qb
3KgLzqOHMjpKK50gfr+outmROm4+kwiHswBNStNjHW3b9iXlEqYtvHeBUJ6VzTbkiMXa2DyGq0Yv
trnxAqbBErgWrwcmxKUnimkQB8VUmroU1DMORzSzkSjaGx3uT04bDKwffVhrtX1Rt2KPw+TIJET1
TqUbRQlVTopeVRyf7XZB7b/TingAfIIceFNr0EQR10iApEzOUGwPpl+dp7mWeTUQWjFNLW5VcODm
EhMCOCyYqi2KsprMdmHGh+pcF5WQgSL5d0tXlPrGZJO7IsG1Sk6E8cgP+pS6YyT1lO769M9gFNPW
fmLyIStCJY8xC7HBaisva2b/5liNB4tVH64wOEB/icT/1fp6+a97enCmlerke+4fguAcnm6/V+Mf
LveOujCqI3y0glq3O8ir36/wMG6+wV30SQwGiPUIDXvPPabj7FJjwK+Xf/T2ejaz6w76zvBnknIk
aIZUX8VprzgQ4UCVJSAgbyQMtweBjmyvcmEJQNRGkPL+aikeDFnqHDDkwE99Q/m/pG7TBOC9aViw
F7+W6dKvBpaMXpVKpGt6TcyLJNwr9S283utILH66sCeN1wcXCxEM1bL5lrftwAiBXKfm//CH8QJR
4mjnzh5DbnDCoPCnkGxUl3iLH2tt9KEmvxOFaoFXOLlSg9LD3jFTOEHuNeImNJgn2tCPNWoThZIn
AM9ooXuSt6x2ERao6oaX41SS5e8mRxLGvaT49/83e5pA/3OklDeEK5APCGQ+1mOyKbhE/OwhpUKK
OUZ7dRU0rCpdTLg+09IS+rbLCAorwLYUyvEP9Bm/cjS7pBU2u3GIg736YksaIKFvUrIEjUscqPQp
qpsNJt3ArxGmg52l+KQdZLh4Z6S8e069NezdoidbGCXLD5Y/mulUIdA+ixIS2HtGKECbtHjcuxFE
4MNI4iVG40jxRcNncmmE45/1pp0d47GUVJ7tczaQS2coGvux9tCxsWgo1uqmjvN/pAgCZ8bm0wKx
zvXXmuwjPKDzrvCdE9QubBpPN+S31Zs6NSNZ5dT79+IBG/g/RvhXUOCwl5hlSd8KBfyvC1Rq74NF
n3fLGqJM01mVotbjnnjX9Zil+yZKBOGIZRTY1xXX48bQL8F0jSFJ7J7zGaJZUP/DgFmsiOdyelqW
kml93hbgWzmQLPjwvVzTDA6PrZl7Y83xFwOMZyf1mLeNXR3ANit6Pq7paDhep5qjq5xe5lSsejrT
zvFBrVwWBIr67o4lcPWhZveQpXPJ0U1t1S5lOiEXlrA9zGvtDkKDjeMHckGjihq4/5gjvndqSfd/
egCLcEipfwGwAE72/rs8e9ZEAH/+n0+3A3Bs5kqxNeEQ47AQ8bbJ8vEgTR3Lbhdn5+V74FrcVpCF
D3x+5x+wnuXC4x0+3+Oj5ZPgLMN5/2sSvSk4Vz7/1zDSESMpqq6ec+rPNxkyb9LFM5b8pdhw9UzP
jDMxxVZzI/Ir74p5gPSNpZmwtBELE4EeCAX34HfoaJj5QoIRvexeNO47KibuauzZZqlTm9O06sIu
OaOrnxiYhrh/SYqezKnyJBED0pZKKMy5wiXBXzVIHIZ02pLhEMWbUeKBgYYVgfhvW6RFdd+j+vRm
C/U2VIoL0rKdNiE0lFbrnFXGvF/mPiAh9KqcJqfy7doVPLjW6+XnoZjoGYeIUQ8R+msManmY2f9h
FaUcQGNW2/V2BDfE2sMJHVonKY3whNkM3jvDzxWMee6xOHPt36BKtCtWgFIwPEvcYlEAInLtmcDp
gLP8yJLzU0zJ9XtpLva7Hy73oq5NQm6s60AaYNUr82fA6i/fW/9Q6Qu4PdR/ZH5+FejvZXlC3Kyr
zveFmE5ao3TmSvyQhN+RCLVj124VQoJsnCfzt3S3xScAIwYFO1V2qtFP6oZp/ow25jZzMr1blmJ+
eHJ9PHlAPF2qGjr/LLrSo9budzObblJGSpbejQk6kedN/oCIil8s79A3ThU3QEvkvzGhokdDYgcP
n7JHqXoNWgUrBh/63Chl/9/vXhfIi9SYtaPqZQmFKpRd0x47oXOsLwLIGeEM0FPmVHuc3JI9d7l2
wIFLISl7I8cSjc7oQAY6iKEz7B9hYj8KnPlsIGvYL+sWwFrwFH/6ri3Wuel5jF+2dKyRUrXkqjGr
PMdxT+yMkuE6h3TkesMI3pImUXBKFMDXqdKeihvB7Mu2mzfFQvgGRP/2T7Pq6f8pOBGs6Xr17YzZ
Wcwas5m9K5IaWxzHan7spKb9H/RO/l+nrGhPyzIMsDkQtN1Rbaqxd0AIgEYu1hPWxQagQvB4PJTx
rDBCa6+TBgMihX2txhzwJ7ryE/GFnzNi7QPbVNJ3x7jYqMDa4GnFUguMS521l8geG5ZUz3rqqvk1
Trrj0LHbudMu43k3sd3F1vcB6zs4vt82gYn0a/tI5Bvd0yyB4/ue5KYOcr6FmaD5Fiom/OmJmEO4
M0pFhho/+mTNXvUKRDcHPXGvzDXhaNZpYCa2NgerqQhyOEj4jGgotL6QWIbHqB02M7AS9RZ8u8pg
7yytSJTVJfUBUvMAYVc8XRHNbi0vFB+jiFS194uZ8Jknt3khmrBZp7gUqTo53xQecJWUNwWqb79y
Hnc023+C7ewxPze/TwXZ7V1aMRjxpQt+XpTRS6Scl81DVCba7VuQH9AtNNkIE7TWwECvKCddj9wz
RzXLPW4S7+sTGTkjRomV9KXsHFpscS9P65l+pekllJjuKJYcES9S7HUe+XNRhF/HYReYPUvcYMep
FffO3Zom911er7jGiyvHv6yxWJOv10/Gx0y1td+uQVTZQJZGCy9NqyN9Z1FJoNXjOyrbyS1MCVtO
kLgTUqfdhlTtBHItFddhfRArAtocWxJ+XdZYnmLcokbIlgxxJ1MGmnNBlIIqyUr4qc8DgwISBP1R
MbcnWKy1ce8SJnUYrLsyora3sBFtP3nwdwU6kbiD5DLyez32qSaHWdhu+NEgT0UTjpwuJV4hkVOW
Aa0YqKJj6AaL0uaz1WVLDMtukpheYiF/WuVKpNfrg1Iaj+BH5QHASRP3vxnWbKZONNtv0zxAp6k8
EkkQgpwNrl5tO1P2SMwGSCN81jNsc8NLGEE2e5EabVMdyAoxQW/PDpI2Mb7w8KhpOIzD9w5Tl6eV
Pdgdyg8IchL0LuYg4L6Fs3uoeEFBq3LmV8+/4os4vvLPTJZFYbsERtT+SnZJMtSRDpU+juuRgMbW
NAH+lcblAUl8QIUWlMzRg6CzhmzZjsUbgjhNXfCxy6m/vDdZf00u3Wf8VJ5wuE3AQg3/mNU5Bb/u
Fwq9pdqRSTDHF29SISYnf4f4s/KFS8evYiihtj/+fewjmn6lGAxHKtdNjZTOve28HVVNgTaOWBfd
99ACNIymx7evYui8KQtaye84XgcLr++ZGvlVRw8lgyFntaROk8+KTVTFP5H8JNkgtvivVY448ZZP
faGyoSo0FuW5EkwlZK/kcq0vwvNZYnm54LuCUNRbKnz6W6yQCRZd3aOXX80B3uYVwv5+WToU4v4Z
XxIazjbIxYge7V3PNzPRiNIZMMiZYWmfDwObXBfy6p9f+/mBBNpbgSSAch/k01CmGXW3p7Ut1ZTS
CPXXz0hAlXx4VSwKK+dTQrbFwOYksaVq2H0toa+zRCy23Zz2mzU5C95++hCIn/ozrewLOW2PygLJ
z2fNA9RVAeLX+HiRGem1LoOWocLcfittvKnjEDWlx88jujYIrlnrJ2Tt3b/iXyK2XSyu6tMFr8Mt
Uqc5EYYXxLcP0/CcgWiDzWvzx3jG/L2uFFwM61CIWOjLsM3JqQSxbKN/FkU/+er1GGT8PzZBZX49
WnqsRAlyMP11Gk+vjHTBMZAdjtt/CZIXJ/SdIohYVmevkwOGVYVAVcC/w9ZUTJOKJOnyDcOtgRiA
o5C64uPl/7PatWriVlIzqqkyH/MLnopkadcBdBQ/u2zXOhrYcnbqtxgBHEceSs3nysyeQvTLTW8S
ryHhKKzq59ZcIhmqIEP+HFRqHe5bNulwU+R9yqwPe82ZF0S60dnjWJbvm7JDqZzd5pVlSgqg9iWZ
aJqKtNKjEjsdJXJknf8E1meX6MVlFY9LG15XjkiXSnGFUFq5q7g1Z85ikenCBLM3OgffROjTTGR+
LHFrTCveOQtMGg/ZKeCrQRWOpMadjfI2ah/38rJlXCjyZadLrAeWHE52P7xkl4viRb35DnF40j3I
DamYAp7jGPUhL8ftDAswc+EetEdaHYcGbfhmEoXUbKnD5v92u6eolTBOqT9FzXIXtwElzL4B3i9q
aE8UXPkkFm3Jx/O4x5/SfJRPJoaCp+h2s5mAhjQXF17UbnEaAjiNOGCumt6OHDMhWiwRTaZYA2wq
86Qr5jIoCspp6s6iBsEwJRvwMmTQs5bLId2NiwfG/4lzQ+ghqv6doktTtqXjjc+6XpxjkEHHLUr7
evPYumqPKd5h0sBFgHSJKQCAxe08BVsv1Zp9tNQ9cPvfpTDtb9y04Glx8tcmijJWRV6a5uK0dtdp
NAsW4CFPH40nlMri+ASY9MoJlYmeOJnHya3pi48TieRO1qOZUbrdsgnte1+YI18Hd2joIDRtYkgX
gKw4LnDZEYbH0DvOs4BU3y9goS5Pczrnd4HvE7vUOtaHdogUObh+n1KJzehv4v2LXy+95XlDIPHa
+8rqt8awvvcisHarc6yhM+JyawQeWJ2TOeaEs3pdiNNlSpc2eXE+GSc8kpK+Or5UXjcY/Q21wmXg
87KxLHeXFMd3fTb7wjzdv/YTljoWt5KP8x5l+K+R+VsTTPIOztsY57h5yJMiW8SayB5RnM/41lGy
ks0/OAWaAVD3NNZTr0j6uLiYSCO10A1dxtnobIjm+rLyvKctGpk1iWHoMfQi3AiHtQraL0yqjvzV
eqyRdrvfk1RM1HhWFNgQascFKNNGlUo0EvOMaBGHMMz85N8plgG+B/RFJTwwHHFTUpC66L1izOtf
BoMO9eZK+xyDjcjKOW14mva7OuWs0rdSguR8k3hNrJ0st1OxNS4bBVogx5NcaAnuUpsH1X2KahHH
+9+38dS9Mvi/hasClJ1tFJqogPGq5jStcjtwFQHmiWJQf0aeZDuCHArbVpNdGnrxD97WtbpCBT7t
25GN6fN5JL5yoHq+hNyy6lIVsnqJweYKzKvAgclEySe/bn6OxakpecS8C5aG+a08A5iXlklJASxt
1sWuXoTSp90JMmQFhcWqFfTd3wfkI02Znbb47VOuv5bcd0iqy0M+QqCabBtCl8jABoPuJst0zXOD
vS+Pmi/+7oomyJe3jTS3+5KpRhT6w4F7e1SuzchDn7aiEw8+3T4kQbHZX5woheAzdHxWfzGLv17K
KNC7cmK9tTAVw68NvMKdDHVBNlMrLvUDK3RpZTgaST0VRb6O+GdabV3eE+G1EjcW8oF4hLxjooKO
BS9LmGU12uxN7iRmq/aNTHfVK0jNgswHeVxPLiwxGSMGcvHzIUld0wPteaEZprAv+nMXkdDwn9r7
gpd81TOl7pksSGYcEZLCBZtpOCax+ZqgioOhhaq96y8B137bf0fmFEq/SCYQDxq1q4gp1CBSMpPn
CxetqwW65GhdOidDD5RQ1SREtZP1qxzzKIzpHCwx5N/h5iHnsKBzQck9xZaAewMm74N7q4/ewDwb
4ulyWl6671S/FhwPepX/fh2CCzca0jaaPAeB9aeGjq/hrBi20nCYE+nliLF7hkaa6d62FBBl7XWc
fvrKlgpPWrSzoEjIPJd/P9uFhwTuoCZofaV43cKqGfMRg+YU9PJaxVk3cnsR3DNVETQKsXJmBvzj
RqmD0cHDTQtv9qPUf6VLUrc1BgoOZuQWh7Qi7BLqhHNe8Ga5zXMePrArLxMClwiv8g0Sw0TDquCh
OQeTU5tdpR06+aV7EiaRSm7Ph2a9vukfOErlFnPPIIg5p1U6rnpkgoNCZTrCWMWzfT2oeCNcKFSl
Ag5NRaV8HPlUzJOI7uq8eLJQdPBbRngWl0bjO6XtvNwocX5q+pikPNqE+4advnfFnlARpia3/09x
CKhH/fqrdWL/dWcrjtP0ffIJgBUs+vqzcVSQHcfW3hXvawXb/Wr3WgTMCu+QI3NL5mWHvifrUlPm
bgjORa8SKKodKkWDBwDGGlDMaOakZwIo5T9vPBQ8o96TiWbiNu6d4xezw3nr1nKoj13fwLwhJzFu
u6KAySkU/rEkMbUMC2P1CNm57BKIkBno4Enp+gZDou4A42T/YOhEP9PnV9F6VICnaWFnjnbP64oq
zZFTQVLb3AEcYCGoT37J+EqYAwl/oKv4+OCXFjRuDNtxyyj8Rw0GZlpCpM43I+r+h+kPkrY3ldKs
dFXXqL0ko4YR4j38EEU7b34udl9TTtvuNj78lzopFMpStQ/+4KhStcLb0NQaTdu6L17XBYXkXFuq
fei2cFE03DH7faSddtpBjqGtjWW/mKS9A6L5b09HrgH/FrRm4Lo+E0YeLA1iQA2+ZWp8Ll93B71w
F+Wg0zI26TE60XbPXcPaNx1BsPBpj3tavzmv26jt6tubrD94rkkx+jMEnFehmoFbxtoREwpckWFQ
queM15NbgPpSkmNxoXTLfu3L4TbQ0obCABiuDtNuMHgbFzUnk9DcT/cPYPTCpBXJHTDpQVQpy5y+
wJ19x+/77xdnNVYUKU0s5l9zeCJtE42MniQN3DnGKo1tfy4FaTkf4EIjks1jETJ4lXkZYIpYKZLv
GEOUgjy6vbM2/6qhu4umpP9J1AU1J9dxxN71e544puDXdfxykXhp3HZ7t/W7pdpPtURlyvWlxXeS
6V6VmC5ykDjzJhdNPgojDlbsL3kbrQzLW5CREUOPZWbuneh6Gsze51MXbFhjxSb0ZevU3JM05TiG
HIWLyebOezrsmWxK5z4r25/L0zPhlSAivpCgstrRKgbD33IxdrSZBnD2pr3F5kIhLvwwzzylUUuw
r0yt1ibIMU3c+Sr2am/Gz+9GhqJS7hZCoG+CFQna0MP/7dS7ogWuRmX60GMna1915Jfd510K00xu
+oe2ByENUePrEE4IY5MkU++1tfg1luOcJI58+Mg5a7iVu+YjvluPDb1sA67wZlHri4xLiiBBxfk+
v27SfbNO5Ffw4Yru9p+0nMF+SaeWczFkBKdQICelz0nUmFxF+wGz8F/nSDNJ/cA149I4Wq/uHOVe
uTFpO7TWY5fJlCqaBQC6YPfW3XB6KifKGkhbH1sq3uSE4UT3LDW6KLqpWprV5LgCu/n/S0YZeYNT
IjqRoEdE7Yodk53Rykp4umY/qLFQO3WMj6mDBvw2PBIolU9Q++fOuBZbSWFqNyM9JTtg2gSOuMhy
1ml+DTGQFFzIhjhp6Rrg3+f9CoF9SKz+3gd7gevThaBuP77wSF4eeuc6sA9ti33y9ZIHJln4OJWV
FPrr5IjA2+QjpG4c0diFAk/VIP7RcdNCE7vN3493ytIaaL1C5brsnYt3RBU+0/oLqSPxdvTFhFdF
+LKYK2WCTXAtcME5yhy19j+Jkn9lOZI7MRSdPZCLTT9n8TzXgkoe4PpovpaeDq1HWdooQm5jUHf1
kA5UZ+6pVw/XFw0cdbmA7lJVmmt0dcBqeoGH17NPwEmAbWzvoBzKcRibBurCTl5zRFtHbR1k0YSC
/VmoboH5kJHQ6eVaYXOsEsIY2kcTBRsiyHYyVz67jmIZCqb/T8OYJOsik+EJuyFj6v10jcroO3vf
y8fz+t1pBfPnEg4DHbIpHxwh+y7szo+e+w3TFx1P7iJDm8hPd9w6nfEI2i3M+pAxR+k9Vfer0ICA
ysCsGaPD73dc4FdbZRXK47RvA1pWKngcZz1PvIj2asquORBBOKG48t6NkyKOw4BvJEjJzb4OB4bd
8hLsVFnh8oiQdLuW8fhHJH/ctEBj+4TEg+RBwLcPrh02t8xCTlyGIYnqi3p6r/MqPgT/y0r9Lr/9
qc806n4kkSAvXm7MsQ+F2KZ84odtt6Xcdinrf7/heiSa4xerogRSKbOtFjfXiJXWf9DA4yRAFG6K
1FT/6w2Iz8LRRYODxO7tpZEx1xb0ogEJIBmoaqGBf8j8JN2LJrgW8ZFjpooCAXB/2c3dMYGADEgp
Yn2Nazt3GrhS4+r88a57iYMlUDAXqA+iSeZVGAXfQqKW9LLgrWKJN97disTlerQxdabQoD8jNVw7
zTiy5CvcrenK3eYyamMpFke+Lfv+S77a2AYp48zv/QCP/RnW5M2ro3DiXQ2s4c5uI62+IigRpi7b
BdCrrWWX129dmnt1D/HUpK0mC2vTKB7balpt6q/l6gM5rk35CrCzQ7iLoBi2ngGIAcjTsU4/s/GM
ze60jtLsMRWRifpgx5oRYdinjYh7aTbZW/pFMxRSwt7FIQk2IMjovYiUD+04u0TwNf8NsDYAH0w1
PIFdCLMx3t+IdjiMHmZtrmlYbsX0WW3mX2eC03YKiKLbShOWyV6UKMN83jkXwJ7yd5DYL1z95IOT
MA12qusJ0N/NwcQBFD2t62GpdrAF5mhzhrqgyceM2cK1dUJ+je5YtP3+EG8YOFLU6DJlQHgNBLBB
DjY7MDmEm0rTDGT7kkwNA5mRr9hO/e04MJcXHYmzNMxjDG+6ML2rI6MzUuHt3Ka81/LNXEvV0GcP
0yfuE0vJXnRljdxuHN8rCy80c1LtkmGWIOX4qSah+QfAUPgn4lIPs4z/J59jK2NlQUHH7zwgaGFc
6OexLNTCqitv3bbZorVyycnY3h6wTd7or97SCQG2SzUldlXhFGF5CWmCmCModO7QjgI4wQM+eecK
orItwL+FI7AYnmNoC0+NmEoB4uAQT7mq8WGmhBPxMLCRGUoQDadMxYYz/EP3mLt7f/kccrR/kKst
PgGQYaEcXMC5xsZg9OIPEZ0IeNIQBRjvtrSAJUidpod0FlXH+gAdWYIjAbBE6tMLtP54reLx8CHL
gycgU+SH730pGfbssNTOsi9XQvlDfIbLtyQ5A4JL7lRqAe15csHGKRgmuWi3pHuAw9MFuwaRpi1M
ZMK/cB5oJkfI20cUxEAf7T8o9TnUKslw69uL5I/ANaor+tx6QMvCj9XsjBJ9MZDiU3aABKus0C2X
Ugnc/yzqTgfwuZwc8jS4Q32QMlpa3fDScDXZr2YY3h35E+iGAEiX5SHjGFHKu3L54x7LXRzJcdeL
eBs/jOtUtmbRrDBxn1J6KqAxdJBWirQgYsafv67BJWx2ncFlRCjJab96iBzeXjkpeEzBluPGHZ7d
LFL/BO50da64vxXHR7qp0xichHA9xvtIzJZCM1WdEx1HHsbu7lfaE1L77+hGI9mHSs6fKYH+deOy
P7IIs6iymSOpdC+M9m2cLXVXdNKInJ32e3FK1KowvWP9EeVV2FTrO6bZDEZ9nvsNJFnZ7MVpsmXS
hKP7sev5tOfqt5yGqTLafHPb9tofb+jSMYN8tvYqnL9Sfp8ucFJnROSR51eh8peU5NYU6FR5mjIm
G35ML5kstlqskeCIIxlc0yM+Sg57zvAneZ78CWRdPywFlDH3uZZpeVrgO6KhTKCpw7u7Pb9Jhr8f
kX31h2pdfzr20ojFumNooW/GecTeMZq/BCSMmnl8m8xF/GaE5qNVXwJWCRo5/VHVOb0OMZsdNscj
gVVvkjbSR/mUVM2NarkftAEt0zrXuElov2YvcK5aNxT5Nye/xqWp667Y/6XF7y3BmLvZp/YNe0LM
ddSAgyZefLeMRDuD55OaOYL3YWNwg/u5CEMHRKUBIdk9m7itqM0fslN3x2vnD02YIaecpTkzhaW2
r+X40uvJmTH8j9uBLDGIxJb+VfUo1G/3wRn51nOWqo+NcavmrnNOu4zdWIiVKVyCm9q7PFnZpvrg
LWQexa4JKEjkoGbaITBoH5qrEK/uLCHV0SgyEN17bRqCFVd6+nOHg/FfO34bQRwXIEj/mmCCgxEY
7m3YCDj7BxGWnuIIh3hkGy0+s+sMUNpGcfr8XjGusuruG6GvlpUrbkF8ceXBTJUeupqBPRoyfGJy
T0u1csq9N2isd8abvZ30v3IrmERbX3FA+cK+kret5Ng/4dTui1Y2LBOYYkD4YHIn69nZhR9eSB3h
bRSL+DdpqH4LQz41xeOI49VYSO4MZJh127iYEHJUkGK7Q2Jf9K99db80ELLPpueTuLR71KfS/N70
ZLed9yDwCuGWbmziBhKcEb53sHm08X5Wx4ChUobGilIiHDa47v+bLXE0JzpWScYO8C9irBomS9Rm
mDNYHOh3x1awtxQsf3WLcl2qVwarWEAEHg1S+qWuTUTbzbYGmOY1A7kmVhaemhY46On3sa5Ecx6g
p0KkutIKNKWm4FHQZqGg+/rRGfHz+nSQkbjkBTPZzoFHlI0Or72rWIMjOeI/JxgO4lhJ5Y6tB2UG
g4I3hQJxZXzvuhTzp9WR/uuFNvAcHLhRiSn7EgU2+a4z6BpNVnRe9JKoJN2me/F5BdrYBpf76uMs
bj5AbnRI7QbUp1+MU4viFumdEpJzlYShtNEpyFO7vQWCfWBknWugwP+B3GObHTgew0QdHJ7jEGEf
IdKDBfK/rvXCPODBZwkoBAr8kSzkUW9NG+1EJL+AGmb8JM2kcoqFurIUm7PJLohP1UlTHiaeSfn/
cNhQ1PBHHIQ4M9FBq2wLT0R2z7GoM4ZYSByCkkUKeG/Bg0XFR+9Klbw6tWpMqBd/Bk8j3TeK/lJc
WMmsZbDsP7rKOrsdKYO+ciyJ5LS7gstRxCc6W53Qw9nkCo3mrae5NY9/Xs3ytRt814sOE/1YWDTA
Jj57x3b1Ue4aDPn1oSsIPh5t7eXTrLdKyhVyIsFr/Fuhmvwys9bnb4ppUzefKroFF8uqX3kXHk8t
fvMewwL/xpYmKRMPK2GnNYHs9X3Oypypuc3COsUhwp5H0y/WQLY5h2Tx0FtId3VJEonQ+p4nxNEr
4R/Q02pCZb32ircPLlfcYFYgvPhuc6mFeYRyLw8w/c2JXIqeRWYk4Seq8f0PgbRg/Rq4lJHeQifM
/yux43AUqLpRRYaTtu/Zda19Mm+a1CEcwQyq0aDEoSRoqxZkmn47SskIfahUi2E5E9waIh8i0VU7
MHvIRZrHOvxLhTVjpNFA6HGmwo88b2kxc7Ypd/SiHoIVdY4fQ5n0LlZcnjb/PL+fHZcZea9N51EY
XuUxP9K+uco9yW/rsW0LrCmAstI+yA5zA2nkp8mli1o4OHFlr++/gK3nDpDcYJZWDrf4fW4K60vH
1Rle6U9osiNqciua1+siIJz6W47hOcfqXzB33jInuMQp2AUsSoVbgAXlAruLTXvHUO9v0TzjPL9h
Xkg7AiG0HD9wSraA4EBM2F6N6XrtpyCGcwWL8WmPQ9VVICFaccBKtr7OU76x8PYzh/RuUU67g1Bo
3CjolPxprmAqW55R+OU2j7qNVeXar3fMm7j+h8wY2G1lsKN21qsif+NA1QBzL44rDSpKYTPINEJ8
V2oUPU4bdi4G8hbNYZXCgWe5pJssiwUyAqDAM1P4VfRWvF3EC+2KGz8GPARtTfycIzPNcMtTCb5Q
1pLY6afPlS98vBXuBsAlultNBWfXTPyW2uPH03ZXNtaKCz3ihBRo33QcWushg2aVo4IIjQYvtx22
8Xkm6FJKpWc93ihy0P6hGGj1UwhadRDMsaGEIRcZHMYEQK4fvQseBUuTadua0OX2cwNlPqBC9oFJ
4P0YA9NNPpg/0AHYd81iUVQF+afk7Z9kRdfgrVESaDL/MDcz17/rjd71Bl4Co792Lixjgl8IAQln
A3fy/HSjIzSQf7YPbxnCnHmOUPDUMZlJRYubXshmnHssz52B7MOvJPIl3chSOOrTIekB/qS/LpAl
0mrbcPCnsYw0n2PYCE8K8HQ/VhGYRaSi/0iUjMI+tY8Rxqo5ZqVqmXxQoLNrnw6DTCslAhcdSapi
Od8L+SvFBy+jFH+sVrKUZ2Twu+2btX+Q4GZxDdB+wOFKKKwxDjJ3w27tiEqT4A4dj15NSNZ1PMx7
b4luGR+C7yOTlTIkgXVUG4+bB95dnzXXHXUzi7TGXn3kmPv8mrf1VX7to6gbvpxKt43GteN9GFBK
bWkDm04pOxvkq/YbtDE1tCIbKhaPpSq1nadZiFs26ysLl8gn8EL1ZnOHKV/qRYHqw6Ze86z130jk
s5ulW60dNxyjPu5zfk7iKYhu5TOVYvmGL1R5xDwLgjuXVBhc6ZoJHW+evLUmQmmeVDO1CuTvLYUh
ilGMyfVfN7fTzOjXwMhp9bDBnhgDHhe82zqIPZmOqhLHZ0+naWNVJEtIz5/gYDTRdxyDAxwonMoQ
5tUmwIVPy3BbHgsBLclXPD/gkNbJkQE2b5n5oaVatSPH/qrd/AQpMn03hDuBqUN2aJOHUqgTCL3B
YcDZEXARsEm3i67YAfO/isI+75Z+N7WPPW1hUkyLAFQoCRrbnsso/me4oQd/90cLXw4w78K3Pr3W
H85/q/JuhZLdFKQ1bHZfJwwcN+tYFoLsT4N8xHq3ioHlgwYFdt1RL2aGsFwGQ6lEPplR5r0vB2qr
qFn8xK2ISxOXYUpBXJLDr1ZLA0la2/5NKgKGDZUhtlDTBgHBbsWkJCYK6OLvxfVE9b55VDBsp6S8
F4NzRWbUmDbntlVnHAXGV70wgVDUXFa1ItDRhrOVDxMgwlkqrF2W78kPGzgqf82kwm2J/WLyBx5U
+Bcc3MlNI/KqNUIrS8HLGWIT0S+G496/Qi4FR/bwDbqmFqhQZDEXvqh6hSACyQlq2x9XDDegPQSX
3+KHFmWUPaxiW1OGqPP0QE54GP9gGEsklz2mfsXsyBRNBb96fSB0d5kMt/ukHKXVDqqgJMbJAg2N
GoTKHYBdZs4vQUCSdfqf4tfhVEQ+X8zxB8GJTeOIdLL/i+9++QIDs8wm8DvgHJ5hiO9fp9wlQVd+
fbemcFstUwdQx4ThY5y0H1GqW0JZpF3MBxJZNKV/j5QEdtwK9LaZKxvsDO/JjLupHApKi5v/ZU0b
fI54oJnEztx3ihAZAj4PKq/7GO70N3ILQYxsXQotGXYB7enJc+XipFzBMh7DgG6RO7v5/rCovzVR
C4Y7l6UE6DsN2za+JzfnxicAgMjYDxt05HDKRgWSzVjM6HBoxd+gy57W2996PAeoSbcXdas/K2ST
9lE6Bd5/NGxLjCoXy5OHWL/nNvKGzpRDyW5E+u0MEFslwxeILOQAFbPBZX2SzV0fOoU06T2E5B79
lfzdu/+j0ddW0c/B5V8gCJgqo7HYC539UuyIWIf//YiRRsg771GbuXtUsScRP69NBYL0KCH8bRQY
9cE8qdVAZ5fxy9hx4hYYI7TUnI2ebcumpYBBcscuRVWy0o7ToDAjQD4K2dYILcfF/6nSXSbHyACF
8qLdUOBIXIrp+z5GGGBxG2673SOSszg12sYIpze64JCULBLh68Hp5azQf1V2SkuK4VBymuSndiYa
wWpwm4PN9WJeGXE9/rLlwi+jORNltf4TyYR8cg1oGf/z/mq1YUx0FJEcWpf1fU1ZUh6qHP+GZg+/
Wg3Hy/wwVwPmJrwfsL+m2WzVCeGQ0UMOyoHZjGi5ZxiIX4LikZlfNcE78t8sxeGGanpn1diRpL6G
0y5jsW/hprotXZ1SwtVkgpmia5dLRdWt9SvIOmpNvWfIPYdHNze/mDLb+gPkbCum3oFeeP/0ngu8
BcdP5NcUPVSLg48hG0tE/a5xKdutiivYBOo6C00Dre8iqj4vp4opTzNe1b/trqvfz+3GKxkaVFXy
euB/j54v8TAF8bmazL4W4oe0JutAYciW6cLSpxLPSB/bAUHuMx19B62imOKJVMR/2m5jENTlYI03
MDq/sijk0l1pYFx52/CyaztzgDGSLw5jVC+htjJ4w1gUKQ4gGYYgdorz/6dnEC0zWaJTkp04ZbaX
KGIQx6eeWk83yT/YxCQMMuR4vYVIh9/wAJKUmMBvRRTmycrvAPb5jT5V09vqNHYG9nWZ94UktXHs
PsGVrbSQnkSfGTb6NWdtZJKcFIPLjVLIDTE25grWeUS0Eg7CGqMqu2EWgKyhyL5V0nwKItnQ+sS8
pWflC2C24O/9AZoXd7aIRYzCLCE8nu75ZOgVexEsvHZR/yIDPBQHwUy08tQbHHVqF6RwY3c/9Bdy
/8Ws4yMlvZ+rq2qxlVXL9R/zvaDKdmt7trSAoSxnIuFHKw8jhZ2dUu7LqAA18kG+bmK4eoseV4sq
+8ZY8K2Nf5fo4oD7fpfaDLhqUwcfajCQGvLJ8/QCqqSCP4I4lhQGr/SBk7s0wkWH6t3YvNCYiM5u
X9+krBJnqXEa0e2PrD39TN84Y0uFqhQdgKCnv4MUKZKhbR4LbqgOTCUylCUc6Yo+emEe4iqEsCKN
RfON3iguW46IAT6euWBQFR0H2Hh5FaQ8Wr2g/zTshkb4g3L40IEadRNREUUtreYwhVw/aot7Yaaz
mBRabbXUp0stQtH5ccpMGyc7KJUuMqYscEOuWY6y/1dvi0VafWXtjYxHEkCPCDyKmMFSefk4ko1u
MZBuhNFXirFc9inkSNFrVA+7oSs4nvQ6MIfdo2kor3k+Byti097oxCnYP+JPdCGYbOGoJPWf/Yaq
GDGYG+4GqtwnYped1w/ACao89oNR7HE6BwhSCUZi0bOLqwSqtlYfjeE/yIstOk7uudRfYx4qjT3Q
RPYNay1oPerjp36L1c1D7BBgjRx8ybMUHgqdczlRASvjl4Xptp4H22BfojsXFaWVL7rHNuPTrXYd
oxpEzkY4hJ/CAG7B9Jk6YMrIjGdThZqwT+QrKjYXDOIG9VnwLDg7c9faZxlo0dq4P9LdnpUQNo1U
YUVnkfsOi60vj4E0Gn5/J3lR7uGp3ruDFUebgzXsjLI3w1VSV4/QFHLpmg1X9fA1mSVtYBwjCtaq
2+GYG6VQAK9s9XZ79gL6F1k6T6V2Mn9Z5qDwIU0DVGWN0RSB5Q1QTnhZ3cIQcpGzt/XCRPHNV0gs
TLnwNPyndbgMFSgB64pQBL0Jq2JO4Te7uRYKMSkMKCe9Rn2KDgqPIP0kqe0p3hsIhS4JJos6x13y
x2bChEBc0xVRLCRUUJc9t9HObTueOYTJbq3D8uDZa+wlbBIJzRC8mogpaUXstmM2xJ/i2Ef5CY1+
9a2L/JJK+vST1Slsude+NF3H1WatR0pXV5sawqPi6LkN9PJr4+KwtJvShT30vY8RzvJ2i/GRaFeV
b95LhV2c4mcqvENyTxy0tEa2dhwSNdF0NKR+vnWcN7o7H6i6gNziLNHQ2sB9Q66lYhmhuoV8NiMS
JB0MYKDTS/5herFhMOmAsLFwq4q8lO4o3q+RfMclQrqJVKPRhfNSK/9Ih62cS7cetNaYplqL1O2S
sMgiEHCKJYoOEyXycuF4XQw3NHSAZhQvBfo+WW3ElJ5XCL7sp2h3gNYu3t7rTXq39Y+DInALuuQW
yJOR+BLZZB+aGz78HRpY0ZPfhufGysEpD81Xnut01DdgS12yP8YPCX4xK59dzfaxVIU7UTcWTD+C
dg5kADd71IwjoROXTD/BVvR7Af/8bCAQ52UAOQcLmfM+tr5wipAY/SFaXcRuNWR41TE4fAtQUF31
gzcXqPWd/wmfinSZgFRsCX8YQ+DAwmlPd3JxbAiGyOcC41Wo+yL3sJEhHnkRuSyOburlIW4NKk6b
lEw6dEbyx6KQIbFtCRVINdgvCZG/h3Ne3uCrEaWcZpH670DKrEoxtdCcD9+sljnKzyw3x4m/vyXm
m6yu6YHlTfIcFj4VcDSP1mex8XyrdjkaVVTmHok+s/244AnTMhLcVroigyydkOtOdITqUlbPZDdv
K16v3L+anTAkMGlllANiZvMelf2iZJU3eMfaVGeCJQpJHv+7EHxLoRX17oeBOemIGs26FsZ3Mstp
gSbKcD9X/acDdPJYUaMkM8VilgXAGtRDIX4r2dnKtxHpw+u5lfGZb0Ev+4dN95FNsujESzWEJBLR
W087C9hGhHZPGI9HUsRLiUgLZF360f3zfDIUseV3nglIX38jClQdynChrWixY7p4PZvTLJbqSQy2
04/H96C/a3NYgOXcl7DRvba7wq8qMaWKvDDjAZfP5FeO6FLvB4gLALlfPvjYl6XXW8INCPrgTv9U
OpAozWJjwJ5i13BXe5k0s3ydJvCI2Oi2kcvAc3kV+z+HYB8emrRDOfV/9JF+fKK/Ku4RsTcNYpBt
9p7cKdEYNIRJJZddKleMltjKX2m02hNanqH5MtSyT2Q0BOZg0Z+zaSGJT30prqZ3VeEyBxskcqZ9
ysxzVmFnKRtbIcm/XKK5wuTnK2NoTLwuIYMgPnr0w4qz1Ge7APrdYdPyfhpV+MVBo7DGa65TqTlm
qJe+FcFYehG/wO+20Axl84ZzuSH9w6saJ4/PM+kyqcDRYzIWbyyp+OrDS06leSY8tev7OI1w/F5t
WnZX32JW3Pc0dpIPudXjjvjQZbEtQmqasZqXbNWFprAdEiEdEuJVZ6OwVgt0RV+ACyAXIzT20ve1
76iMBzakpCdqcEzwGxBItzA1LkGeqWE3JAQxk3yhBqvP4gJd3Csc61wRAo+eJiyxYFiVNzln72OG
/yinr3eQ780vWz89UEf61VhvDRX71lFelEUFga/VfdvffnmLBo2dDh7oLtIEyPl57gOTBVKKPm1O
eQZzI9lnOTfhgqvfK1UQeoUWmLXiSwkV/1thkufZzQ3Cq8kP6GY2yVSa7JSBBhFasvVh48C3w6n2
Hnu28ggXZxUgOAmVFZ0l6qJ7bp7kpFmCqBqniF2OMMb7HdGXoGvLM2qbCdlO3GfW6NGiC9RbD1/Y
Ah3LWolBXfONjuMYd99tfocEE9t/RjGA4LqaxOdqvYxHUYhwVDFKYNNfJEJpSGXMwDEV7b6Gwzi6
DyN3fZc0Ddlhb9FsWwUm991I1mA63XPPXkU+/MLr2edM0MknwOo1+L0fUoOELSH5puvHPnk35mUn
9lnTvoWLH0Jt+mhGl7oe5K0wQD6bVlyXXakeMuHfFlpxXLuCYcgNMoXEO3yGLnWtIG8mn9NEMP4O
5FhRBrNru1mEFnvEx4zzX0Qwhca+4wUEiRqg2lJ7EPSZU2mXylZWQtqga0jnX8A+u1gpCdmE1DsV
DoMfeR7DAYekmoWy+DPolQUoWoEXU1PFHjdS8H3hMp4dL3B9xG6EnF3vHR9VKC9KpHLNhRvY/wPX
sZSYrySia5/fgQASIW8bTMLILG+4LBSt3lxNZSMXJRM3KS2JHf57RiJk4Iday2zMagBs/d/gXxDb
KFtQDVU5ALu9ummOAIP/KNjREAOMEO/Y4WkZy+USmWKkZEz6V4wVbSASOcoR/LJeQXI6Yqx/3foh
CfAdIItDghNllLm7q0GEL+ML8fZcRpdFy/kMCRUCpWTRurnyXHVKXOOUVQeB6mi6VfLODwMmpzPJ
57OLze6bs3r04ucwzKPF2bClRIGPMeaF3qSIa7o0PeoueroRY4fk3a1TP16iRQfUCSFelNfjJYI4
fCj1r61crHVrdc4RppZMuERstBSD0yyO/G0WFPqZOJDajxFySRY/XJtwKWm4riqvLA1YlbgJVBV1
8DdCzfhu9NcRoCU6/hIkiEieQlHbriRD9iHvjd4wyLmSOLu+ZIE3akVNcWyzYO6FN39BPK+QL/0D
U5/SQz0LV/72ff38HTu6YOxqXSnpM6gTLlK5ADfGGKmztT7AEYZdVumSRogvCWds6QqBCE1b52Np
K0991mK9Zrt1YooyClRT6oSVzVMY59wF3OY1Bevy6VXbiOgYWnjJMOm3ogOeCRE6LqqmOL5dVwB0
2kpnwu/S5l2SDE/51McQBhN6avWLIOAIqL679aTaBipdy1T8BuWI1eReRGl/j2WpYdwaL9LBoeZi
BeNgSobtTbiKcHr/fxoyeD4LfJC/VwgJBC51lfOOfo2d60g4oCY3i4UOJgROhOKX8FsniX5OxSnU
JjY/uDVmPptQcqEq69QTzJSZ914hD6vNA75XrcQqaMSRZNNzRge4Iu9fwfMxUQC4cGGF/QFP7g+u
7RUNzJ+OUOdROJUqIqxQ1AeQD1sJeGt8ftrsyfOJLI8e1IaniiqegD07Dg5ybqukPslQbSL4Pous
KKaZPQ6A60EDMZrjs7DokUvHYtsqYTR5DTUKMnt9wcBc3aQXm6qyXxWkKmNFgnP39UVNO5519PLW
2kjcWOai21EthIURwCyg8I0a9eupDOJD7UKqouYOly2W2+4tE8kLwWj5NkTuOrfyB9nvjKjaKpNA
G+57OYPjT9DFwAk31uG1sT5IhW15T5DKqZZFqbIGcdZHr2xTzSbZyQ4V4VSAxtnCUmiRPirtQrUJ
3WrQ+rEfuNEPXcdr+JxL5Ur9hnCoPxksYPqNS1tuPqPEj90AqyMuejEI0SKc1S+RYnJJcWF3Lpvm
pcw0foXBcmcyGfur9Zaq4cPt9knn9yqYltG4HLyyk9PIN2+dvPWX0izv6iU9ebrr47CjxJZhoPOK
+oxsUI0FGFpUmiOyVZPgdJmy9y63Ktb22qUgL0D+omh1ONwl+3/MCHjXI2covMEVYeDPGETqINLR
4smiBSAveWyNGvhSF6lA8Az8IKhPGtVqDZxV/1wCPaDzu71pVfanlFfypFlJk1/6nuNY58BxrXA0
3btqROrDaJhaqQEJ4j+lZyG+QKVJ5kosiacWD/1RhtlHXovA6lzvABA32uMiHcr7dUrsojlzoJhO
21RtwBMM6vWCFf0CbDlYacuWSJkNbwUUOpEgz0Z96/lZ7HtW3U6oBbIVJnoNUD01zEK8BUvsO7Zq
RgJt1MAr1SO6TNGuOvQdBgwBVmNtW1uNS5acPmM5R/rT4zYkLV94eZHJutEFjsl7UcgMN3ksMOxQ
pqbyodVUadA/eIhnB7D3KPj4V9A+ce2hOCUIaOw01wsPgtQWSAT9ruHn3RPDpY2x6zrtUeuvoQaY
o81SPARh48R3gH+1XDm/8eLHt43i3TRPjjL3u9uF8iz96gbgUCphJ6KxUeyNzRiD40QMrxMB97e0
5NW3iZxc+RKig+wIbMtyE5n0kTXnNb+iBVQ9h51OILojtdy/Z/fG+fUaueFA2JXNKp1jpG89CtcT
W8po2GHAs7dewedP9fgC28TpyRNNMazQzHqMBnVdpA7xN0CZArvzrTouEhtJfw4aLaSRx9VqML9d
qn99v+lXIiyESDGBvZKjYBeDFTSlLl3FZ/Q5uG908aaJw8UquNwUDcnAfrjqv913+ucbw11lAuXY
qTljjfT+yUQYxiXPohL2PEEoHKTpnFibN9vZ7t7oAF64X4Xo5dba0Zd6OW5CXGOwLhO9CbRLZAAV
oeutofW20pvxosPVjFAhVFQK78jvF9f7ZaXG7ve+bh5hqs0ccYySc4gIAeWtHB72OdDmc/fTL+Vd
t/YWAQeBdkW/aVaAeB5Y9jdN+g1/9Zg9U0wZcDh4KbTuNO8eT3ZhUAr644IOKjSZcOE3qwxNsd1Q
LMBXsBbincMPSb6iKgFg6k1ZMZ7ZY0sFwDeurCzK5aHz3IhZoN85OUP/mERXQrttJvqYKf6UaEuZ
tIK7uZQx+srKeuCAp6pJVgEOwo5JxTIMFaVWHzraP2cWZ8iVDqk7WYPHJ6duiDkXk7EaC61bDSSy
j+TdtVmuSStTAsZwJZhQeY2xqIf3Rj6YLUoDKsrj5nNXNHkvqbPZ9fBSErnQOF/J+6SHBLRytxVu
+5/3z1VxGNNmVOxV9Q9ct3uDphIc2tqbBI+szz4YIPMnGTKl738eLmVb+gpFKLDT3oWlsVCtEako
SBrcRZ/Co3ag4KXXU2OoMGQgdam2WcT+zRyKEpUrj4toUZdCoicQjsMujYPVMh+Y4x6sjasGmhFk
N5rH65fLuJKUZBUPHLFRCZiXlN5BQ+pBZRWjmBmpvWegUOgy934blE+eG+QI/GyM8FoKtum0aeEm
vHqZD4aSDoYafv6XvsmpdR/MgmwszOP4v3O3L1RFjBFVKu7N+hzkJf3D3VIQpJhc7tEAuBzPPsfy
LfxGnCU0pji6HkO0E/5bgg5hktTut6MUVTl8xSvZ5KeoebqpGirz4aoP/Hd9AgaL/mZ2NHdldPLK
4BxlbtT/cTn86AlNdSqZHc7fRJ83m6q2Weq1D2hXyXGwPLGwBZLAsplqxHdCdZ3JhgpxrC4gfepC
A4wlWNOgY7fPFvJQUyMHLpTnQzPBSvIGEVHXWV+KLDTtgOacB7L1Lbx8wa9XWaw4cNtdpatUkNtd
pPV6VbEG5xhz+4zH+dUDYc3HPJa/vdJbjnJKb768EUBW4wmz2k26teU0tF7VTvE66tzoQ2t7rwBY
g93+5WlnjN/ynJ1thRynpF5aI4GgOnIaWUy5GoD7vIcsgbLu1lslgvAhcMjR2HSHY17+1J53BBwF
FTVs6C3J7fyQYDzcMlb+V2HuzuwZiQ1PrdOCeyR27hi0OZLnIrDG0FkcAsWKDRwWofE2Ddf9Je+w
/EANJSWbCexypME3O7kRTmsOiSO8Ktl3spHzA3LN00WZQksxytVcROPZ/1eOTMHcq+G/0koO+2u+
mQsjAQ+jVVXL66cckjRYRt2QgVuoYWin8hKHpYgcv1mnW0xKF9eEAJaicFTGCdJPkHzX8q5hoPzc
Nxx5ZVSJwXOxghYeMLYuZPfoVhNurARxHNLFjrQPmEGJDxC18lMSHnz9te2qpD0VaQtVQw1PNMBQ
5eNCUWhfHR7+wjOLj8BvZ1yYVtr2g+/HxceJkQYQfpZ694kHzMebVdgr1uPzCif9F99R0+5C+gr+
tEwg9z9riK4aTs7ohw14U1unHQcOvF+oRFtkSsNxdkvyreG7nYzcapzxOYuPKmRgLyc//yQVDRCG
y6Zbzgc1NK9V/lXdHPas7K/THHEUVl0UUgGBT0ECrtF8CP9Mdzzs2OvH3ClV9efEJnXy6fYdx+JM
WaBEZ5CIGfOuI+aXMz6DiPuv78TTgHe8J/FHxaGorFaX55HleyvE5O1QSj4KprSgbnHhetb0dHGN
0L+ndXKvPjCD0jSzSykIeVQ3+ZaWI44aCWeV2xpHCCDu6l3dekz+By7/r/UZouGzTtsOzGT/dMao
E2rUTpSrNI4UyvfFrINkxTf73wkInsiTMCLdYKmm135HVVTszyAFx3gl8+esVIZeR5SFAuAnBACX
w3k/TJX0j0WXFZWjzyU2ZoHQEgX8BLizSOZRmgT34jVRGY2OOZlmJUPJ4J02xhV0Hx7r6o6735iO
H+fe5O3cMtLS6Qf5JlIV03n4lNLM6sJaJUsrNw/4BQ6nF02oHtbD5WjkN9Fac08FxKklW53WJtnc
T7MNuNHWatcyLLuouN3pz+fJBZHoR0NMEIpvjI89NSQHQxsx18K++ITZ97e6S9ixvIOVjj2bIQSr
Ecl9JWFXz22MdHpo02fnsAnxXnwlHj/cg6nkjsC1IDp/4SMSTECA9GY3/aSbsp5fAv1qETXYSvKk
RwY6/EpCc3wy/ZVSmZdbPlCrRHfOyVtX9eGzpAhYrQ/IHYWbHxoB2H1fcpI3f94gJQ43fjhcP9Sd
pV7kZFVkC+rFbq9FAl9XR+SdUBmop22SPiePcbNgiL2H+iIUtPiLZt/RQ9Gg466kbtyIhBk1s2aw
7uq/SUQal4NKI/MHE4a3eVHMljkZOlNzgxqJhqteUAgAQRzn9I5ecqKzY+NKR4x0QYW6I/v/KM6X
ETApDXBzA0Wbjb7prs9wz9PmozibjyXJE4QkScKmikt8PXU61ckYCBqCiD5EJAcaFmKRWrIMQixv
wxkSCuHPOvl31cXs+gWifeO+BTRyBqgCzMYYdb7Xz+aug/Yqp370xCVLiTBodGjC80Ec5P5OZT8n
4I7rK6sm44H+c+npjxZffGNbM51XFVL9SDcEsn5hMAAPbfhf0aA3Np6GjKI1/ft+cVhjmiNj2BZw
ZRvjWPkP89/iFokowkmiwQE6YyCSTco/l6+dqER20mwJK9qG8z1UO2fJW8nIt9oHeP9XNzjBgkou
gxe5glwwE9sueStdsIbPMDlsWdZDs+aYFgALA/Qvw80w5rB2uBiTf8ZGnMev7j6Dop+XrLXWtCmp
I0/Th2KGeO8TSTqFxxgsl6lk4jU84zEN2rnvRAhWRPSz1XW0fEV3SADQrxbnipBuakcDkAksRcN3
mhMsu9pDmzYG/JUolOgh/PG3VVH6jXY32E8B4GDr4sSibkNnXLEwjeEY/O9CcF8u36lfn6bRRhJF
0t9MVBcq5U8nsMxiI0J0SSI9KsavE/YQtY/Gx430DkXSmIR44O8AQV9rodVZatELsvJmolOKd6pe
JlMEanB4DCBX5dxfjbfdvGx+g54GHONbjce20x/uwKNak5Ot15k9uOeNSu+j15UcAjBOq6eOEsx5
wc7ZtlmP6zDXGaZRkgPUgGNo2BfIGZoFlFaUHL47lWyAwTrcy3VfdGiCJd3EmafoZzEGQtpWalmP
zKuJByFzC15YkUBM1/BmPaW5SAsX5qG2wjsgnI6MHalScnA0uP+K6CKlac5Q+wLjqQFLSM54/1FY
8l6zKqJfpRASY+Y1mVayvFWzGa1PPSAK8UxUPJPQU3CFl9sXsgXIe0twjmHwC9rJFiiu7IGHCbao
7BxbzY1JI0l+XQb2uf1XwW8gJzZZJjfXUWoFCD/KdUBdtUPQJvl27ADLREAv0bpKFme+o20AGOxh
C7TaLqq4ICK3HPZZ77ENtgTlM6n4O0KHC+o27QuCdQvcGKUaMiOiIeNNYWmkzI/BYsdYSIZxzuo/
nYjy0G8DXhIdu0aU9gao/Els+iyIw985PVEHp3BF7t0RjTKBA02g7futrpgegKGu5A5Xfx+R147m
HnPatIWBipT0oUbkgU8mhYSbURxDZVih40sRbg8nVQb97MKZnYZTHSz7+7UBuLimibGFG2LimlU0
TgRN1UKV0SI+XgGY26Yv/lpbvkr4eZI6oXA+pj37pjrHezFpu2dkxbmg/e93exFviuFDuLfpXRAy
hEP7vCosJc2chhT4Zi4FpuJTvF6RKeQIpQ0Z5JrY3yrDBBQqQ3Urt1Dg4YnEEml1+kHQ97EbqDAz
My2XdUBU30yrVp1dZCMvPYsAr0zFLnyCcW9AMtJlvQEyKHf2UWIlY7uXv6aRr6u5wcSdkjC0KXbi
F6vBl65xF5TRyho3hoY/Ks2BmbXgofn5gxT3Y1jDGf8BWCsw0xJekvAU4y6x0q8IW57tc8ntyklX
xYRviZ4q6Rpqdc03iJwEqNinm/b+FBVBXA/K3czkePjTh4joC0znOtQ6UaZFo1YaGT+v4dfsQHXy
4ed57MW3uZRoOGYNL4Ut7+QuwuMa6yfaSDntCR79ADmRi/p03ff5DUftS1aY5Tqe/X07V7AC8bLg
VDkIxaNn4HlCwlXMsC9KqV6sycLdWprPacxP7Tpo640mHoFDsdzQuFEwiQlkcTDQ+0qBbpYvWlcc
Y3w+cxjG8z2Dq4bypfNi70Va8K3b/11NMC0WJPtMPq3Nwzd3hEg30t2X3PhHSb9nYaK3YBVY8dUE
20ydCkE9Q+A1BsNLhJHCFDXE9z3kSsGY1X3ciEe+nM5CMeSaXwDVYqKwtT5sZTfDQCeu9CGiMsBg
Xp5OIPUBeGxVwB96ysAmlj+Xl8RAAJ2+lKSgq66D6LT0gufne8Y9S/MOEkN8IQiLfwoi7N2boH8F
gjotonMOUJ73NsrUsA5euzQKwnxSffmlECD0EQ5h4MDUNNVscCVDClRMOfx3o00Tlnol6xvRgnxi
koL/s7th/5RxLEp5dqrbF2OBvq29a1yGRtrw8O72TZeqniJBvAsAUvSYqsFavbkYKpxsMMjfRPfI
5p5XrLyNQmJhGa5zwvW0bk7uIP8WzBpS2Qq5tcQ+rorW2Y6uNe9cuyVhCKSpA/c3/ZIMEbxIfo0o
pXd3qs9n4pEiDeXCMvxuj6iokeU0mmNbRN9RUnwrKXjVnXHD+CCBa8woyryXfD11gRUlzrroasI/
TB4ry2x2VEu3iiQe2ihS1kT3HB1IpzRDsRvSyl0/Fz4Q2XwwHC7iUakrLzgith+R4kJRbKp0HcUc
KcaWyjf2r3hP/3njiUMdgJ9A7SRk7iIrSEmeZfDmWCge4oxmEg9DTr5Es621pRiMIJJb80Y/PVkH
M2WDXnZ8DZke/TLSa4dcfl+0FnNhwL3uhUIGn/upayZmwbT0ErCGai0qUIy0tgIcJ0saXq3vIlF/
6hB/m2SGbLyq3vASOCe3qW+yf1m8Kx3eFWv3xMa7IJzjliSQZh+GH2lStlqDQKOsB/6IPi8Ow87f
unI4n29EGU8YhOBvTZDgVC75qp1EykAPlr9+temgbfAttuobQ72WUP41ndtr7rSNTggKUMyslfT9
oUbG7GH5Bcas7ipVz2EopE+RFed3daX5X9C7VbDRgtPNteVNqJim9DXK6dOm/jmK1/RPA8CJwAY2
63FgDJnLUZ66cMFxPZc9pjoo4pt1zgB0veARZkS9HtnSDokZQesCKlJCRHyrc3yLj4pNKyHqNbx7
+7NQ7YPet/D6AKvQuhaY5mM3EFY/N2E8BrL3nSQOcgsDuARwNWcrikCxZVplMYodayIbffwePycn
7G6qEVYms7jD4MB2+CRldXEvbjx5DXQDMAgmWL4UiwIyZh45NxuLUxltTFfk+I96ELpKvSnU41NI
cC6cKMakupUqJ6nU5EXR+fCe06b1ElL5MYUtrH7/iF9zm48W7CogL/Tqe0SExBQHzEuxjWBQmrTQ
bpkMsM6ozy9dg82NdeLhBp0I346EaRrwc0Bvcd3CqpCANKHQUjUiVU0I9C/dhENTI3oj5VYPSqMb
SEVn57/KRvpRW6UtK6BSXf1nOEazGeZRVwoTHH8BMh3xgTjp93MGlbNZ81eRjK19peDo6WWwruuB
kNnD80tGiUfvu48Tkv99QqgV/FmJjcxEuZbri4NMrxkKc0bDKvFaivTXJvm2mAgDfYe4GI5gbzar
biOhi07VXHxGxmaRLtXWhGLXLPSQV2qKm8wDCucr0ZPZa/sJX0FSMfDnJVSp22nqS5Mu85aro1vz
fR8k3bKAv1n8kJFVDbxZrIp5VtdrIuxQjmLoSvAaGDgQLxxsxBgIHEDRDEHlBEreQCxcR2FYOtS8
ascGBohmIwFv3gnYuU7nclmVD6YKRfprhWrj5dtbO71rltfbvbshViHToZMa4IyCJT0fO7ku2K8z
CmxukH0FXMTf8xlKFDa0PqBvHF7JxzQB+y345mtNVULWaDHNt9mYQXwUFO2vZeBxAD7Fare3wqWq
kpp3BqAqN+Y0tXhk0RGWxg3YNJ1Jqoj+F8XXSHu0i7YwdBrdKClFsELsqHw90JYiK/pykf2V2CjS
LrrbommPjQOAdrG1xdeMKb2RrgYOifii+ht85cOrxx+NHtrNqvFOQNpe7ZHaeCBUrxOi5Mep17U0
D1YwoG75SMzMYruV/G35PJLUmuaV6XRwMPSg3VP4j+/Otoks7Wi2Xny3I2zx5p3iq13UdTFJmomi
jbvs9gqM42DGrUEsAE80SicO4Kt+J86Wbox4whSofgqRc71OC8aIpOwqd4EYc3f4XZfWsJJktpTl
Q/jiRmRMdki1bwF21Gj1lPxMzwy5DKx9lMW9Afh3FC9JxjqjGK3Z3OgpHJSh9x0JjPHU8U32YpjU
TpHpwfwUNUB2Yn/235k4L4eaPuqIEoex95b3LM+cSxPFZi/ivJoVByMocBBmpVXeJUwFhG5Il277
d5TZfH99ZmhRAHPn49/KIku1NxnHQ1RCHbibllRFGfRl92LY9SZWNPWtubM3oP5g4xaU5O/vCEXu
ZGwVmbGzgjek+Y0WOQUOAsEnyQota/3GsYXUsJ01RHaTGc1J6hkW381/+eewcrL/+xNREwpPTjec
BUcFGe0aWM6j9hijVf7opN5rNnUEIdlq7pEfdBteBSjWiDeTuTkZlcu5Ty//7ssi1YsROpR3Vt3C
INWL7ehulM8QU/+nbz2QRqNvvOobQIfRh8SP61d7Bcn9nHSj9UW0sugyqyTqjS966a8z35qzAfG/
VP6LmbdfF0NCNeRX6aXhW5xyANGEq3KWu6Jji7VgMAhHkPTO8Qjh4YzTrrnXXAXLQuWUjjzZN0qG
93lYUq2ig9Gqgq9cG+mBxaHSDoaBcXQ95VSNT4Kim+bOx+vh6Lgw49S+TiyHwFgTD3w/htAfOeJ0
HwbB9Ll/fFj92BElyNvnxEmCIfKWZ89WNXLUJ0xwJ/1XuOhVSppAGACz2SG0HFGudY7MW0OXy8sK
wi7h98UD6vlzlU4w5Ip9gpen3/FKkt7xMb2TDCf1iyEJ66hGIIbN6thhVcsjra8YNIEQ8GVaCO3I
5bgIb5QNbmT+lYuvDy9tkoja16Jt5IZP8n5pWlb64GKu1znJJEvYfvQRssesvz7xjzS3kBoMhUCz
pNCB9x/mj7FvjXz3OZVStATEYeSNQ1l56EwNs1O2kTqEfqvFqAfzlFV1/FYyMMekweSw5KK7KnnC
zpPcE1Z4ieEzSwP+DtFyfuEK0uj4pvhKd/0vP5sgEBWnMJhbi+meuEMq9niiV/x+xPN5jtYGchHa
j/UqKZB2pZab7Vu+zivGjHHw6BaCBFN9m2RWTnWSSCpzcZsusqBpefpXb2kY+I4B0OR+UcjHJ4cR
5wgBkQxMy7xhn1e40iKBj4ZnqRQ6UVrjRWFNlFEqLL530oRoqZm7zHlaA/XD8p8CLtzcDsYBWLq0
lNjxxa084GA1cUPummS1XMvK4jk7KLWSsh4ZED+XyWjFgx3myBmFWj3g3ZOIlTnfjLiFFZPGmfc1
Kt41GKhT37xyC7HBRDBTVkolxS1b0JXP931yrQWVQqriCkGsMqkw8h3lid+de86FWAMhwcE7QwBE
dzztAs306qvHHiYsIxF+J8cfA3VfPzZZzrA39mll6S1s3I5fq61f9zwSRtlyohMvbY3Df3GbV+Ut
uJ8N2hcggC6LE2BrnYi7hl/bLzGkg9EONBZl7L56qX5e1HFudekI7r9I7g+TtOmOSMkM1w0gKPM4
uEL099rYNJN4qrlYsOYOIzob7qTpZnquT3oMllCMrr1Va0Tr4BlE69IOwju/cquENHSDZjaJ24aI
nogivgt2wYgf5Zb9c2HfIhoyf4/wWrt5Xs4G1PuyKS5awoIXOk4ee7dD99A7oiIzc+mIvIrt6LxM
3UOX+0Slt7a1IMW9QnxZiJkdrTbup6hcjzmR2hQywC8/+cBqmVBV/vJFstIpmuYd+NHqqTrr4V6b
a25HZowaqdw0rY/WmZjGaaHB34FrT9BHm3UQ4xDk0iKjzXDYEOi17x6pDb4gE81grAdhU1HsfOEl
iLWWtHCO3PYzQdM2X5HFQ7/nK0zu7P7HRSl1ur3ncA8+UyS08xp933kUCzHzS0Iw1353xaZztVov
1eBdNNl5lx5YQxjhqPybH2kh70w8DrzQLasLrahp+wupFGdUKI+9EFE0zQJi/AozVPM1VeLXXhWi
9Nga5AEMBjGn5z0OukfqNY6j9C+2ED9AbwFeSryW3roWq7MVAYuZ4IuumS2BRbpUOnfsF6wKb2+q
tDqJQofb+bZOrcZQDJAzVxsOMFnc6U44bX0s8gCqVnjsKHJZUgjmvGOhr59kJTO522Z+lD3itWH7
hLsFZv8csTkoB5ZzrEhWwr9G9RaLP3fAgPNJgd6hMIGmIanx/tHrZElN48KDIEnfTcRoLjqQEAKK
fvt29T4/MiOuMMXZodzmlD9M4sbFt+uixnsx8720DJsOr2uGOs9+W+KvkWSWg7Oc2fU2QJKeFV8q
85wCd40TXUvO6n7Ktwi5yLZOz+hr5hLLgrZqPe4zkkoHKtH6WkXksw1jA0Wh4yZVf84ycSvgRxxI
LDg4bE6Ld4Q1LZaVsumJcJfuOCDX2K44nF0SZ7bQ5P7VvhXKZ4e6i3FlcUF98Hh1vUWo//IEhnYQ
SFWXRmXzG732s8zgaecfhoc65U3JUhDci6T2DuDiqg/tia6wp0UklpmtNkZKTyKeiAO2NGrm9TYU
W9dG8a7jpMCjhhldXEWQHpH2eOdHWRsEMgbEmWgcOog4KKNnQ1wG3HOmeZ2dfwGk/1oBIz1/ai1k
JDwQIn34D5S5nue4K99TD3E7PhjNIDCFpQ0RZJvyMLkEPROc1nuRcNU64NZUNnc3Tx3IXxxrMHKK
f7zGRdew1ojhQkoVWUyWfI6Hfy1cMs2vZLnPfoAsGJWr5GzBTTGrUIu6OhtTMQJcGFxaq6N8Wo0S
/1nvI2+QZxtZoRz1+5Y5ty+NWNxM6XGetCK6rW84Mp3lx8Rn0OLDBbzVYqH8Xwhta2XTYvyoybJA
qjCaF30w+WeWtOlwCFS3jyaZFRT3KTnZNQ74+KylzFeSKzWra38z0/HpqefA3oCj1U2gtPSUCGzy
RM3leXkj83l42SicOCw8Sex3asiBqm0v/ESgJvwSUJelqUeFOfmdyOQVOnhAo8gqqvpOkEOS9Qrw
sHYn8WmYP1FkS52hUprOX4xbE15gJfEMSUDnIkGxgxlHYkqls4VQl9T4l7eS2GVYqmCGzKbfkQrD
W+SW3+eve+mWh+L8+PLY8tTWmsJyn7SVhdwtiBQECd9aCfhiqBgFX2+8lxBqB60yuOduphuXUTim
/FBNjS5xHWkiBMp09o+7wbY89Flee/WxhEmdk/4dbzNuMWrW9Tiuyq7Px0Q+78DGVQUgOuwwVVzR
WH/OhcziQLr/DJy8MtREX9LHOhvxnsoNDXN1zsZD7hGlEcxSfGKKx3s2Iw1k+SDt5ZYlzaF4SFby
xQg0Qy7HbYGMMxypAhAO8IhbvfyCT40SZst+dy6tlZ+8uvSP4O4o4qYKhzjFYfzcRODEyMmA+LRn
lSWOhnFQphkeg45SpZommpOmruXnsiTmPo4SS0NWFd6+sTKyEgmg00fMbqmoa2ceI/MKTjQhwt//
Gm7WWChD+LmFIJmmGyNZqgH4WZP6mr7Zp8BFNRRvqVJZOZuJ8InvYcTXtd7+7UJtifoLkHzaQLEY
D9ine0sn+7naSctumVcIBs+8xUvNq3p1gsfca7kQZuXo1obPRCJA4YsCjUuq7uQFOsTLwebP4KHS
tkKog4o5uydDQGSXmiBfp62PAFmC7kMKMw552VQmt5Wghrml7dLaU9S6jxKRd7+GueKZhgnLa3m+
n/32l0YOjRl+61r9Xlf0qgxevdjqelJpZO2fwufb0o/fgU3RrnM8sCl2HOFzo6HGaAElThTEjghC
Vxg03Fgld8yt0RPM8ApXWNP/2uzpHpnLNYK579oD2Fxrx80xAX0mfTYXH27/QbuJC+n76orwHQQ+
W3u1US/+OyJdk118puF+EwpM7GJlXUzW5pt40tc7N5KVGYhNn5GcxL3vPMhiJBBBfwPuO8HXmM3B
s0mY4lIxkwWdzt+YYuKoBT8Lzj1KGtnuTHq0Mxnv4LDsQWfRBvuSYq4fRPn4cJSDxzbsFcHbD9Vt
ouQAyV/X28uMdq2ntYEc8mtC28zDam8c4K3OE87vMSheRbY/dT9Z8o3TUP+yo+R80PiccIPBAM7D
V2Lj0YOLXSKbJfPU/XXEFHneRfSFlIz8cBNxhtCF1m8aHqoG5UU4Cun8KSJ9OQA1mLHW0iC9UBky
wc062SmORyrys0dJ4d63cqg0AlpLSdD12SM/aqmSaty93yEv8ICftz6Kq707zE2lX6OPIydvp/VJ
EYoz24YEFC44WCUf3xjZYozZ1EMp+dGbU23DcJOsEKWVE1Oh/OMNVgqpJ5jw0APEmTT8ibbULEP0
xioQHELAsFFzeN6PtyxAzEcPXAtCRdlNRHfAcWMzxZ9Qp/NW3GoI1TJlEHieqJl46AKyGmGqx22c
JohHh9sFBuWBg55vfP3vPD/FwQBLTaosjKyZhoAcXAJ97dSY+E/MTQLJH7epdeH5X4ZNkuMNyXUh
41vdMHvlzt0l/qIWnf4BlmMR+vtoUFjNY7kdKRolduA7MM1dU6KDlQj5bS0amadVcqNXW1Kka09J
7LeEX8AaijK0hmgfuMusn9iALyYqCuQ7CHuG6+mzBl+p+n7mzXkGDR3wJYREIvj/znk9IKFrE8R0
hcOhh29jbEMihlGtTTRjv+y/II20SlbyjcAbBXOZejlpRbjxwdF719u65T/Fe5AZ2nt/7u4uwCj/
MHcWeiN1Bg0+JQ8jPuDKxzk/4LjZGNg07RDIUhtsic5BF7KEFqSmVglHibDLHLjm1GuYKp3ecR8J
eRcHJoE+c9p9ydxBNHSGrqEVrnP6n87p/SqcZvOU0WjWy9HkTvhqiE3gZ6WenuCm1wg32BsYHrkj
IS8i4NqFNIs9YWuzAELACZfR/dxLawEOmxW/G/JXHEOJWX7XyyXh00FRs1kesa9aG0/i3cNnJHFd
vbUWuZOCxAOHZXgN9tDJ5FeMQA4o/fDt1sQvgtmtZPt/wX8f3HWAJ3B/zXpjzeOFjkPxtPTrhHDL
HvpNgA5ONJhTxW50rGXze53nQG5r98yyConqOcfjiTHePF8JzQHfQrKxwI872atV0tpEH6pIU6bp
nGIiaw/Q5MgZP2tuuA8spNUkAMSYgp75iaNDg2iiRHrvlXytZDetGHHYaZfHD8/VxWRySRg2vZTN
30qoVxK4xxu/Txq5mrNT8E8jd1/RX+Mne8FNkB5T4algtejSkYKLNnTLX0AJ3jnRoKnHPrcs12fP
L4gU6z33yGq5sV+2XkSCQ0e2zrpklNAPsJ5BXOEx/2X1BFzPG49bIGfHdfE4FTe8ghQYthT/X0PG
Wodbq1NjLb65KMjLrH/GTiewu4y7g/wcGV8X2BZXdFvaVzmeuboAI4iBY6s606H3M6gsRIzT+qu3
+zjXHDjg3HYzr/Cvqi2XPoLQk0RLBWPmMDFv+5RGJobVD/nW8jKGMKBevLiqzykpQwTgp9N5CSLM
yDmE5jE0Z0oQsi5l+6rE3lqy8lkncV5J/p5d1tzuKHSRA5tWs8QXcvcwj5zgQnFpd7UBWKHcLugd
FDtr4L4TWJOSczomGPpvt8Jbh4y11YVg/ZYVL/cuHDpGiP9e5Z0+YkRCWs1ZAPMDsZ6qSQwEfH4g
ESfDxS25n9dERUGB9yYHXHNdz7bCx3QbQOQQPglvYYLPBb7nppCsDCC/DJYFf3EJ9c7TUMq0kEfC
3EZlPqbbfOYhZfrI7E9VQNtB94TYm45w4LFHLy3roGzuDPGkTy3wSeVZp0DRqH84tb6E+LoBh9tk
uCzOtP0wfAGyjvYjvwGTnQxftfsofY6BYle93ntJ7iJRGBCCmB0XtmWc7fXZr9zfuAwJsn9ZtmrK
GfBd+FM27W+uSWwMqi9BOiWjMdQMy9+5ka/x6m+qUBPbGIoIOIX/V4hlRiAQ4+n9QM51BQ2RI8xh
YiLYrc9YOzzP0CXuCn1E25BCIWpVfUPxzDJaKlcdXv5nBFs9H8XIwD1bzIpkUf/HPu2GdpT2tann
hmc3jf/T45hO8qJXZYPkd3/ATFExsjeXiHeFWQiLan7kKGcg/nj27O0V1UPk/IGLihvpmZk/CtPR
WPtMh3A6LibTRbTXwyTeEq7nGqZX6av+51gskwucGcByL7ncq/uIh8/agBBQ1GMLpMRYMeFHqId+
hMV7TMiOwYI3mM/Se3VT28eiLnNrG7uGt+QIOiOxR5e5LgkdRJXTQGYo8ECgkNkeBG1wg6smDKLw
LR/H/99gj379/QLZVfZ5ieeTxaX/p6MU3QPAfEq9xVoMmSs/AH87bLo3t1QReqokpt61GBVbxz4F
D3bXJPs/1qD0m8GTQkkkXAnHEllfdJibZpsbQo3MQvmvXvFAiobuPKIsVJeHAFnRvrPhEp39vu8H
8Df3omR4e9XFHsjkeal6Gpn8XLei50/qiqfwHk9HJXCcBPaOeWS0LSpXCqrY6olzOACmgdB3Ovt6
K3YWt2Z2J4H8rplNzYdDmB0doxt8TnGkrEDXGK+crwsMSLsRf75XqvlUv0j7JaDpvbdobc7tBE5n
muoxXNi98bH/SpA2cQ/KnmpuunMxFBWAA1OKvjEsNQEN7rao5anb1IYuhtLKVyWtDFIyN0ldW/Bi
pPllMFWqaZIsWgXSOCgey+IyizqHD0qT5+0SmbsS+GPEdsluSJDD6EJwOxv4blR294iXN9hOAqcR
WeItmHtmPtohANmdjz09l/BJkrjxpJicehqAUBaNqa9o4+meD1gXEc792MLuY6MtA0nTIZ4pabwu
L7d003UoosGyk5xHvRFFPov43HADmcV/GaKOST7njH/IMKI83LPVVxsosPEFfTYCFScnemPHPVBD
3BbjccjiCH2aklb/UJXA8VARl9vYHJUJqeM0fAw3Hf13kSoQk9GdQGDqXw3ZhOMNzDr4q8aeTwPX
g+ZOSvzpJJc6u8tiommp3sTQxlKNbeWrEhh7BPxjzeXJz8VhnqC7rsQzDax4egcZ3Wvuecrfx0b4
f58xg/oNhzN9Pfi7ZAi86tQa96RlpgFy+xU260aA18iHTZg5cybzaP35Ax7kv/9mF6fUBHCipf31
c/KpLduaJ7ly7ZJ3vGadL39NZWH3O4OdaPuGMP205zeNSB5+vXb6yrcm6G1Ke8gbZfdBeQN1QJ3p
eK+YgjMITVL2avHCl2TmvI+6c6qGuJ+887aT1C6PGKvgLumTeNVk5Jy6F/e1F2PgZbi3LkkBoc/B
GQbMADJG/IKiQcfVc193R/LJdzKeHA8CB1oDvO+f5qPTtYve6NMrIqAj9oIlePCvBNCGEPVaDAfW
l/zv1rckj8cwldpUjQIhxisQyy6meVSPu/i7o4m07qshf5irbuDUPrm9lCJraBfQK5iYNrr5Ta9f
7HnE569fsr/DWFJGm6D/ziy3Q/iEHtof9cesGfVLzTkuhFVH5d//ztLpaq9peVU/uhL0gDLznnjI
XFeKd1OvWueWS09tiw8EkXt1GEUgzlgsP8zxclqxKUzAkuhNor3fj8OYrUIdmtR98UA1ff+gVS1+
Q+kRZJcp67zfYBGV0D9o+JjZtBn4+GfI87dCp+P9JZT0Lzhx2W4/d6UtcwRpSQ6VGQymlvuTRsao
zKS3SKR9C9YhzX1MxOs/V5Ij9l/oS0V0Ftjn2KdcbdGorJ7ARW/o8jlp3BUJ8VT7N1Bxb0DXI8Jd
WiQPMdpLQ0hDgk9rZN7H38Mx67zEO+q3qVS+i22E24ZF6YFRCcZPKEQ8jzTb7FVh2wkckUmEjB6J
zWL+i/OozxWJYkqei9tuCRiXPH6FLr9eJEff4rQusy1hzIboD48i4WKjeWKzVywaoaDeYoru/L9i
75pMrDGCu1wWhdz3nG7LMqfeUIOq1siZWhtyvtOP4VoDOuhUOHQZh4VVaYISvyZvtnVd4k6GRHDs
emb/Qldv3bY138EtrTNbeGHW2h9BQC8IKK7PlRIQfVhBxMY18fA8UkabOVW3oXvQfUhMPAg2/jwT
H9NZfwklIoVO/hcf+kQSvhFZyx+PYxwnTd3Mt/l/lMGl8vtPGaYhUChtcE4C5HapWrMGRfbGGnuY
5q+fZFRyfCIp66cPZ/k5iCkQYwHCWHI+bl5aqeKgbMrz8YfvjaoA7GT7hoYHn0wvkss+WScF8X7C
VjEDCpt+VU/r/rS2EJRiRHm/kqsHHQT0F5RnY0fUR+i7lAqV1RyoowmZYOZ1LYyZaatzDl69wu4J
NvYe07iKdGeckiWt8mf5EEE4/zFDBLcCFTvSUb/doSy4dbLl3DoWjOFUePAceNOzp9xghP6A8dyY
mIivWLw6QdKnh1UiUnvl4ZdCkmV65t9qPoiJzN1mGcpXnJDlw2fjNGyePHDne8rL3yo2tD9KtzWc
ataxwp7aLTfnjm39w1FRXQBX2hRPdXCqMbMfI+kDdIRCYxEjzL2naMfSJMBlFEcGjGNL84q1xVx9
lLRB/I20Syw8TpVIRWZco5yLTnb5cM6yJh+ERdCWWo0mRZMWqG4jh6TP/HcNuE5KqpobNlfqYv83
0+tEVDk1TFkq45DDDOe3V9t7K5Gam6ycciuyG4kU9GjM3aRepOkdZccFp5hqi72bfwMCzcADMjRM
+Dzjragqr4BU/5cqZH3FcEz5WqpPOgU66HZnB9lXmvPLw2R5qPgpY4B68uEJOrxKS8XUMeljh6G9
2yyOuhCkobIUY7DNk0Gxd7ldG3JWfP9Ymki2AzF4XthO5ePmQIFJFDsK20onatHpdXK9OaTRwzGj
R7b4w8PS2xZ/8B1R2cEQKSvqFKW1j8P/Cem7nVn8B6pHHuR2ta5RxPvg/5ab/zC3T41svjGOkwr+
CNBj0ZrktJXkSIngXVageZdjevV7W2d4PjE1X7XdylwXEd+mLlNoMcpf9I0lSqK0p+GPBvOtocie
WTj+ypMaBJfimpHcKD98jA5O1X4wnsgKuq6hk1gUvSeCLRAf7rdKJuOEaYV3LVaNhvH0p4hz1z5q
ZzIRtHBcwRZqkioQS1xOASuynIGDvbfJ+rp0wrcSuAsflp5uNmKRMNAlvCklz4hF+XMntEfPWEqs
kJMRGxn7vW3tUOLaXP7k1PM4n+Gc8+Kq1BDiHUb1zmX0FmcjJLgt8K9gfWcxFL8w7Fv5C7Py0FIf
k7aIJxRU8o8CNeLtpo7EXDLT0bwO6slf8xZ5NC0ONIQTVzxdqn4kwMp0QUMmHa1X8xTQGKf3jMgo
n1YAzcruO90Fsq/+Qq9KjPeuQE7Op2NHzfi9MRQnIy26+iPOtvCP6TCaFi+eVtGWH040qQ+e57i9
axV/Pp/4Rn0a41p3/6UHmkSMtVoC5rHyMuh7NHJzyJcoBo8EsVwWg7gAMHR+vd9SAXl+l0lYCYq8
/F+JkSPvrdmLReWrunRWm9mpDVPVW9PwlzGzfKQABua9DFoCQDuPuH6w7gyttIyJB3FdgiJ8BJ2k
ObafDBpRAtU1OohndwDLzdZHni6GFzPJU+n0Ndou+wRrppJk1wxo+1jvUt4jn5OaL9cpc9tteVOO
OI2pme4GY8wZa3uu0kKiR7pMjO8qZSH+3ot1wtcLHLbBdz01m4NdsSSeMXSdcQU0wGngauCWlupr
fyQFi39TSSxKaeFpJFkkfHwcaNj0ruqf+d2uy6U1FykwTCMSK5S+0mL6S66x4Nt3AEKUL1ceuqS4
0ewSEEbQE1R9DsvVCGaFM4A3uQ/Ydt3QggaR6Phs0ixa9S28MEmNTuIMWOJVAnd7rAgO/GKouG3l
4nj4qdeM94aitPMeVq1R3mSauJGSI/MpFgcz1MJ5GBmxPe0iGmTQyedPLGFHbnB2o6Y9rtEM5sly
fZAwUiD4CugwCV3uX3fp0S1QDKncawSpNWm/GxVkvLp6ltKgU6tQopE4JydF9eGukS6UYKdh//Ni
nj3G6Dw/QaxtvDdusGtr+EMvD+0YZ3vXqN9aSL7yO7WUSdAwoWAseQzIGKqpwax3K3PCXF1YcUiu
pBvhIUi41DMLKHFIMx9LjVuggUHc1AmaNIMZfRAgMbIAp0/rtkFRLkWYOPEH31NDu0Ln3knSwscJ
1vizF7cNq+HYxD2sHkOWIaHU2xUxrctffTQWqzNvu0ElHeD6JgxTlNQerOCGrynXZ9t1pgeC2Lm/
k3K7F/Nvdie14o/D772M+odcgCdWsy3o5wS/1AtPDKd+d480PUNJu/JSZy4Lsqi7LKOi2GYMxHWE
3TQrVnk7oPpgOAuB7tKuBWlhrm7BAq65lrX3oDytj0Cy+wPBUw/6QMoBRbHUwwVrxibguYu4Sfly
bzqXeoA++PkWxUII8JUw6gZqRhfIVHJBVv1Z5PdojwZi077vvnEljZxoihoB2EPUyeGbKmr+YohL
XBTCMQ0LN6riT9vAwLo5yITqt+YZqms2NKG1FcXyugrWdoTILfhLZP683Q337PsUcJuN+lZyTTdL
V33ZvV+mjQ1ikawuFaUZjGE1UA0tgvMbNvNsVo38cdv7fe0Hl4VxKcdKPejBdmQHPUppBZXo14bE
ioBfl5ZIbDpFntJBlhEzB5E4Pg4mUsJ3qGxpAfWT3dNBEaosoROItxbCs9UNO1x5+hhZIy2zQKc6
mkjdNGypwBOMgqmKQu1AUI+RCGK7rx56CXstj6GN7C2y7+WnVWG6R9ScdYo/JbqPBdX/n4Dt3fZq
b6pSHQSAtMFmsN/8MHX96Weo+SSoXn1P3lw56FLrGfmAeYPwMmsddhtru2EEDBxmKNOaMyvpcCPy
r6IsrG6/xtRcl4oyZddoPO7RoN/JAda4rEgJ80kWasaulv59oGG6bCb8mgWIMDe9IXyyM0c9CYgz
cP19jjf2mbUl2LAKmCNPvNp4tJh3xZ2UP6D/syLLRlkbCEOJ8F/d76PeiwUmlM0brdMLmPaL4k9p
p3wdJnJjMazOsi00p1IAZr3+hMMYxp4ONLs4QXBFIW3e0KYsiQO91PsyVrqxk0AdWFOKsAavq8C4
pvjDcvY/2kz/aACGU/cMRlTY40yELyug2kovpUlG8FGhGx73jPPb0434Q5PsF0gUeKja9g9FEbgM
sW+zbT7R71PpSMFYuyBBdvlUf5XKfGOUyKErITBrl+1GPOLGMnevrlATT4J3YPNc7Iz2vpgacmGe
5n5ytFvfmG1DPG7URC2XyCoRER1mv+yx2Rg7p2gYRy1R48DtT/BYmuVCg8QKklotklajkB9GPlcj
hcEuyePNNTB6N1oaXIsQvZsQYaSmaGZHS1GNJ8i92IrohQxz4MDEmhWB3TJQptzdX6tJxxz2F2Dt
H/tLPBZT2AV87RFXVVtl4MQEFmM4aL3w6nHBA0gcMPBH1av4F8iz0gC3tefdqcK10GtDpxsU//HC
KnhiXfgpsxESoSOojbJgVdEfBxI9yb1zWLrVDT140QqObCNfBOOjgTV55ZtV0fWtjc1MHHYv6aJC
VQ2zXYzq537Gf9B9SuBZYRmAP+Qss+ZXtcLiUMhrFx9zFw1QGXSORBAyYUqYBDaX0zeg7cYmBPFN
GeKecpBa7S3bDh7Qw8mt6hdZ110oTxBRSyTqKAJCvHZicmgfZqb2+IPxtStVDOIY3FOWVeZq8gd+
77CkTfmDkOMb5rXrvmuvZ/HQa4F89pnMQ/rfmTFvTXmcEnnnFSjqqzc4sRu7KwUiTYSSly5UpA+/
FhVVBCN9Pe65yOFl96morboZ68qAc11NZSoG71kAGP4B9daozWTwY0dXi8o0QcrzAw9iqb4KD44/
ObjAMzzaKTWvERLUSgSeQ6wDWxxDanFcKapfnF3p7a8C67k0d2BB12azonWpoP5vP4OncDpWf2Pl
xRU/dEQbdNjkhjbpzlrWpFHDa/yZOKfSw6e4rGxduOScFlRTM+jbkiAvuASLK/tQsM8ArXfesgG3
7bmwWo7BVmD85kXUxFyt/Rm2UkaZ7OdVn9SWJd3frXz1T4SC+MC6HZzpxoOp1SRqmu9X8QFUuacb
NHyEOpEA3HBKJeGt5AKIYfNUcEoK8ZXxtbvN+Dl65tN85tu1Sccz17Elqbj2cfklRMFjWakNH3BG
4DxUvmjQmiOARNwV8kF7h7O47sL0HmVqTgxDTaqQSVZlLpbzdkgONddvuo64kwcheCr2a2LT+43W
+wjETyyzPOxy8bGtMU1FK0rtHETxikbXd5Df2QF6wtk8y8bch20+qXTz1HXK1Sl/WIQ0Zp0BRTK5
lqNwdlhZ6O7SRlYuJxxt87Qv6DQSNxTN5gfiiym6R3lzbe0LyHwxyhEt82jIbOXTake3iJ7YStNI
iil/twdKowLf16UPsP6A93Ol/0oCehEyrVG9m9i7mZdfAEY5VRJqJDzgx8vHpMjNP2V/B+t2JU+N
PMG/Io0SIPHfqnO9HOnS1ZysDOORsA3lMJsfX+/dRf7TFAZk0Yxhvqy6+s2gNtlKYMm7lZqfmrwU
YzKvDacmzTB820ioolsELGYJfQRU1/30Cj2XQitXF7ElBZvR7XMSxXzd0thHAjFsY63JHqjfrKEt
Snza1s5VHI2kpYGtwGUeavTkyWo0uE6cwLTovGNoIru6jUR/FxPUjuqq5HMklJLCT6U87aruYdrG
ZWenRCg7MGiN6H6u2skGDBf6OaBx/GZ5iRBsSMNSogNVro2cKcLHWiy5+8Pyo030vDy39Wn49poH
6dT7B8crPGWKNMv7pfZ5IFUB5+R7P30pCnAZQ6C4VadGUXxDvpTB0beSWlon8Qtv7BxlcnvM7TN1
6VHT7YJdm7Y0pUuBIhYWNMmFZSjhw1pJo4D9FY2q+Qsrz19k/xHj34wsa/9v6GpbLSyIzAohSIvM
i/iuQakiuGvX8Z4DjxM2H8fPA0s3ZjpGhTuNKW9Zwqg6PEnoU4EHzGqhnjs5jC6sgyqMqOfLMvuR
+D1bWfXZZz3aahTJDuhhNDB/mCYqAJ902CC9vIV54GPN+QBrGrpzc4RuKGMZhqSDoZOKj96bT0US
nSLbT/zsdcgr54Pj39YKd+Zfr+N5TDM1S9oovSXaZCdAG9DDyX2gREkhmFDYg9Ontft0OAIor82S
iPVD6h15agJiYn1bKiGpeY+Eh15wlf51TiDpg2YCrtQItlZg8tQYAMqqsLtjQ8m40RzbdA6o9IHC
VQEBKl7xYd2LFNx/l8Gye/On2rxyGP7xw8EqbFIorBGVrnl8JPptUBng4GmJfCWVJmkMcZCdUbvP
wkzqNCHBKLPxJ/kfW8FcstthNEcvt3SmtdBJM021DVO5TwjWsXQhAFNA9HbyKeGOp9+PYTCf1q9m
p4xz7kdKhKA0LmglR6QM3LLCmgkYdCWnJk4Cbr7IKDY1+p79caO8p9B2ryHvQ0xmf4H4Vf1HLoOJ
Dj59yOBYI6Tas4a0OOegC3ooGBLPcE54Q88erV4ayZs1j5S/XlHWVYGYO3qoJfB5nDzyQlCqLV98
DWIEU2o/ptSI2RTYdSvveDm2OJtXRNMprpUxR0uBTFreTRQVkkCT5IvUAL4eLMw7a9BwzS4fYIpJ
KXStP6RdG3bblIvlchp7ntCRoXGAcyZcCRSe3ITsfQwvff5vA978rASwuTNG7VO8M7Oc/fLwUf0/
twGVBIT9een5dimB81PfFmj9rMK8IQG60wYw21QO0K98sqTR+DYn/KOoSBFGdmqpWqXnToq6qZs5
LU9yK4FuLSrJrmwpGy6BcgPbwUT2G1P2RRRuw2ChXY6RLs5hvA717rqIsTgfI68NLhh4JNp+nLRa
8A9Il3MIKsSz06LmAv0azf989qjE+3i0Fld9OEMtuMmfbjJ18XsMMuSBRAaxvtKR73yzsOJcp203
zLwhEceyOwmqJ55FwIrRtLd8TdN1Yz2nu7UTspZN6jzc6NuAo9ypydJVDN6eCSX681kt4c8TXmRx
bp0F97FrAOlSm1U6M10Yoj3yFj0mn3VKqn71/exVumT3mHhB2f/r8DKC2gsYGRr7xUb9Q1AJN/BL
7WIoA5jbtg/LBeKc03kIvRm0+qDqxtAAiP7V5xFmLqbYkwj0DJdiHEi6m6L2DXVupEDd3a/kaMFw
R4/tfiS5fU5Kl/zIERLviSyit72s+9K7o0r1+reTdCsnjnxTFIWwSojYQ2Xj5dBu3BHVMrfZPRSs
0uBzKYWUQxmksI54fzOHTizGTu1UIkNcorQTQE09xJR6LpO/PtWycaAXz+uSLpbLHGoPz14AoS6v
a0Ztg1m/OymLOiWxB7niCZd/QVn52p9nf7+R/2FGROQ9yKPhCFEEWiueTJq97MVx9/QX0zbovt/T
Gi0leBCBzXEPcMagHLuYxVkpSnv4ei9XbBO1/nUqhvlm8nkv37eoVcjA9qzTMmIN8ulxqhzTmucf
RwGvaLoXmhVpkKSYxIBSKOb7VonlB8V5BwcpOsTVvxwo8Z/fd941+UDsRY0WeeR7P90YWgIdC5hJ
UHnxxNvckQP7DPd3njr+2vKO5U5Xl8N9J7PrFeeaZFjJ4RTE1I/8olcYAoyi+msvSxaKaymYDGSr
/tEN3jdd8LhgwqrRU5V2FLrGRvcftC4EHaRCB0CNC/HtUC0zLfO/PJ9et7gzi9xi1Maf8WprdKNK
xbgE7i/eq7nLOJcDWHwJ9/iyeIBWALb3nyZM8E+PzZe1ExAtORhCxXn3bItHNF7Wk4QsVS29zmyo
PpBwogtQDxhQYcv90DUjnDru+o/GRP08dTXJ+L/BBiAMKieYQ2/XmQ0gU6G0CxYBOJclnIU/mIzo
JgarhQJ4J6xuM8vidVMbW1BuvZ4FycfvesPh1UKTnGoMSiU6RxXZTe5dPg3dB9QHMentHLH8C+5g
2b55wKUkKP9RvqFavGbxpgKTN4eG22TSuxt3JkDq/wnmXRFgGdkZfu4e0YfJeeit/14xqs1uyphC
3R2NmKBPXlXBMbtsA2zEnNSMAXtHuUt4mLhajWT3/m74/jXSA3BYxU1TLWIFuTNoCc7i7x8JZuh6
W6iuIRHx46RhkRHii+8uzy+iu6Z5yREaSBI8mY28fOQsIkhERwYjtVOrlx/7XLvDudukQ8AmF1Lm
FjH19MVJfs5fTsL4nvXaBic8Jiu4zykmpedEtKGqrwzAm9xNHAW1W8mDjSXRc18Orhl/XczwSk3d
mEYx7JkMBjZNAQUsmLGX8f9M/X5HNl2hGCsPoNBb5FQXzA9P2MD7tMwG9cE9ZuxkBUAPfFmqjM5A
6gPZbGUjSDLi0HnQs0B2Kp0DSqvT7h0yy5o1OGLMUjVnE6+SniDdN3sSudzj/rIl3RJek9j87GIV
pLjjnMKMH82OY1OOeK9ctXHA6xfOGNU2Q+age6fghJcFkM/DsyiefGVWupBCP1vPtp/oAaVuFbP/
Vd4rHrLIBKhY1sT/aZeqkw3AVEhe9mDu5hFJhoaimqJC6xDYqIlEpKEC3X/8hG/vt0ri5LCep9qx
66t3jOuGFIs7NlXWlhlkG1G2Wd0oQqTPUjCVXUdSSxwHFBdT6uPkTLWCyZga39DZIcF9TBEeggOE
fvNTMQyaGFTGkmQDSkHtYHh3t67xs8zUB8bGjdOnN65Yyr8EfF8h/ZHvfjQv40vQc0/s/rtMUbrn
m0FyApvLPYDsoTRidbJieD3EuG+dh8xJrPV6/oL54m401YAuQgTyWjyeS42ewPGfjteWIgk3eaZk
qxKjSbaN524uMAZFIfsHwhFt+ev6zMYf8MlX/ldKSWuh6SGA/5ZmGMI3hWSGODe/j3X42PWkTI5f
OQpGR9fP7X/1LW8pvQrnnUHPgExc4TcjCxvyI+I/7C1fpNMKufPBh5b44yvg+bnao57hL73ZVeZZ
M31F4ZvDaSwDjsU7tVlbfSvMCfn7sWuahcILnGe/GaHl+xMvmnPJDFXOFaXDj5VRAJ4rAbbzlHKs
ZjmmAZEzGPjJP2BqLLiLu3yLL6diQrMzo1KvkDsuQfS8TEMPlzw7Sg0mqRkTXwchdKIsL+uttACh
nK5blADRyW8+Vo+jWHbXipPL3EIY8G15jPXEZCmHVxCFr7NOTZNUcXXwK9g3rhSHl1N9qD1xbWe1
++7CaZmovljS3GqpAJY8qiaJ07pjVam94amfKUuhQUBFeLDCxLjot2d85Q23MH6L59SWAQwq8oGa
/1WQ92yOg/v+OTzyx8IK1B4LW6UU4XjyM8AMnONKEZ3r6arL61WR/no37UfBzvavMGHuB+mf8dID
TsMzbk8hhQM4owQkOdMA3hEPfYyBYYFnDx0zYrCEcb/wnqM376k9iy97uGspgrN332FO3VVKDHNQ
QmixmQ+prd7mgJVYEQzMzdTSRObMFHrrymZlIOp8QE9TPY8UPOWwPjky1iOd5lqqm9iEmskMPG/v
7jb7pfJ9HR1XhkWvJjaXzkAWhgHkONae5TJ4mGX0KG6pGuFRUq9PEoZeN6AOkA8rm9IytuzQkC2b
9BEVnToQCxWX5Nf5cwe0b+e9DZskV9ExKVHAkknwpvRhFM4wbVsoaX6TV2MxEgNX6sB3iWK1r3KL
pYV57VvA0SqYmIZfBh0DLlHx1SI1HCvAE3Syjngizfaz9N+CNAeS5XUhJq8TzVoB0XoYxD3eODR1
zDPAM8QjK7GwssXhp+KGk2SvzDIFGvbBVPoPKQ7R9kn4eaEMstMeXsFOmFbWZACWrRTpkLALuC/D
ewJtrQoFOFmTP9PuHWoC7Smxrr7+y6MrKUxnsMTpHVJtq9/6qX3KVJt2uYkhjoOR4q3GGgMtVKfj
4HBh6ck4zbaP2cKUA6Ak69sY3Nhz51vv+mXE53gpxHW+iRH3KdFHyZjmCQLB5N6munrFY1SPJVp9
xuU7j0dQsq1nc16zWZCC2tTFa5I7SGsSBVgVICaa5aDz9246hlhUNoWuMAOHDQ2tA2cuFCXJ+rJy
MCX4aRGTE0JswvmC5rWYEUgb4ywPRxvNFgvBGNdr873J08uLoXHLrCKu8YLBj7tyAobCLDs9Wffg
LOsxaUwpfuAEGQetR/8ZdOOW8mRfVf6jebmKv7KWENxAgEUxrdNNSNveCo0DoaZNJPOCrYGuw8qX
w0koZ/sku6Tv28KNGRKZbKpA4kqiQTGDyzs0KsvCu50xcR/JOpBrEADkYYoPcLkGSLFOQ4Y656cO
V5Ouz6ErPPPXylyyyTzJbXyvF9EjRfPaz63qN0UsbHmcIRWEpIOQsXRFGESE5s0uwoj3ZMGLk65N
1feLYKgXUUeOn9Hll2KmErN43Eiz28FcQGXDalPLaTxJzO8RpkznEAcC0FicLE7Z3ecdeJZeRsvC
8FbVntmMp7Ja/JKDSi3grNirckrh/EF4br/Cxee+vonxcWn006bc1PwidoKUgLsVfd8cG/L+92Cv
U/BKlEEsuLNd1elzc/OI5UFdqlAvaoebQQjk7ii65aoGANHw2H4Fyr9ipB5PysFcygNxZbZJuCj6
nKir54nU2Oytbow/AvowISdw9FilOLlJe0/HvjOmqA+R1+hzVfKCGGXxA+72QmreF4076vgckVXw
//AWVeT/qbQ1/DOtnrM3im6FwVz1IBzd1YakxLf7oP69JdCY1JWvoUTY6/I/5S6F+XlKf6CepmJi
jzs0irsGIXo5pzpdboRnr3tdJbaTrf+E7cEh0e6ZDayIxEunuQCGy9L8zS/Q85SmdO82+sFZB0nS
40+ijP3SPp7sjpcMui5v2rs5gYm7I3Ya8+OSTteXc+TNAOegNyOO0JroMY+4iJcBp5mcq/RVxcOb
fFz48CRHHd9g4zfCSiHn3ZUISmtIQrXIMhjiCvya+3WkaTYwIokwHtehrVAXJobeADhUrL9z1i0V
i6eENsIGnX+n16zeAyoorOR4+PlKauvq8N7wHuj7jOzuQf9onkJKgxgYyUj9QrHzLI3fqa0jkpsS
728QVm4VRROupkB8JmTjtc96/6Wpckhd/rxGwLkWZyq+OMgs42PhP8roUlY+cZNlxiqQ13pLAFMi
ZQZnI2nD2kHSfCMTMJeZu47maQ5wT6CBVZnt/XXc56+81sVYbr3YbvR0Aw+CWvMvjszqUDp4VSiX
lvFpvhPML4DSZFpIiqgQEmMTAyID23NU4bDVI0xSfBq11eIFr26QwvS7j1O9UWY1h83YQ17Mbl1E
7Uksl/gJn7lQcZKYyjlBFJBcO4CFJSD8SOiTpEBjgc0KKQZqwGfOYwfksWwTK+lcRdC2ihcNr7Wr
xSMhRVnCI9+Z3X9Hw/yEwlMjEoo5GQQoBa7WstG2vXdmKOMl+CXfwe8nEdp2ZOlX8PYsT8eFuCUH
ZIhVxGo1Mo9uhAzk/99mS3F0THJbQHE6bkfAaynWi0RpK4ipBOOsZowcuOxA0tmTqgR1IsarQNvd
4tnJpGMzauPkvmrW//ZwHQp/42lFkxMOI3BRs/MGNvjAlDDbH1fa9WKcyaT/StBdymYxFlSZCkpZ
pCgVvrI9U3mAjNBfVjAEzfTD8TbeUtp2OexiD8s9eJgt222EUAGCYc4wskcHQlfd4vBT+nA/xgMy
rd0xAUvuSl/utD+7vccksR6Me/n7PqZrkQLXI/+LxSPs/o/bTQ86jtHT43FeueFqF5wzEwu/alSr
aPCbwr1U0eCN94VHJ/mPFM1s6xNYLezzUHaODAnKcgtZElBDtTkP/wbNzwPz6HisQm3jd7v+N8tb
5SHHWa/71UrNTDgycDw1yqTxfnPPn+mCUTXbT5NsPQmTUpYsAuiC9Gok8rEaxA7zOK4fLKLwOj5I
NdfLYddcvnk0yiiH4pD/aRA9LaLeh+jiWmDCCBVydFXWPuYSrMZeuPzNqWKzuI4P+N3Ic5vtDQzp
sFfp7zTwJzjBXuQyE+CakrXGEz/1YrFhwl0mRk8q9DyLXSO1vSEMSdUMT1wCieOvBumEb1GMESHM
SOqLBCDW9gTsHrDBsf8a6/B0tdK1qkitrKVSuwhCgrqQz0h2dBhEeLJpw7gqAxDbVAvDJj7SCnbO
ti6bIaNUMSC3n1nZmCqGzUQr9wHneD23dtpgA8YQbV7MsKQaRFVhLzgatku3g1s7cC2d1IxKxQiU
KqWjm5UXPli2wPmIsMejHh+7+AbJqeEHsYnyc6nPQ+B1huS1ZQWI3lLAKCT5VmwzKi7zRq7FaWWk
RNwhP1SSYUQhfdET4QgbR3COVPsfXlYHFELS7vu905yAZtJLf2ABI5dOtPVB08XuBS8eCoUmgNGC
Nzw1ZFm1P6G8fRieF0s6qSDcpY/nqDJy3641wtN/RlFtZytz0BjBbKD/9sKelQJ1D9pYtdPSN43m
y5Hw2CCjn3HUiDBgiBGdNMX7+kEjN0FUxQQf615UEyApKsyG58qsvCTDepSsncd365TYYdRP9fA9
1JZ7HIIbnY6HI0aKigOP0U7KdO1MDvbyc7jbuhCieSWGOXGiQN1K2zlUZiQYXn2+nZnUmEymYxYa
jQspBnv3txUq/47uA5WevgdcVny8EUZ8T04QDnxWSCpeGl69BA+mt6PYEWNujJvlTrgpW8xxP2nb
6jff0GBDtsZPHW5mZJiGAeygYroPnF2zmfLuyaDeJxBjOeuQKcNeZc7qVH0iDLlqtIxU91KUDNH6
3/JRFPojmzJaEEfOLPlFYwQ635WUg9PQ1kMAspzlfI550hcbcCetkNAblDezMXSEPNIc+ED7VOym
CmXKjbE4Bk4hliBakOvbdnULz1GSbaq0H01oBHFBntxhaRBpVjuq1givnaaF0OIEU1c5a9CAbrTu
sn7/5X9xs5ZFnCUf0dFP3HbkqPB95zuWtJfuxNrn+9xwKu+eGU3S1Rx3ZB0M00LC5tFrDnfIf0ZD
CXmfh9vA1MzcCfaMbqUNSI/c2SCK2FVSELXj9jYJOHcKdOjjYLvnER+y/ua5DeNfgWWq2QWeiCTX
q0te5xwe45xlLJvf0x7HE+Vf+QGQlaMw8hSXKjut9i14vBSVUuLDlvJORWj1HXsUwNI9+SagNml7
UgZATt3Pam9aYIFzKRVIQfxtPltbUbkwz1LqWUpVAOeUt0XK/8yMVf4FPWYQCBVDul1hAtIRwsQp
vn2T0z7XRUkSHLuMc32Nt2PZ85I+wABLptNJDfAFHR8J3kVCVe5G/0Cml5cTq/YcRPGXTtUNeTEC
D74hpRTfRszga+bO+yvi/cUVcax0jp4tvhoq4lyTEIm9sFxxRFwed4Hln4nYAyThqBkEkScfTgdg
G3FvFGKTPUgv/efZ8DOmVPuEeOD58Ri/06VHy6bR0HlONV29nBdxp7K8NDPR82hRT4wK6eGQxtht
YIzrIcRz/AZ7fwW+c18UYT34FqQKmP599JcA0ldlwRgcafYYjxME3sYmCSzG05iaonK2wbPPNCpm
DJ4X0doN0y8I5DauZIrl74HLK13OW1UpaGPi2OGHuUB9vISD76N5RhHzyu5OKctG4E+N1rt8Mc9l
EYpK+9e1Csz5ZF9BdmmGGocdP9nOCQTQYtkf8nBtxdfeIBs8rbUgwoPQpkz6txw9aLs7kWsorZxM
o4mBeF7q73si0SwJzEHw23tVDbc+0O0oEq7snWiodMdCLHqHJDTIXdxOl40qCiacd+MM0YPZFrGU
LJffi1tKFVn4cJoWmciJWxjvimCVS0Qn9n+nC2Gjv78QIHFUlmIGMQo9PWZLKxEtNU+KUPQGbgpq
rQ62tqHAUTiUTWuqLy1z4sR2uh1ko32o7+Mu5yw9f2gHItkQF8sb0zhWxI35H6TUHxaR43yy3Ox7
lSu8ix9CokGhHvuz0g5wUV0iE1AaGpRdc8SI+gsiSA5eN5+ga2GpWmlrc/FV3Jb1Mm9GVi77HVKP
oNmCMVVQiGEnNhhkNlCBAXAwy+NWHbYsUANFv2bsvmp5tIwEqnl4oUpSBtn+D7L93P7qhBO4uENZ
rpaThUNJO1Q82imiGPcBXBgCZp1Fhi6ZyA87aGoEZbmhklR83XOj8pIESQ2MEuf5pL5Hq15lfPx4
ShiPjELRuf8LVBXP6IFS2OodiOpnqPpVj7iWmP9ctniOB7hyLTpKwawgOF+Keui3N8lVZrmuz6SW
guVVYUbTcOSSoBCEbGHmyIcR4OxxAjZDZ6vWzsSCVCXtdm4agWHmgqBwFsaSySe9UMMgLs4ivdFH
bw2AEGnnik2eVwWAHQcVenR++4J5xyXXs/X5IUg73kZUFlBUBQ770527cGw6tRQ2wlMsNDBeK5R8
j1CMrrHYjkbShZ6x/ggWQnbJxd//nYEYEF5RawVxsWsVzYuB1XEvysXz2pFpp330KPHTaEDaGfKe
1DU4NPAprOa0rYTo21A8V4joX+CqoY365VKsYFFSNVNVhWQZSZGbKehwMjxZ5WAcuSakiT7sZY5b
WgTO9e6C72Hmg/B/hQUtKMveE1+eRUe8V3uOZu11T2E34NcnSlHY17RRiQNT9fuRalL+KYM1u6O3
WgGXKVp8kvELqO+RRt3jnbBqN0B2zTk0NluKDk8J5Qmfwcw7afgvpF8JU5NiRqd7D+ZMNiovpRa+
+TSbx2VRqFkFmBecGleyGh0I3P7fkDM8aarkz911a3DKIfKfcbxXclO9u9Vf+AoNWh9R8/4PR6OP
ubpCbWC0efWf9YPQtIWvf9Vlj9/lwBqkI0Boz0RJiP0YfE3zla9X+wc0fwCyXbIcVG3ZzsdzKTnT
vB9E+ntT2B0N6nPVoB10vM3X2AdEGgmQOVEhOpIdCqttZnLbdCuhx47hZcCK4yWGabUZwfxlY0n7
O6ay4wFugAbRPBeJ8Jd+R3Y/V6cosSN2Z6EECWlyOy43jwTZMG5+wqfKGDPM2ORUsIS6W65823T9
0n7hMGc+1eX/5y1b5rg2Vnj8rRSv3w9XihIimFrKVWyBDCkZx5SqZY3TimIUTHvNwA9iipK4OAta
j646BL7Bml2DFOVeZEIqnke01BIPoUDtiRFpee3Wf3mqDMa+JSCWiougx0silx6goZXZ4MtqsZSf
E5lkgTBPiVxD5cl5upMUTYn1Ag6dqEu3MR6Cs+H5KkaT8ksNLh5tRciJqajkyXakmwqjSEQbqS8g
apYuotCiBIkgbE11iMYyWU7qrR0z3/ILhpuE9/WWJb/TRwzFxSYTpU0/1T0hhU26OAu9r7kHy6m3
QXQ9IYMpIb4tM2yslNaEjMb2kPDKcf03wwOmxIamccv/z/OH0ryV/kCz0KCISq4gEoyYL78pPavo
T800LSn+pudYtRJL+1ebmwZmXvpxd63uANg5J5zhDA0dN6K+UN2ZOLrZw5zkPD4sRDqCX2SfEYLH
FP7Dc1GMJlZYnct7BJ6a6yxmK/ZfdkB1+iElTz0brC0RcJm1jAm2O2GBxTK2geYvFkj6EGMw5DuF
G53re99ZitfTXX13uH0AufLA0mBMD0kJZPaayqeVIB8lOEVnU6bIhWt6Mdc04ypNvyoLFDWVhpAx
P86+DOKbYtk8+3Cd8EJcKd2bsNVpngOxVsScRDXNefPWVEmiRu+08O66/vHl6im2YhsPedWDnSSW
2Rh1kTwUURM3q7brBAuZHPSCdJ49oAACpzVgRDLqTUFy1l3ViQq03ZDxn8YtUpXLuBJyXCKbF0yb
yCHZPMj7RPfWqQ+07TB52kFRrVzeg+hNnc+z20cTYgE46KX2FPWiehmF6DTTYNORnRahk8taaMhc
9fcEMOdeipmTqcBJ5cH2/N0xvVVGAmOhM7RoZtXWxV4CvKiiLmZbxoqH5tSCOUBXgzChKMpId63M
R2GdFmzC1ZhaJwg0b73gKy7YidaYBM5YJWJINTlgmPWP3MM3fW9XWrXKPnZYJ44i8kkkcYi4y1Hq
vTflx8nwAaD0LSMRGCpNJ46X59d5uXoGFP3FO+mXJZ3/aZ5AVmaOFmrEkw0bANcQU5HLBMSbmbSX
VIzSLMW2nSdQjduazFACjSk+FvGd3DevIL73kSyM6rVrB69Reko2PZB3ED8hcYdB19L5+nwasIFo
+mQBeHKRMZeWF9yPIfcvj6EdFx2As0SAJ+YWNcaxyHP+1fkhERfd/r0KBNvqmGVgGZBvugM6klVq
FVQMMlLlEQVhZpB7dpgYyJkq4lwJz4InrOccIWSuETwFH0ilbSizPEXlTbT9IOdZiEuvGPNXbW1n
ZVRTk7m9jliI7N9duDtUQtYUvMzCFX5zQkT0Uanhc1A093/me465eLgtGPDW0VTG18GtW58FSv+8
sSAfaCO0J+TTEqwfbHbw3wW9PBNxbTdn2AYiVO731aGKcJNhkjpIgIC8b+jD2gTniUtSPBmHX+si
bGqt2nQUbujCtrtYpHnR/GjR82/ai4KCZN/GMcfWxDA9TlDs4A5x0Di4r/P0oX2N8hOvYUIZrNrD
fbseETKwmqnwLTHWfK+JyJ8yj6ECTi4burE/hWsj8W/rp3Qxp4zAfk2CtZL0JVYvrf8jOF81++8v
aRE51RVrkEMHzQr1sMhrkcG6zqJ/gZMThGq4788chrw6CQGqH5FVJ5TSnnkfTp4tJOuLIVyS2bBj
Zu02dilSjGHo2+/NbM4Y6m2tdgmO6X5Bzi/e0WyBiCp6Orq2yIS7yXvaPcM19EOPxspl1B3u+A1Y
DJ1tsr+1LF8VfJQ5D4g6UgJCxCM8ARbJTmmBBN3DMlc8kS1JDGaey43o8ZAS5mGo2q31Puj597pO
ucyGxzbJ/9hIfv452S92ERuhEwe/cAiw0ChvHiqj8Z3SSs8ciS3CRbBGfth9fWulzvGk5AJUHksT
71V2+/pS1wiyjlRmCiJjbDy9slqp/8M6BhopSkvlojB+h8kEZ7w0wjbREghERk04nUPhSA2EwOET
W4oWy5QjRBhEH2Y3j3rq+shKR4VsNU57SinEQ9IokZa8FMyu/LEg7HavAvS83IFPYZxO57BslIC8
R9Mz1LyfkQv2NP40rbCRkawZuxSJXTVLZeKt0lsLn4msTA8ecfywrgZBnFlPLWZV22fe6QLld0sR
RHW+DsQe3zLxa/LwCbJAY92fmZQN74GILq68k/QSFHVhYYBfR/sFDxPjt0itGXQkkoqpa6PS4QDE
qKWimBpFwuo1Wg660+Me/QhzwTQvlYtXm40wNr3c4NKz8nIgTspDQB6OSrUfXaNe/Q+l5QU7AYkj
x+MjgJGxhv38os5UGtXLO7dpaVI8jO9uLq5YF9qO4nwNk4Sk2gAD5WpmFALGm4+LxeWWhWYtn4k6
KhI4JuPYAjEywdPLXa08uxOmdj9MmW58C1ml36/11YJUr4su1kdCx1FpjWAUud5LKIY8cx5FKE/9
Dt1ABxtRxyX5b9S7Y1K/Zfwfh44fwrDOkUjf0CYMqnq7DezrlzuFlukZoKFbuO22yqRafRQQ11WA
b7b0WNZK74UN2HaMHdL6lhjhorpX9dG5vNIC8Chj/C6x72dB88zb0X+waZouJ/uQW78uihX4r1uT
uqiqAeASjbXEaNaTFSkHz8wUT/5+ZWJu7vpPsdXX+4zWTVrcTktIGYSbgEXPTNhWPGUTafQg9Aoe
gk0EXgsFsqklPF2fgyiFdhUX4JPt5pZ1pFPK5zENkgRl7rQLYYMT12XkOwWwSBnooSbTdxsQWS31
ACXHVsRqjr/2SyhJ2WKwqQJqJXfCH66aCm53V+GdjEErW3S1VKK9QQhvy+p4h7+euXVvO7qHHTIq
OQrTRfjAGKjkvFlGdVM/Byvgox0aLSFAhNAoHu62/tuXz9cbomx3z27tid96u7luzTSdYEKRiDqc
nvbNiWNQ9oadEQhHOy8gGN3QEd+euTwqsfz9bxIp2ruHfRL1XvLNipfM0SQuGd5/SGSxb0prQZqo
78eRdmIqmIZOekMl81tj2dON8MKpRR0zE57cin1LCrnk9W82cGNGD0H/JyTQB1+FY2fT604wvaR9
D+QsN1PLl3EzJt4sqHOWGG8fwsy2lto8ZmNFJXAHMXqDeWbB0wiIIja+EVxmPuo96Kizj1Jo2mgd
dWUfhyNxejlZSSlXwD16KlB3kcJE+ozicE/uqkZtk1mjgIgriS7E1kP6y6ftgzFsgdrO5X5gwGLZ
FqO7j+QJSHEpsiflciyqqq6UhD/xZzRoWZ37StkS2tvyGgUZdcRYU9Y8Hb0ZUBKbt0zulnpc0Tbh
sA2HewLWaD/6739oE5bcTiiTBxSQz90Nlrtm8iJGZEs7yH9HJn6FedJK69D8UhjjNLZlK6rvM0Iy
J8+I7oArdpddxEoP8u+kz6wGUxf7Ujlpbj/FANV/jjj39Q3Ax1qVu7eXvvhkvhiGocROZeQtVPGT
kEhC6pPjC1E1lifbvnOgIK+ws1FDRNvZanEeHr705HNYtVh17+eT7nho7/AL9fUyoXePodsrF2eh
lRDRUOBcD2bjy0nUqNawPpdI87c8cRT+g2GTRwHiGoZmrzjlCtC5pf/lZrSPbo5SE7lnXb/YwumZ
oP8WJhSIbrIzaeJSFy30q6EIUvobgur2YfyXm0lwNmAuKWJaE9XN32mj5TTSxlN6UWH4BXNDaX2w
tug34ITpE9nec+xatPfzoVpF75VWEjw08N3QNgBDT8nZS6kti+g2Ig9eoNEDgDr7+EFbdT6qTHop
3dlhCIny8q2zinWlfU3NHuYcv4SBN8RCkZcvBacsag2Kh8RkfLXa8kBum8gxtEXCXzYfeLr77o8d
tV92+7bNuzqqFpqpfHInUAF6fdDFkf/q1IfBgL0t/fMYmC9x5MmkY6+2G5xL9eoPQ3lCbHXFCVyM
LsQKw3d0R2LRuIy46sv/50/RYN3R7w+zm09I5xm52YNYtiA977VPu0HC+KPsZqKIT6PLe9JkFx0U
hEfGRRK5AZ3nJRRvVP6X/9RKc61eQEcvXNLrsmkDvK3YURskiAvscF+j/aL59hO6RxnNApAwNK71
AHDILl0BKl1hrK/TFP3xhBr1rkh4Oq/KpyfifIPsQ4mPl8VWUn3N1cLQQrGAxYTYzHuvwagaT4AD
dFRuY9VShGar1k8dE4rtzfPB5Ef7l1ePhsThCv21hzEObF2d4cIar8oEs4TxatQipMYEGic+srWk
OTzELWn/3egMErwZcJNQ0JWyBqFgDc1CoJ1+rO77fQZZBZZHIaNg9IcvTzW+ZbtQbtGryMIHQHa+
krZvTuN4xkeZ5OB2bk3bnewAaYceYMKXok0kNjiZEVNX/bebypFdjQKX3CAkNqjAOfxgMSGkaE2O
JP17xnu/i/24+4gLBYmy2iShMTOTmyOw8ExfLfsJyjUM1KGs1N0w+ewF6NKs6p/GOTH8NfgVNPBt
4a+jHr51dYchmFZ7Wy5vJcqpWoIooVC0Ht15emSAedr8rlBO8S+F2a/7qcjrWOYceadKCQmaEQ0L
zVE9tbqttiaqATGZJv8UQDEA/zP+KkmsxBA4IY2ABQtC/dFZAgjfwoaZgVolm2oI5/VJEp9X2rLD
1ZL/xKy2VJMIIYFoGEjmJdnyzK3ZgCNo7c7DfxSlO29aSJZ4Ki3j2IowduoYLll0VnIvAoPUp13C
lacrNq2yfISG/IctSz4R1Eyfggc0x1Y74PvYRlbdg24jNYR0TWfjBhnyI5cvr4V9gWXp835TZL2V
ieyndwmVQ46KhILJHNp1GihoAlqO4oaoFU3X1/WXTLEXKpUVN/53NUpjak0ARx5eMplyfJp6JHQq
/Gr3OzHgmlo5PgwIOYFWI/I00TWkQDLic0n+sl50ijmNvyAzd+UWL4SX4mdcRdwUgH6NQU/1aHQR
itdG5bavG6Cro+iIlhrMWfiLn+OSqj/Ukhv+g0tMNXCYhDxnhDkDHxqSoHQiJYGsrSiS59cYtQhl
U70JEFEBpmSZpcu5kXUxQXIEnWD21TZQSz8cLYPZom6AtjkNzda74RnmPA5a6PcZ0YHYa0jdNX5u
IBgix5B/3Rex9cOvh93v76Pq3QlNUbO/9tESUVxuOo6uaygDMgWDQkatPjZOCqUjLPE8O6dSMeAW
l/laLN6QjEC15ffhrAtPiEunDq4UWIs4JD8yWbjsTnxaTlIEpBZyF9/7Vn9ixngcARZpcWTsiQj9
vqotvi8N9Lcw7MrUfFhCMYI35IUT4h6tENt9DTFLEwgcoAhmBwTuoLzuv1XAdKkmsMiWskctxGPo
ZhuKVMnlTJZyMrBnpYwOJHZpxsH0xGzLXdSQnGLorTuf/ALwzRR9cAZr5VVuh915B0qVxAlFVQ+X
dpZtlPscCfMB1KRT7BLuH4hL5DmrshWzgm0SQzOY3870wAFGMp25W4+C5SVfKL/i3iDZPRkb0bvI
wpRSlONNds/TdPbhoz+rUK1RE84fHNe03C4YOJVACjw+MYkXSu4d1zg2E0pXtuPfPUL0BsMT7hDf
/IIiLIVZPXgHC7nsWlxabJItbatJ1jn8i7jw1amteIZceHh2PTjNQKB6BLSl94DVDIDE3oEVx9V5
4k9olQ+JA1NhGV87bYGZP5W1r6r1Qq2MKfkpYU6Rorp7/4Z7uw+VH6TicjLkoibqHlJD+sH/FpkD
Yb4Q80OV65r/vn/wPyiM68CQM88bqz5dNVWQYc4AlI5na3wK303A7DfIqYdkdW8mtQ74zC9NSsPr
J05egYlgvn/H9N1kh546bFi4bAl1m07vFsNj9BNUVmD3XTCNC6QxvyLklJWKBPVxWNNM6f65SiUw
ItSu6Hql1gkU7FAcCRYpljwKTIR0j06N5x/UqucMvfQvv3ufTESyR+Qmg0iERe5mq1leZcgsiZFQ
1LZLgALsbDVPo7fST4AFcTC+BpsWnqlNSzL7L8K6QWTBrZmjeVNvA3i2jdZlQQSo3RuLqP4YVQ2a
U1+hDNUr/SXbboIKrUSdSMg15jxAwxEOPxDPKlmmtLSHAer6H3t58fSb2G96kSJ1plPNkEj7qFsY
GsSUWUXto7/o2JeGsKIv9w7/B3KqZK437e2AejhqsjY6nhpj08VQr5LveJhrIsrEP6eLOcvE26zg
6kgzpbsZFvallISIM+JQcrnDuNyPowq0OF2mCpGyxWSwWKlEOJ10NgWQ3gadygrinkS+IYSoa/sg
e9tLf4rYgre5lBl7PT6bFWTjWNZytC01vFo6g8C6OL6JFvedEuqtzQcrcII7VrtK7NCJRmJJukhW
lUbGeX/OYCiEcSnhk6Oc4hI6R6Ei/zqnXs9l/2eGsGj5EoUQW7OUHKjY3RbYzKspQa83J403dT0r
Z/Iz4WMZNHZBZlWuwmgKeAimK8bZJUllEBoE2aH8DSHUe6MBfJUiZfSFRaJ9JizCSkhu/rLiaZlI
9ZZxnclZMLf+t2v5Z90qxHRQvwRmVyV3g4AyFduD0ocyK1Crt4WTJJJ6n0znovH2uiWnFR85tEyF
K63PSa5TTKHvh35t+rwS3qrjC/RaXmh55U8vPmOjzjEU0deTamQaAXJr5tKaCupaQwisP/lCrlQ1
XFR43fJoLZIsNWfm1SlcyNjawhL+QNdgLJwsdD4BmHZ2GjP+dHRgav7fmjuj1rp+8OoWQ1k3yil+
pywi+KdlGIQOXMCH2CNmcDl43AjbL5QSwJGIdaoEFVVJQMxS+T2bbezJfbyncbFjpesFieYgzAKi
5ut0rAvXBDqzUwBi/W7ppXPo5fR+FpY0Zo6e+/5SSP/fmhU0K3+uiYjGU5YmaoCxx2XgAcVznUUl
GAdPNC3zpDAgfpixR2zb3NQZ0djVG4Ve2mniZfhvVG709jp2VMtAtG2lMOouxyAK5Hfv4goK0zKs
qqubdMBLK+lLjhLkDZWwID6jquMkVMUzXLBO4x/LxxIyQOZwcVKR1+3O3YZISUnOeHF8Sgav1kNX
sd2VGYOUDAhzLoc8crTgiN9YJKo5TvA2P1u/xe6tKigjhDSzVyoaKRxenoSRCjTxFUiiBJulEZYt
3bW1OWk8Kgcau37vtwt/Lir/H32j2SHKkk/n8Kng679PItclIJCRP4WN8cI6+DcDUfpn2nczazi3
znxvQy9QWeSr2EsXvZqh9PIsc2qqf3HYUlFijDCeTmmMAbEKTQNEpdytLXGChOOl7ZjyrD8ybo7w
a1SGeuYnCrw5Zg299lEt9WLJUPAlQPnO0pDpMW2sm8x/qNFD4H4fACzca3upHMstaxohHlEpgSIe
SHtWRvefv0cWlRjvNs9aJ6fk4Y0pLJIbqNsXrTCI0ekm2EeiLRyhEJM+kb0BuWGvWh2tnkpJV3jJ
UyTo8txl62VdjO1zo6g2l/OITEtl9tbJxgABk0t6snAgCZjVKZjQzSU1aZjwIQx9TQ2Y0DOontyD
f7AuBd9oX/ix/iEOVv/FnwOIXD6D6FpDIW3ttSHZBZfr9+GwgykeiFvh7lJBLoi2vtSrBdYaU5Jj
iB58sLSQyiv6g4Yw7zF/AlB/mzx1UGhm0aHohpCAx6f+sy5cy0TRswJDHnpsigCOviWl5XEcpI0H
Cj+W5r2sRtlBwXMFm8X6KrIwhIKL6Kg+Gj5gX+gC0nqVytWKsW4YQgX/h+X52tR9i21WVvLTwGWL
0MM+7CXOUMp+6jTvTwaYepJ8rcnEFXq0D6TZcRJhppSLzzUjL3Jz7MC7GmYqzJ85ErtXmjLlYRzK
IR+M1uRYlkm1myN3sol67PvfKiK4TpN1hHXFrV8C2W/TWLISiJbeoeuYTLeOlR+KnLt6KSgoa4Sk
MEy41Y1zZ64/IxMoCBFsTetCl+eyLoZ7UzDHDuDkjDfteBuH682atSfU8TYOzQddOSHm7ZuQHkDx
1k0PtYNjOLiIXU0yS8XXVIqjaxY8D24hWwYoIsTf0vHoJiZNnQzI42TxiIvk3E0Djq24VoTgTzwU
NqL7/85SqfaqspXJoDut7omSbN97vDJz9fJ5ZVcKeLuzs6T6d4rAAVZtIr697esha1sDHr/Xty85
hRPZRuL84oy+Cy2XrQcWFF3ciW0+I9xSKGdawCj8Bxg+TFq17o0ZNJGQBdHFOV6a3+sV9Arbr//Z
7lJBqZgP04yxN2dkEHvUXZC5JWhoE5lTWBCzPRwqd/hPPrU8eW4j7a0WZwfQBehx56mCFYdFLf4M
8zw9EfqI4yFvzTmNAUZF6odJeg8BoEfcnb4Z9wkd+CvQMnnym4BPuehFrPjUSfFVpT7sglqW3+r7
XTqVMSLL4sMNDaKbIAkqNQ6dKONWKf/7faiqpxh+gjoveU9iNRHZXiKJktzCXOEisRD5sNT2CKZ8
f5i7RyZ+j3dn73G/CSOKEW7Z5uzmWXHu++y1LBm+cuCzA+1q8iUV/A+jVB5Dhasiec7jjLR/YPAk
+9LgFeNGzDnFk9+xelqzd1Qx5ZZNYBir2mqX+c4kIrM69JRmT2B+ZFkcccicq/NEUkjbzrOnfZqM
YSX7aMEeEImxqMuCP6bVvOrfS1n/O4tCRty+vmFpgVde79c07SFDoxHEk09fIeRVPraXQIUJhsyV
7aB/kHShkReuazfUgC2tW3j0mTlZi/OdlWh1gStX/bt+cyqqWf3z7zsk4h+7O0Fmt9Mtt+sPRGC9
t+2TbfE6ntejJsKiTC7C9RSqS3HPhtIdLJAi44LnN0+Baw/KpqTELqHoKjh5eiLvjbP16ZGJE4sD
eAludn4eR32PPSTuYlYjwVhQlXoL8NufC/PnFJBYDITVcbsMEg82hzA4ZyhUkFfGhXjeUbHfDZD/
tP2VI4XYStAskj8/qK7XiRT8b4pMyWhpNkyRQX3yXhPftUUPO8pOPR+yw64SruasH2eUetA7OvDu
RnQtE5/Wsf11zIaXw0wNorNDPTu7+aRDMTuWzRKq/L4W54Xqn5oQie+84G6ENXbqAeRfJgzsqdtQ
iZcuBfT9ZPiv8AJ/h50OsFK5JKoRc4bpH3CAaXvwX9XWmFOSFKcqmdXxDKmPE1cteYB8tfhrAaL2
lNPj+A+yZ+lnB6kvQ05YyeleC4v7EPPbsU+6dCK56tE4K6jzX/+/zMth7XwJjtxvJ/j+lb0UhHbr
VnjCbaOtBd2RRTYQgBMQRLzfwsGNw7SxuELownMG59zpEA27/7r3e8XdBlXIV3Fk/GO7eQ20nAzM
K0RdS2o44BTs3PRw70XnWL9udn0/XVn8ZMeMg1/D5tkAgyPhukJRT+1E5mKxofn7H9sxz4NGvHPf
+SygIQ0oTC+qesFFA+1O77BPtAxphuPo/XK3VtqUzFgqJDO+q/nclyclXM3TZZMjAOSuBaP9clJa
+REky74SdhwhIsIWmKRplZAAKe0ipniDhjYK1BMR3swf9st6WJTy9PdSk0lMYeOplxbEfkPyTjX5
sQFYlteRseNdpL3Cavmw+64horpFAskyzg03VYdhaAk4xthTaKUaC3DUliXMOqh+by+LAff09XPE
3S11mFr0Qst9PeQx33iUGoVEJkijOe2vgK7tHyi7VPsP7WsUn/MZLcIpJOtKr0vU+gDo0GtdyRiP
sxlIwt6QGeIJx0dllm9ZtNUa8WIRNnVa8RGMkG92+KVpn/PZymCMNeTpnV0wXJmKmeGCUumRdVUD
x5kSXH5WHPE2Rr03pUXbNc0GV82hWvWzk250eMJaDLIM5U9uuUA66ZybWvJBdTe/XeKFXPh6xA3n
ee0hemEoEY7odCo7egHxkRvQA+sYTWBYa/wtv8JNzYoSE7yHeeWNqQvnUWBJKWlBp5j8i85h7G6f
+AelTHY91hDGSjfVyZyeVrLGRKQBKpCBSYRcayMM1gt+sBg0C0wUI3y8OktvnW1mmTOmxdW2IvoL
PpvxVbx+l1tm3FA2pHjrKub5KfExjFjUCeZ1ww9SpFKbhWNG5Ws8mkGHt6sEHni2Tu7hO/2bNRxv
B1ktXh/k2N3fLcrg65cUg1fcHUhCWcZOnMsXvfSLPonb+IkwQlQxcvhbPKzvlg1W02xgvfxWadfE
nFPgpdxaah5rPJdXSVPofQWDaPhxBhDzG2FjXQ7JJ+vRN8fbtHQXn4jDoEy96jg1aFt7z9NMECL/
vP7bHlO9JANOmDDhgEHOF69qy2NMv/KPUYBjS++1aeK6A4WfUQ+XyxdUnvVlV8PiyI9KD477eTPe
13xi4BGTTRn9aSmQIhn4USP2GinAAGcwewtWSDFjQXKAOjWCoMJMPKMkGyKWAU0atecHOku2K1d2
kvQCshEFHgLxn1OOZYsG9bkX601tEmaupN3x8uMyQ0iCVmNPnNqrtF2BcX6NBtP99L7pfSOjRUDp
fSYPsGGA7Y90N/th4AYdPEyBfZ8b2z3ChY/UIeC8HUet7aAIyvn4jsa97aPF5mVeJRhl66i4rlhP
NmXhYW67EB8VoTucliuG1l4XWpCrZxxDCfHsLfvTog7AxB2dJzxNjyiium/EoNpGzpUxwi2w8PUF
RpFCAXQRTNgdG/YleNwfnUY20SI/6XWl7eHvh2nSVjVYU52/ETh+I0iYxYNPQuhWEm6hcc6sLTnS
wwOOtVigrf0WxTVHb3/Ek7XUxAW1VPzRqHM+yxTbfkESF8DbsK1BqEV0xRyMyU9Y29jd0nIFub5l
a+GoVAjm8U7t+ptKcVizb8juQyzwgSlNVBcqpETMf/4whf106ZhFmneKsOBa/YIebloFn5BuO/XO
j4QFrN5y94EZIvxetvw1+WV37dw6UMQ3L27Rkw2j5RXeBBz/MIrfLxviCszBL3alQedPe8OkS/Ea
l6iO9rP4IyeiE93/cEdvB24Bg9pIbASij+MYeSBn7TkfHzpq0MMBVEQp7MZI0gclF/IF89z2iGZe
FjVYcGv5eiWNq11JldNXbIDNY45wSsC50enpuyVuFb8PgZtg1E+hS+nk6+51v6hboOkYlGBYiwyH
VEYZ+l+qvfazvb3WQfd6TvLQymZXbnjmZ3u3ehM6H2Mos6PN6E1+LHTnNaN7LArUSVUjwt1Pr/rf
WAJit+rEYKkTyp9Ook9lIoacHu67MjrbqgIj77gStw6ywEvsA/UtGJzn1tXAfc0r3jnph4UbnysZ
X/Muy8tvirc8X9qC1A4ZpanFElF6qYPxfScleVTioV95iWzmzDUnAiltLIAjJrD73BnFb6Y7SYt6
t56Qfux4vk1bpiRd4Ebjcbkkn8c/ZZyLClAwVThjnbGmE+a3KSv/4L0v4Sx5H6CkAEbyLkaKom8N
99hUYlQcQoK5X4Q4AONeBUtmQsWXPYzwHK5QNdHck3HZ8F/lyextOGEJm2v6pmSwS6ioiGXS+fx8
2xMcER4UFpJdDenyyFxCON1hS9ABH25UWf28sIpOhUVVuTHmtjTW2a9SMn0LWL0cDtwlTTnutnYG
EQ/N0FB4JOpPguq4JYYC9FdZf4NVUK1WRKGTksFW6cBmeDbPcsg60UGi1ylIAsD7kOS2KTRj1+4Y
iFKMUfgUFVmlWiPTGaq76YAchCXhOCxoZn7l1Dfgmk9Ijy7+gbHJb26253FvPkVqp5BeYAlRwOrA
JuKWYD3QaUqUJV0Ie01sbj1P6AA+KfSbPb8haOCAmETztGwj9zGNm2tox9FmnCuOECHxP7ozCUTU
weF4UAU0+4Nd1pLf9RiazRJxg1ZrZ5PIkb8vzOzf6/oDFXTXfOpAZSyrs2LKGJ9szXGlAMGNRqsj
+Qw/CO+vG2D7dKS26LIxvg1gaC4qCjBpJ45fVhV//j+ZrwXgcVM/5scGjzm6m3NTfiF7rJnRtR/S
Vhl5Trlso41DcGtHFk2WUrWKH0d/jWKvUbrJm1qO9H8g7pZ3nv3cfFz2oeF2b73D5iANfuQNX/2G
dXVdnFEt9fISG/mVjg4SSLRjxdjUJQdsbEegpeLitorarM8NvIqEvDuJObbZ2MAhP+QAjbt82pSA
C45ogj9HmLwAuo23A/WFfVBQ6r3jrm5UbCvhDtfkv7cr2/89dxpzKYsvoZJgIOItbeyY0gEZXHJZ
ZOTpJ1ZzQbv0nd8QSSKb+WfB7ySmJSmFlKD7nZWxDO+SgiybcPA0Zf8N3MXlmNcglRa7OA0Ch+2a
Oi99jbTREevMLZpuJOE1VQ/L3VKncSOxMNxdE75Uamw6R7eBG5jbJQovh6LCdhxPT/BvMbWhAlO5
tVvGmA2EOZO4jssF0bxsqEYIstG4dYBhyIseKygFLR/iHU6wS4qmydOppaVR38QmN237pqkMfFF8
s6RqGbhemfuz1t5UuXkfUswE3NWqQUGN83av6NbE/V15UoOf8QZ/m5k6hGf37Ne4edXO05pY+1Ih
RgfxLrS72JBZX13MzxfzeaRgjBHPcUAh7LkgB3TgsiKmVhF5oeRYNAz05aWgF1/nohkFwCbqNBXb
uMSL3dgkxpqB45Wnj3EirV3mJbnHcffTKkb5+84VLMNeSeOHbQxl6U8M1yM8GM9KNbfzziQWStyU
orEtwnfsZpHQHlgG3wgDSmBwAhi/zY06KyukUYEhIqLPHbhntFVGKNXgMNcaowTneegYadF06Nvo
1X7L5hmS6S/KzoN9/H4GV5famxeUqCp/Id0USuDLJ74ODWzHKmIKwOFICtaL0Nt4i8J7X8a19U1q
FAc++RzY/oqTzaOOx4dN4iKD3jNbSGe5xQZ8bBUmdInrKFNX7ttUCwmTLC+ew8njVPhI1fQIb/iC
pzyUPRyejPQlRcbUI0VYXDgeW8raD74y34AuDTs1Ph0S4DslVoRVuDI8q/pWyvGZJV+MGe+AGHKk
HiPdDP59C5dlv3oU3F/nT2lXLX/ARvdbH7LvNl7TtXwpdMvNjXNYmv+iAplsZRxxBRT28ZLRaRmT
yTkb2HWafEuBypatMXglVQI2zvpNSCKzwwezvcOkJMoKs+mRSQ8JIOpScvNW4ObvhueWxzOjz74U
8RTtP+iKp9qtSHiO2PRHC9iXCRXI4i7IkxUITPN9bZpEaC3M2fZcBbbfJxHQpYQxVxKzlMTbR7Vb
2vodYjQUHAgb18GKImj4foEFjDdqpXkMDWSswAZ13W1IlDWmso292vVDCjRcexIqJ43zkBBUTp7C
CueZGTDrda3SVcSWd1vj4/dccaWeAoqDeOxnMNs2DgxjyGOw0F67RzqTNwRmaM1ZyTHzukyvfS0R
7S8ISjeMHFm2vTM8d8NmG/C5IHzLQktVsp7a9dYqZQJFuW+fppw9kYTz0ysVi2xyJuaxr8FKL5Wq
LDl3vOtTLJSn7YdAAQCGZvz+r45bEc0smrKXZPex8gO/6YK9hSejJotsjVlfQ8DBONXF6IE+mp+P
9qOJmEYfwjvKzyF/kyRanu7jqD6lPefYOcGkPi9oubNbcJX50WGUKZa76Or13zR88SDSs5pkgcVL
dwQ5pa+V/ApJ0yckCWfGo8vhKWbe1JkDTxHDiWqnRFXQUOCHP8UIGfWhsUZFaSF4VhXhGGcL35aF
AFnlwPmIrCbk2I6l6D2l+YDvwRuO4ivRO9aJy7Eg2qXi4niLOTue/3f2NMagh0IPYIzuWoaNlc61
maOwe+shM9kodXE26ednIU1t9Pxfq3LIZGT/Tj9LOg+uXwdPDQ4alxPGn5x4c2j9hWshfkKeF3Gl
PbyX1axqJZRW+8jyfwtbVfl+mAnbctrr3moZpbkNWK5IKFbEAs5byF9JKakSeylPocmecE50aHyO
3xE/dw4EUi0beBLOQkIApsZWZI3baoqbKkt2dg0wYyAnNmUBP1h75NGYRsuQ0IkR3aH73rzNsi11
U0c2KjKM44PPHm5fGNDkSgzdKTGdQUPx+eQK/JgpO7eEx574765v7/YNYBpFfZbE2qAN1uzkAbpj
YpQrG7LOp4MJbge71xUyO4Gt1KYJDU3OpKWC/PI+gzaewouWzX1yIpqCouK3v5fxCml1uBsQk4/L
heNliOEPbMKtS4whPFbSLeOSQ/UYBl7ZjSat4G8JYCPRm8HGlLzm/EO2mcCttHLgptWK4KOHdRq2
gZ4N6JEqK9KXGa0+5fdlCaCWKYakSyenWWj0BjKL1K/zZHIrh6CXdqLp2rHTkHNj/4TDqWYfx1pn
OoY5iDeYLGF8C7WIkBaTvL5CRy8GjsdW+pq9DYunfy/uNJBGjcIzGKv3Fw8JdDTUqFEb86c4A6sI
/7Lixdn3yCsnYEOe6Q2k6JyGj1dN5xp0h2AjiRcI65JWAT6eVwXmQFv022yuhnLLP95K7cWgowfh
IkVYaISwzh0dtwstqZ9d9E1/+dvJWo8mxAdlZGH0++UdKyv2Q4lWu5caPKTYmY3U3GWag54gWpqf
tLMA/0mF+aN8V5vS/lvXa35eQwaXLXEFXIhODoJZcK2xkRoaaYoW4otQ/ogSXt1PqMQ/1zQEBCJB
eQe9CX8zcjq/JtIlC//8v8FsrRJV0RqHLFQvVrNtckFe1QUFc5My6RzZzdszgKWXlTi9KZ6vLXMw
b3dKNGP4qzTVCViTpCZSGaytiuO8mwd4P7aYLB46cR6rFN0xbTKZaHonfABv5SCconMeQDvHj32A
jDXBZ2JpdiA7GoKaiCY4I1aKhPjVeKzKgwLNwH/E2Pl5rp48sXh2pC7FZZjxhssUN6r7ey9ZhA5/
wpt2W1dql6AHAAPERgO/7aIMv3itYpiDERSFwxlNCYwsFk03HfOs/rbdbhP3eA5mk+c2SJd3GbmY
JL993Bj8yauB6FpTDKS91dfhszzGmrU5KWdMws/dv5qtgJCGJTQFUGgDiKpCW/PnCXBx0zqJ6fTd
nSnKUs9WtltLE3bnvQ9NEWtDvtzUXL955Vn4AoUpH3yp8o/088KO3pCUmbBbqe54/hGFKisPPRRq
eg2rizQwJYkHFmz+OBcWYTyE/q0lG7V3nJF4w5hKluBUtueYrRRPzmPG+cJP/eLKvOT/rP1y+Sol
tdqBaRhP3axxcSxQBRhH3zs7f0teBw22fOBL5x/lBElJj+b7EhBc36YqX6RI+nIIXuLgHI/epGY1
GD4gq85CqqXFW6PVtS1sxlyAjuB+ia3h8appIqUv6v1aMoG0D0FIUusI369O1uwhmyCXQnfdY5z+
Sn8QXLJMrsC9OCQM2T0nmGAFFjE3JGYNaTH+iIyUlT1YfVayAZj0W4jCrdUFCPC1wiV8LPLeyRUO
8O0ZMxHD53Ro3BIvKCJJO55LDa1lmv4c66OdKy3PZ5c+EuUInf6kGczmASORsc27Ycokn31PUbjv
VdydW94VwXgXxtL1KDd3cDHhRkvII0ws90doQtROVI90dysjxI3HwDq/Num3xKVbc3tG3VdzSRY4
7eon7N//Ez6UT/3bcNK4KRKGVT5+hDuMoh2/pjHCuJqAmIeCDXd329nWzhfDB22Gjj8m8Csep7HR
v4DgJIc+g0SFGSCrYOX1KcmHOyY03wHLVJaR1e4iepaDTRejaO3iLLDy5gpIyB/WcqGAvM4j9gSr
d83aQOuLl5McLBxA2YQoErapIysm5KFFxb4J492cj6/nI8ZZL21foZgwIkYrMjTxb5d3vqWowhRJ
4E3UySkUyAt6nDRb9PTayTrXZyBzNXfGtUiwEFPnFWwpm3xIOG/V1IhI7ASQFXdWUr0BxMgawkxP
7pPH6aVoZvbN4Yp7jj74L6RpqthV/BJLv0nyHdwMvNW8KWLTNAPQus97+Lc7dXT+m/Wj62jaRY36
w2F+a/8ghrcqH4ZQuMV70WC+nz6bH/kZXw3DedeAoIFqYJwSwO0MxlmGLgSvAvzD6AqYvY13u1w8
LFXdtLMdP7Qo5CfAOjYaUpFkwKQdgZPA7DROCwJXaqEUjC3qsdFB/vS98RZi6ndkT4x7vN8ox1mE
fzIuWN1eTC5XQsH5Vc+KZazDwJvw5plSvQsx8kh9a0cRNKtmuWPQoqjRlowe3VjhduArbH+woQi8
TtF+lz+ZSfXXNDZ+NtT+bD3SkpaojYDboKTn1sogXXVGi4AOdYFI56fKwosfmF4+AQ7mDWj+TUaf
SOTkJHiee8Hhr9W+DRcsGQ63PTi+kf91OIgxT3z1L0YMWqAJzoHdA6+nXyhlI4Td4j5clBD+0XkS
ZEY8kN6Klo0BGrM8PrdkFqtuiv73n42DnegkF5YBGADOxW97jlolGBd/kDUwCYizXuj78G3yXBd5
FryQpsbJcX6UhJGCPPgDrgMkHr/YMerN37JAGSDhZ50y/yTmd+4l2JBUKPKFcuCCP/9h+B5YdckS
w5Lt+R4rEzrJt69PsSA3o/UuLwU7zmYH9b3KTeJJ9It/fCiRwrztpg67VdOG1LrhhfAvKyAZ8Dr+
HPFRmS8hfVr9Q7hengk5J96Un6GeUpcOF2KuSwfFlPTI3h/FfvsnKblgcaHBpsi/67XgtYQ0lkiV
T0/OEgR+KwlftwCZ2hdlhc5NB2VhMnu7z448hiUvrV8DlnPXYHeOusR+JVaqvggGTuLO1wdSTuYe
KB9OpgPj7rdPe6ndGWcjnqBw1WnzdEN4PhLV9nN4bP5gn8VPnsdxtoMZGzR/ZfCLOAJbU/roNAQS
AP/iRsebKsap7wDfvajHCKsH3VmGfsT4qtyGxa97MHSNhANfLZryCa2dVc+yO6c49qDwNBVJr79E
0ZCTd348Ww4puacsV7sue5PXNyVz1KsbmaVOd5lv8tZZxHvaJszwjnK1OasySy2/OPCa8Zv9rLIm
RSemvzyCMv1OOrfcUHW4AWAZLRJwzjQTMDMq9UEF9SWDas5oiWHXBWtAMHdPphwOnCzpmrfZkdrq
x6CnQYAWW2QyqGVaVjs7meXv4GAx1Ox04sHmxn0LlTORBYj7U1bqhhQ2YfWbzoKZYU4ooHUsliNE
mYDRa84cYSYdG4gpCzW1xqEJtG1t9f3VhE+mUal+y2UayxCP7bHwxrp0lvUh3urUm7gW/pyCvkC5
iVTmRfBoRfcalHacvfa8w1E+O+2HUX9gHSId0Ix+S6B13zkDxZOaUQwFoz+hL5au7AjT2RaXMPM/
mkZQFVRDLKdh9RDH0V3yoOyvBp1HmWi2VsF/P87EtgWtwcq6yLVYADNp1PZEH+RF/vuWqh0faaFA
mhriVo/S5S57dJUocjGTULkfRyH7phvXxa6C+C87BIOTiIMA5bDnnAlpZYDbAQCzDzx/HLL+mH31
0Iz/nceAD9ArGrUUDp67L5flj5C8gvgLcVX8G83Fccf6ZT4TQiWTH/gOCIFpyVQl6PsjFr/PTUDE
YzzDJdd0CeeJSzBC6D6si/2dbnpaMqrGewceHlcJkfVFHqO+FCMogvpbhOSh6SKoElcefLL0QCft
8vr2y6zvy4+S6otgp2Ch2JIxYlBbRNDois5nBTl0v5EYrpQjSWIjXMq1b/IKWIQIRG1Z/rJhuzoq
5ZCDwxCjE3irDVTA1oPQKjM4AUt9HndLKbaZQcEVNLeJFWo60tTP39+vDtyTX5AWt3HGDjZhd2Gz
RM+3chU6gTqR/n6Ywjff7tmfqrxsby6wsT2Nf6WvgcFNYSEseD5DYJmrI1gY2RpB5yfFxTnQs0hf
s7O5x1pQRh4rS0lgvAhFHHJA3t+Naeeae4sYJCnx2vcISKG5AA4SWmnggjk0BU4Af4Yp3WFB2dr+
LVdapacSYVls2SGFaYSl+xJO2KijTi2h8G1MiNnMRjracXoWe8M27GWy7GVUSVm2lgcO8W9Mwdfj
dlJqIlzTnXuO+9Qj1J2K2+RO/k0VUSpqHqoMivGvWd2i/uXrrYrP8nDgN05pEWBQBORsCiSO6pPO
LuV+9HNqVqJu006n0M8DYcc6bNyTIpbU3hfoWajGRs/p4eUyMNv5CRY60KCmfYL1JzdTD9grsZxk
uh5Jf3MbUJ2+q7QjwvzRFWLyWy98n67N+dyo0bPzyaGNclHs/kmBZLKGwk1e/6rfsXCgkgFmT82e
+Rvzv7OKnzF/yfbolbJlBOpCIbKQgjnQArLLooKkCi/Jm0ZB6IKEs8UJatT9MzCCR6wIrt8a1Cdl
OSg5LphijIZxJp88l88InVv9w1Tr5vSCyad33HbdUzKSS9FZw3gI5fAu4R7jJ0LqWIOisIFDe2mm
B/yc8zKLFNB6w+y9AMa91UkxD4pVf8ynDA1GIBBbeBVZK6l+wG+swm1IlgxMf56s6EutGbyCUXTL
jBIXxwxYJ/JQkBAZGFjixT1IgrcN8ZYlCpG4bTiR3O6qdS75Tm6ADoaql2biqsTbDNScvsh0eAND
N3XMdKzvbs2tx4Y+IQG7mp/bPJJE7s8/y15g314ERKVfbusueSjfjetsfgwrFryo/+ALVBAmkX5k
ftPyl34Iu+PpqsrNm4kLj9R2naL2LpXOOu591qUQwXlxu7VZKpzmB1ORdsKp1owGrvOLjiFiGlOz
n+EYDCprNWU9UbutZnEsr4DbusA1qXjzGxuuAvxiAuYbQrjAtN8zn41Qt+ixrg8PMzY+7Cri8jnk
FJhm96EzzczOqcoDgCFC72jSS6XqGXCS99uEUobA2ZelRoSR1xo2RATxVDcwIZIQDZHe0o8Fz62a
j2Xnle6Ma7xpaZinc7tKQVNUrTWasSVyipCf7j+Pr+h9BzeHdMHAxkR6EpBaxX6KPOeNI6tRUSaU
KHqjhTx0DfJlQi2NH01jt1Y2h51Yp2Cld8BAdS7Kc6KQ6dtWvsm61U1f9iil/lIMQbKhJkRqeNSh
VEy4EpSAy1KsU3Wy2shgLhTCboUSy0IWsLUM7xy19Bs3VSpj32v3x5B1JVoXvl1OjV7DHPDS6u9J
wKwlJEDOUkbJcwQpigmDCpUlYuFVpQg2vNYhTrajdaLgkFnnY0UVq76wgxm+Y38ZmJAjT0jEY8TM
FzVGE2rGA++LxEFnTOVR+Ymh0gYpBVjzaMK6eNMbFBcf6QuksY4b/24XpYOo9qgEIS+U4dWEkSM8
6rSxv01IE3I4f6A1qtE9gEa1TFH1+SDwuW6o6z0Z/TWW42zCYlWSTYa0e/dUVikkVhm77508aoe5
IXnc/UBt8XbmZ3zbax6V3T+MiJIz+abLW70+85AtDjWHFiKhAGIM1eFuP6uBRxsGG2k2ZqKTaOjg
94dnmafI1aKv7kAyO1zfnr92Q3NEvRBHgnfpqAIau7z8CvN6v8u9CnnrvDUVE63AEsCn9BIAzVSa
EJxFlJtie2pKQCPAnkgu4i/JJc35dcfAkwyPOBXigBy6hNO6m8uM7HB2vVMajTWaQjfMsOS8HP3w
ncnKXsugW74IpkrKFWmJs2Ps+zjGtSNwikKXsYFTNw0mGLcCote5tY3HP+oRit68lFYvTtBepFb5
NNzl1Z9jGJSSRNAjBviDeOsteOf6kZF2t43i4Cg2Ln27w5rNr0R4yRk+GFiCoQYSv0LbFpFRqldx
L2hmZm02LYvcy/B+ELKsmxOLVEP8QWlGHXDDPg/twz4IIzdkNRqrwW09OvNPnDueaLtjJ8UhKeaA
R+/VdaHOpVW8nFj5fdjbcy7uBT7Nj7+2CTZUbXjNCtZ4pSqz2MlSjr/we/FshXuotzdOOutW49kT
yis6tGxaziDtsfKLS20qaE+9JEwmnM8HdWl9jvYYx0H0X946sGrZaJkQok9VgySTSlL2GE+ICJMP
0LKv9wbkS714ECTwoXdZSNvmvQkJplRzeY4Eh0O6Lu4groOzo9wVeGHadYoG2SC+3M9I3/JvL93l
cv5TFbE+vbHn9vXNgkJ9HhJRMqBRBTLsQtxLxSyWNcyhGhQxpOMouW7bMr/9nXxX+l1bpECpTgaa
8H6uiFr6anlo2FlxUe477pXWpkHrQcVXj+YMA+8d8SdYfQQtUNgaekhn/7nHT70piwtAd6jB1Px7
rMdd59Ia9iTjGP0WEXsSUpws9a18N/NhtDfJZx/KoFA8Yrp+ZsG5IklKacLk235vhrjVliyLzNNR
mdh7PcgV8ms5p+nHih2jk4oWaSmU1UfH5wwbCpHPePcthjOnXxfMdp1K5tNZVqhBgPAkc4yTwEBF
2UP2YUfwFPKeoloFNbiYiLu3gbwHeWWIJZV7wOf/oUPwJo5zhxjheNquAe1Yq2P2XqxKu1FWlP3p
mtlfLdpCMsxOhhNxoC1QB5SpO1fwCz5Sa//nkDfSTv1UwVY+N2/xtXKVp3uGobCnOoB8gH28ec4T
8aObuPaiL2rnv7L5AtB8cZOqDdkrZNZo7vUcCWmcz/GDaAOZK4Vsv5qt6oTvkU+Ptia1xhdUoinh
GaPDUf7e7lSolR0MQbydYYIesWEEj/dSjhFFK5EQKDWr+aO1k041SRNZSPrfhhNBHcddg3J0x9Kl
vVq2VnzkANfpZ6ai2kNKNpbusH6IV429IBCPo1kNitnSTC0W7Nj+cdN3XcEbZaLxuhxPsiEhTvV5
MaJcHzqu8+KI2W7MuVA3rE1ZtYSwqETeTjtcaXTe0dSAUVs1eya+VC2qn5e1lNxDQu01rlk7gAeC
bOycig7YXc7a9iiIGODvVmWXQ2WR0SYSHGwZ2BJDqUEUvg5Ghfo76jFTKH1nkHE8M0KrNGbdiFon
+3+LTwkWqrQjboV5FTB3BayWP6BJHSvWqs7HveI7CW5YanxAW0DolioaCPieohKr8etuDqMrHM14
NeGny7D7+FW2F2jnVubRSn9ywy5AVqZbWZXFkX9WKh3UPRU6lrd3UvenmnX/nkrO0a/8jAaQVoN/
2TkK9RbI5rLgK5coie0BZ6Vmvah+ntO+heEMDZHPAOMV800oD149WTL8LR9RDtdX7w9JX4/Os10Q
YRBs2bpqlbpeaPHgqfeI9Kij/nqUR7aWlFxIv6iKBp7Z+IwXK3A/VYtVQN5Q6fMv4AsnmlBrMH9a
IZNFdvf8akkRxwI+FRFGJYDdh8k5cqGrFE4zsMRG61z/flQWtPCrGJROlWfpeReUFHBx4f63dqSI
CFOMqEyYTOLyMrpARaucpFqwiGfVdpBJ5y6Z1qnLw5fSm0LQo+FBTEXnM2c87xhC2TzpDp3ckfvl
phGNCPYBIm1oknuEj8+QjM7U4ozz+MVa0jj8VNe1AhUPpA6VKe0SgUtM3GyHxFy60+e1SS9tTmJ0
cpUyDg3ic2bN4m3Tst73slyIlgEdSQB40/0K5xL/j1qkyU8aXDt2BvNFaAbku9Kzk6yLIyGgDCzY
ZIyTT1odgCwdG1JLx1g7qodWcgaUUxF0afjBujNqrShUWMJtV+wifg/+5dkuUgEO+Y9CDiBQXhkR
rQvDMsLYvGKTTeRIhmLjPf/x1BvyR6FOeJMWMODoeFxfCAnzP/9ODkXA049n49DMBTUkNKrGf3Oc
REW/RYBWuMqIrDsGH0ptj5b5DkdhXCO6WO1zg5+WWh1E952K+4L0ZbeJxwltj7YdFJqxpl9DH7kT
kVdb8zCjoqefhy/rGduoFFp/CYFqe7/uN2R53KeZg1kA0CyV73WsBVzKojPx4qhiXNXbVjtZ1gUs
MTRTu3H6QITSDIn1u9YlyOOk3laT7F0MgpUOntmO+0S86qINKFYd5iywCY8deB29xV8IsM8xxllt
4BqQm4jl/mfuNveW4dh/fDIHr0b/MaNYN9q8d0AoAQEU1kKQF7LKHQu+zicVytq2b1HBl54BSuDE
n8/Od+Iqk0CWk/v6faZ/vEFRR+LCNs0bHv0NrlFn2gxG6GPZQdkFXt8VKmX5HRSk1o6CjSdvN9nC
mACmswjrmWeqwKZVTfnW2KLU/h59+0RkHRHYtRwFE9FrZqzxYZi8p0bpHOJjoNie+it/8NjV4O75
Ak29kyhwHO8MOl4O/bwKIIKFeWPdYQjy12TAjA/paxgePMc4Rp//7jlT18d2e2jbechlQHt6ZYfJ
zOBp10Vhs9tde2ugC5OHmz5xFhMLYccdG63FHQx4xZA+A9rUwW42/QSONfEDXuci7sqSHlJbSm7e
vUgvGznsO3g0GZcN5JG0G6Zh5ZNUNE5p9ZkH6ISw+hfwSqcQPB12U1FTSi1s2lpSX0VJghd4Z3VF
VYRUSkm6GMwzQxlL0CU/a/qOA2NPTBxdWSOTb4Nr1Czljx89m0tKiLoDSOVi0dBDrp2HGIoN4sBh
VmZ9aNmMln9+j0WKfG4Z2qpBdEi2nZn71E+WtOa7C5jfJ+N2mn/Q0Yv4rG5Pc6JfHXluG3I87Y9s
OFBI64v0sUz0LmR86daSmo+VJSl+QGO5aTUdCCHgti3vWucdasoCKfeq6ndKMq4ReuYhaf3G8Ez7
GX3/92JM9S9c/UCfj8i7/Zr7k3cjOAW6I0ZkVYr4mgFxuDcO5SeHpv1FR2b1krecf8Snwnmo8f4C
qebSZOqPRBcxXvayCd3u2Xsrme9M89usHoAwbpDjaf8bKX+dDLhzz3HAH0b6xFwo4/I5MYfPCoC0
8Hk5dpgFO36E3+0wWzh+PIQDp6tDEb3J/CansGBqLQl7EEZib44+cvJLeby5xfLBXEYpVa8TbXIE
x1dcCgo93W32S5AggqPaU/quotlCrvnhCX5/V3U+7PFH8as4OnaYkPDSHcjCD/GXap6zHkDAiMFH
N2i23jiZ8+09ozDtAW+uX9JUV4Q/lw/6AxxaVjhPQa7G1i+lUoDF78OXSkVRMcDzz/vKFsa/BrwY
fRru87K/kAJzffwSbCZopg8wdVOMrRU1EIghEqVHJwnPXaiRQUd/3mVfgfm3icSD86qVLFOkBbEs
xY4YDkcGOQUgivoq0WrOaB3of7W9yXZWYTPF7ojWUhWz94JGDJMtRbNUGLAqMn5euj6CeEVFe8MH
o7u1KoVdvAp8FypsIIm//ncfHA4irhuR8dPnU0M35zky4rB5+xHBdgQJR+v5Uv2WbOHTWG7QvAqy
Alj6HKqJADqMBRi4DuGLbPttfRRTjKbtPCRWwC/4S5k+LPddLd++QCLcuYcLW9/QGG0EC3DmpGzq
RM4cw1XKtVKCrgk9fnTA4O6697smj281Hfbt1EFTelPeUJ1zfw/z2OHoaSKxKMEWsSWi+mMEbhMZ
CYdrioil0HB1st/soAiz/7S9Nx/U7aDSYKhNPqQQRrduNl4fsXxVh2K0D5biL0spQAk6NnIYbmc6
EOCV3ZbwJ6NZMT8F6c7DD0w3u2soVJb7VEd80qLp6QxTkqSpEdHXxt5V961Iivua4L8Mbb9FzUvl
Lbk/ZvjlX061wPiXV8PQ60686G/nLIe3o9ak5wn0YIC++XBOkQk9+hIrz6BT+Jgkp5Gdv5DsNeuC
OilGt4RC8SP2wnlMx7dn156DpfnyRWtgMbrsBIelzZWsrUIglu58Qmh2wDrtOnT3q5OWp86NCA/U
6BQANvJFiBOnMoI83o+0CGtPtERCuWtzL2bT42ImPJAmuFVJyeSuFk0R5oZr/8HfE11UJlU11pxa
7NpgPmiSabg5HvZVcpWrUU+JLelE+MrPFJGEAzrcEcsA/LVI97kxM71Xkvt+gTaec/Z3nDnJcrG7
lgQ1B638W5EyroUxHB3jwQlEDYg7ZW9dhx9U32sBi8L5vGnyWWspa7joXw5bW/efFQlpGASG08Y7
Ivfo9VQLMgR9ITzZQ4KMfsVUFQymntf0Ke2hIHRmfVet42PBwq0EZFxxr/jfY08tn2WR/ktavENO
b6zsUkcTOkItuLzpnxU9UYYQEshb8Effh+HPFT2kQbUfUn+qqDMISKjif1PVgczEdFNr/uO9Az7I
wziCSb1r2090WUBwFMb3InhQTQbiyTH5C9miy45JG2nt55kAhNlbd2H+fSAcbbdW0CDew4EzQOMT
krW8liF8sgKS3sCZEOmPpPuEHFRq0TxX/jB+rRw68m+idQXGUVM1l0DEmJ6qCBFSb2CKMgqdZqqz
TWk/jybEPbVbZzRNZkG1mvLybDj/9vBRXQ5xnSBTCiMw5jmgmWBScrbaFoB93p6VVI+O9MtoBQP5
5WJpecqA2jJIRhQHxI3zhe7zVWS7SFTURWWu0TR7cP82IpOkXVNnAIq0CQba5bF81Ulu51CHj710
WImeSy+KrzAuUOp34CWzweb5tNjPKZwEueKNy53UTSsAJh8A7+vzEjyMetcLAELeC6OFywGOTk6K
C91Dk3uDU/Q1rMy703UuyVBnfNJ3obtpGpGbx2USRqfIqLcLsRsokRoKh17hSIlaIVdy0hBDl1oF
MoQJNgp7e+sdC4E2LL13e/cv0albN2EYXK8ee4szqFyj19grqtfMh4Tvzf9My47b821DpbQ6M43p
kZaPTPl035uTTdaxThOH0auVoDFVR8Wo/2geulXZOalCUXBZIQnsEhkcultaiYJELul1NzRTi54G
VaIr9q4ZmQh5kwjTxt6KwHQClrlCQH89hx9TnqqkdnWTwVH1H1fOQFkLo5t3K2VLa6idf/ALp0BJ
0JAa27q5sVwqQwbJJWSgfjsrFIr8zysPZ9J1lluxldVzv0pJYtNtOpAkQkfQU4AJllJyehK/VI7+
kIRoN8ObEhm3bhwHbqrGw5QVAT7OXMXadgAaIJi7FgnxQJFxDfPz9wh8RMgRwUD5bF0zED5eMDEi
2OgDekHZ3pdTWo7mNg3d5aGQpcAsvEPDGBJ3dnpesmMc2zTu5Xdz5UPO87Kt8zGCzAD4/Wt/6+tn
rhh2Tt3nwWm/4cpXDS6lUgUuT50dVlNDnfLSsG3n1l+WleyR41t/BVe88mB9xOzE8DbdBXU378jg
7AO94w2uoJEJnXHgDo8dMWNqgkJ3IaV8akikKyQzKdvsyTUrZ9OTWCITkKkOFd57wvfLMjTn8KD4
q5nvNnc6g5NHYQ0VWgmfoVfkUYYe9jeULH/XVu7Ftz9HkIi6nGbda59QZXjRn5TS7Gx3bJVhA6xd
6fKIuWGbtssfbUcdECseXbhRSPtZnk3lDErCerFr7MC6e9gDe/mJBMbyIu/vS81QhJitt0KNqT5L
x9UbXKC7dAOJnJP4N0/Z7LBFRNPheJSqHZI0o6rLbi+L5Wiq3j5llD9Dse5VuYGF1ven4ALatSUi
8PHqTcSs3qpvHzYmQyeO+DdiRucEZAWzgFoacls3k+l4jOknXtNW15IxgJN/i97bj4hVBvPaqa8y
XU4sdN2sM7qGTEJZ0z5yOVJSOvkSzPYM607w8WHlhqON3+cgfUznd0NL/ctpfN4ayyM2A0XcglcR
aUV24viVtBMLFWs+YaG3gOwe1Jb6IFGI8x846rM7OURi/jk97By9VOpsPOw4rWkrj3boB7MuVfMW
Jmmel1xwPF0oK1BP7rIesr/3WxpV4LHuIeHvOZpZSAK5aDjkRY1ZG5QIAv5ecCwVELXXJkjtRIjJ
Qn3PbUGVrUwWA9zKDrV/wvMQYU+GJzPE/9+B/owovNN/iRDP2ob+3OJEgaNJfowfuGllJYxPooUA
9kOH3CRT9cOHwOD2vttLnS+GYKr8tjGUEQiyPe+e+HqJUaAdoZi0fjBfCLoTN3zrCKsXaUE2fSlb
kCVtOPq7JxoCZkfxQQwQ46OqlZGxIuEpieMGW83iPmDMI1MkyoRoE4phQJb6UYV23VjOsDNBZKDZ
G91T9LMuiRqU+wVwWZgACYnwsLemsFueSPQb90+UFMXr576ha2xpOliNpZ0jTYDAOKcozx/NJ4cM
wC4iccP8irjOxYtVKzG1dKI+ziqwZv/9bQZBLbV+5N16Hcr2k1+yslFR6gp+4V94e1iJoUxsRmAs
kBKeQRwwl1je7jrPzQvKF3W0a3KPY5UZ1aVzyNh9QLHgokcT3DCr9ptMWkRz+l/+Jr4heabVzmb8
CMuUHOiybNM34hFAVp1scLnVpaKppCieIRkoxAnDEK2fb5B2cC+MjPQz7B8OFtjcSACgTNsuCdTO
QzdARhFe8AAlMVg2WBA3HCEKrynMNTYAo3Yfnn9Nhr3gQB0y+MotmHTVT1SR6SZaf33WNYz4I4N4
dLkwdsi5OKSKAt9I3rjET8sZGWidV19mrVsTG9gvZsWrvhEXYi0BWyD/LkQgVz6ebhbPhgCH78FY
PhBHaTtHwz5oYwOxVoL4mMniVUybZ1DUrPciQJ1E23l8GaKlr6bCjiqLxGZhkf1Kh8e1La2pUQ+U
kQrI+FNAUwFvt7BygvyQCP04gasC9pK0X/oo+kGp2+S6tlxCpMdjR3E6Lt/P23KVpIlh/0TNUxHk
HmOIv9SMNtvJ90Kxb7bo8E2Qlmya1vNIsgp2dZGY/P6o1GX9YHL2NK/lzMUmbO3lnB6sVH1ubh3q
gIo6Xu7DqB5rSOJtLqY2SSqtepQRT65KPeNaTFURjkP0YdEuprUElKuDgkaiM3ziEHgKzoyDR92n
JwI0fP4dj3sCsaGo1tqiCukJ9tR5dU79FCGDuEAyjM2xBuaylAP4iJ74Jq6dDU1EbNrN49cPAzqh
TGfPiPxfQ8Jj9ofT0JLTqdMp8Outbf3OS2gu7bw0XNS0xqcaD4+8eongMKr5aljKH08XN6DCXA3c
dXh9QSnOBV1r+rIY2lyfw2R5aw2+z2vX8ZqCLQM31N9Ma7XzX/r6bC2Jw6aQpJMaeXpm5CsqTmFP
Gusx5pYSeeImUqWvQX1yU9QVmAlNuIWmTwOeAM5xn15/7U9FnlG5ASz2RdeccaGQX5w3Kx6h2n+9
Fuv6+sQ+NVoCf5JQ5KIulv9RliEH4WtaLTG9YlTq9Bk2wdiWfFe2kVDbYlbM+6K/mH29/xwOcbST
PqnhEjywifBUSxVy24nPKCeH1TR9azOdMdhjzrjLBzo9PZh3n65+Sa14+rtQXJy9zy7SMiVXKfKl
1HgNhXTRToOiNED0WCLz5QQj0CAO932AvV22e6o4eR9W0dFYp1UlxqK6hp41eR69th4kincPUDD+
Pohg83YU1VnXH2s9MxPfpkZMOATqgnrYYwMM2/GLIMhBf7Ba9Sa/EAqayab+BEagdk+XCK4q9t72
ze2GJTSBiNC+u1dihgZ1HTiDvTZyEb3ZEd24JRsyK035uH4qhtNa7P7jvBpZJyVlAex/eNeZE9+j
fjtuoo9M/ZBJ/4R+vhrezIIbpwczKop3f9zdNjA+VndpvnoqvfRZnyQ+syOYwOY86VGS5c4kUH+a
pftBEdtMZU/UKNVsiviJorXzge9zoguLFtFNLCXLvcoAFk+pbebR4HtVwadxfUKSTK1QW4gQ1qDH
rgSNdz4ph9K0vjNjAMMlk6u9mhFkOM9xtG779sxnl3GQHU4+d5OoolX67HxGiepRWVT1EFJWxOyS
1CTC2rfr4f6rWCisEKO7403xrIULnBMiYtmxGa1JEgclWkP3/6l2ttij/C9ddEkEyWhkzBnGyVjp
/QcMOtKdRgSWS5lcDiRTEo1rekia3wrA6OiPkSBtgv16QilTn7GZZK1mBh9E4nozHbNiIHTsZ21l
ZYSNYU5x2bcHKpc4DgBn6mX6DxiAAUWEchmNP7nf9919MFBaM0DoX+ilt1KHHomrOHoxO+0hTGOm
RZA2qtlnHcFISIQiCaRMGmRegW8mUrR3lthIj5mpWZHXVxoFWJtLrWmkdJrMVlj3NyJ8x4F5cvGF
lj7qrTVT8mWo074gIQsjY/CjZn77cZaEi1+Jn9GfHso55dhC65uNJNycqXaNbzJ98V3QdeyCGLxx
EuktDAAYSDjesMOjNTUqNPX0tIJcKfX7/PNm9L52ZGHi3DutpO/NwCn7xidRL2QCxef06n8+2BVB
i456n8gNXZ4ZZ+nF6btL5/W2gXaeXaKQG3JXa+iAW7HkXGWCs8Br4sbUXo07We2ifH86Ojr9MhLw
02ZPaFv+KHJTDpgkt2QjMkIMV+UVD1kxzbG00+EkvscZojweKAwzAv7VvsdVRk19yoGeLzrSSFLs
uTgVJUVl9DTvDLC3biaq7qX8EkB5dBe3kVbd91X6ts05dg9fNpRXHf8TWpLod31n/strSjWsyzH8
wWJSTP3xlTQh/8rnWUXhWwYvQE6JIP3QVrdgKb2JJ4INSAN/UFojsDBHaLP1sFxLz4qvaX4kVUx1
0LRlQNmDjazKn0hm7tUhcWbs21/EdC+vHHu7DIZrQeUgt3ZN985C8Q/A7bAAiZIeKd6XjzQjtAOq
C5QqAco4hxN8ZmhVfCjS8mXEk6laPjNELgE6485bEt5Y5g/Mnrk2+mndNU3B0CavfxlBlNNe1B4/
frEaN29MMj2PkyZfRMSgFTLGcMgyZaQPJv1kmYRxVvF1Vd4AO6xzLSGj4+pcDpTnOpscfO8RBo8Z
FBD/tdinxFnSpPPdrcpQxst3bAyXHb+0HBHdzwPrl8t1L3KNFksIBnJkQXVzuYGxtKoYIyht8K8+
r2kGn/Rn5fGc9i2ssIAzPnq5sp7N7nfa+hSHbhZ4ekr4v3urL1UFQB9migatsz+mokUl0CxUdlXK
mP1rSxf64YdEOr5Ld07wZCZjO65c81Squ7yzMfQjv4HDaLJQDEagH5jEn4zprPPkux6/Zeb27UYD
vR+QA9oj+RQYtlybMIYxmboK0KzuocQi5PjYRsSjkGqsPPJ/fPB5l/sCecIEVE1Ly6+rJ+4Jat0S
p0QHx/FwZEUpjHNI5/oXSOy9V3ukHMSBk37rd4RIxJVSjybHien0Vi7plncx+oAmR3SnkD7piXL4
UjL0i8qFQipRYW/mBg9Kzug1fuPD4AO9tNnPbMWKNd5kZkSGA9x+bVZ67kX7xxjrU7U2PYBTKz4m
poz+Pjac6HGmiz9zYdbPSAbpgD1cRFLUQdO2zjqVOJQdu5kCydc8ZIJFiJKdh64rsSYMkqnfp4sz
VzbrMGDZ6YWDCbCPkXGPf9FnCi66Rt5Rgrybd8Cc+J9fXVlbh7s9sG9hrxnbYQK60eGrScHSv69l
g8Npt6qo1Ufx9fFHcHEKmHs0PurQycnToKqvNjUcctDn7tsdLEWt8FlyOLHe5A+iSR+L8gvtk35G
cBbcFeoipd10ULQcNjqSux0kh8WShf+GKbJSxd/yNnuqfA9v9BLDH2bh58d5iuK33FAmto6m7ZBU
jSeUILbk43xmb3NXN0jQ87rAlVrD3tmr6Aj3Q8XeUDr8he+WHKaYDvM/QRIuJWC2C+hhaVmIgn9m
BbTJH5JcyocSX0WE49KMJLn17PhPEnvtfyRre69aNr0uFkbtfrByX1m+wNDiKW8fV+7P2FPJ0bNF
u/U4wSFEZzdqSAoRzzLduB0oAHkY119Jgo+16xAnf8CLFyWvKz2m6pXEuH3ziggyigjEwfTWJUS4
nAmxjFOG7U7Hi3MTTWN/S2H9HOEdQhCNwupQnfVCAuqy+UtT0z4N7vNypkYdFYJYl6vKA3dvl3QQ
D/tmmGbKPa9ApZQqFYB9i/1/sI7TKi7Jv5KcYhwBSyTcZKnfe4Sc0FjTRP53amL7eToMehg42ixe
z74mLGEsPVRGjfxdNSxQ71EVPj4DrMiE9ou6dB2w3pxChDL/HCvU+GD0ZS9GU7WEDRYYiUoRmkTI
t4ri50b5QI28gYt/B6tAau2wgjUzSqCU8mNCdWxgWkI7Kxe1nKrEUUy70RM9+CWPzbFALIFQALSD
kXpTmatRNNur5GP/Tj3HQMdN2TwRYSkilp5GT7vX8J6I6hJ74eTAfyv7NvxiwG/K03OUbavs7Z+3
DRnolI0DItatiGzqkJzREK2uKVuU9uDv/z657MHAomJa68ls7SmZOzxDlF813qgxtNEVN8zTOyz5
OCyoFwf2/kMuKVrP/iDZhOyjiZRq3WBlYdRvFx0oGC4CA6SFG/YdQ5X3uo3tWX4kgWbnCGX3ms6Y
NdD3P19gwig+w6CM5qCbcobnxzycYdWjqJpeV/kjD5Y6vbTJXEzHmMFJTtOfVOaqNVfv3D57J+eg
Lr6te0bJYglXt90o7js780RFxHvkppPIWIfIKXLEUBc8Boj9hLtfao1j2WlAV7A1bHoGqOSX0IIP
32aAr6f8zwbJ9Qq0G45zsTEiIn4pZE+kc6MX2mRy0aijXSOP8AKIkV7e7zb/J1lSRoz3HKuGuw2y
fbjkHATwsIPqRGupCvo5lVCj47OpeGwv3ZgKaXElEL8r5FyYV9ILgoKQsOOJIXj3vEBvTu6qkWSy
QMn1hswhNUsCsTXyCNbRN//NXv5x/CXtehv14RO4ZIlWIQeT67NQB5FSCUiibYEhYpFjDIaDyi2A
FxGdBCbhk0049cpAwzvguRl7MpWscJicXLHgzj7LoIFEnTrP4ueaj/q90iHXO3ieL+FRKEB4Yzi3
NMK7K99RvhN5w8bEAqY6hs8Frw4rYqmEwfoNIACIjz0IKzeiZfAXwV2f0qbQaTRSEIOE2Ns77jEJ
4R6k1MZAYzm/nBc10do9p1bap7wrf37prMKt5xxiVV1o53O1/rUR/Jj7FTZJ7NbqSWoDQTyUFe4g
gmdTxcBryhCj0YHqSOlJliN0isWDILN/RYdAkOgBiqV/tU0Ddw01bJ9lvjYzrHSQBA/Ljo8H6HfB
E0YcsJMKsNIuocS0TdoQa00NWkLKhbzbA108Ns5x5DJTkuzxuW0tDkrQwIybkvpYl0osVmaPdD7s
M8wWyTJGTfG/q0DiaurCUJ33K0yzmxBFKWdg1WXJcjHm6VHJnLsQKyvrP+TOX/cBxfr2Z3MQI+6t
haAz3H8/TC31ZuGRrqPk6ZIYSzs5htPP6qGHO5XbT5fGMigAMn0JSM4UQMIpxYZi+8a/s3jGGoW6
LsgXMTtWYJc5p7rfBYGI0/ZKSi7ns9S8Ble0oHiA71+hEp2Lr6iVzWWqZRbhFvUCdgfabGX5DR1j
n/l2kjD+Q+L/jtJMYwVKIv4XX8moZvt/5i7WplUrw4Zjw4LrVQW2RMC+udXpOrzM2WaxElJvirr3
ojGS1JETdGtWiFGaZYreBWniVhbKV6Mj5iDNA69uaxciSTfwOV2rNvKwqClSjAnqvATelr3swCUp
zpANpiWMhQZVjMpaNjqaBjU34/64okJC8PztMYy6kOVQheUjxuaSLRTGTcG+XrPllfuROzRRLTMI
+w589iYJnyavgf6HRvNKAYBtwQlIMCRHztpBhHk2DrtaiAfKluigIw8J31hXXJm9h0RvdjxtD7UM
/tycjxofpo1ltWkfrSsI4DMpu3NHJFIkM2EAOWdfD7SWZi1D6Ygy5Ej9xpJ5HMo56cVuT8SMxu/i
DHNprzu3KB8gnw6nfLm61vOZ4Nt5J6YkmefqtCcjs8DXvfOWtFPfgkOKgMPL88jlQTTxXKRNScTL
b6THG4oqVDNAI2BPWyTrHhxgyhl901npA/0PNu0DMjb/6ktzRDjapYN/OlXSgaJlrWWup+am5xLN
mFO5WkJ5VvUDeH47BsG/Z1FrJa6KdncZq67Zi2f4iKdjNa7o06dm2xD3zh+XeVFDnV+1RuDpeMwO
1z/IgeEzZH+PrZYOgPdwKOPL8LdubpatRf0rOnrAinRa9BYxI4iOqiG4JVgovsWhV8mgrDdELiDP
TT6K8+ZKCsKpWwll2nYwwQrdzHWl0oaGDXYxjgpH7w9fMrW1bxYGKBCNq+8fonea5bJyLMjJKGUD
UvohBv0wCbpCsBco0bYXbEsiQuGcPziVLrOUezIOpAVXs8mW1gzgiw72i3Z4V/tueSen64KWOc5d
puZ72yTUfhXDRWMINYLjKA4gt6wUoq3854uPqLBPR/V18HnvGaPKLJyFIG6swdj1g5VP9cTQK0JL
vvAuF65aFNYb2fNLi2Rn/vEzCPz2XLQNM2/2OQlMLK48HwwImarv8nqoJV1SIEyLV4cH9ht6S5YE
Z9tQwwVv1BSUOXpJH17vQcjI6k2FdjLMYNrM1KzmKE8zum3mmsAuwvcXaD3TX40nmY2/rbbxUSef
lpSNFLvf/Lcaz3Rr0l3ikv1rczf4FCdT6kBRk1Nb9oHj8tkVUASn69R0+Ui0GrlFBjGkW4tKe4D8
AIw9MumxSrQXILmQEQc2nZQsfTZ2B9V5F2RMnoW3JzbT/KN5+L34kbru9BXQtKsIsFBUjI8BBCNS
ZLC6QSkqRS0F0oOiIyY8TlIVwUGBi+TE0YZVnp3IFORvM7eIdiurc2owu/FGqmgUbJoPqDmBnlI+
7S4TE44jLrGORa2hWwg8KBbjvQfyQTJOACNJzdZNC+fhwAk7SJUUgPDf5WdmwK+LlPFi1QuSYfwM
6b0ld6o540CiWC4wg/nUY8N8kT0H3m/jiXO8pi2Lh0MnS96Ujyb6P3KIO+CaudThBXAnZvOEAmXy
w8ma42m2jtGW5Ox2LW2Aj+bg+1g7zRo5rZUhBitM/aWll+9wJzQMVaRPglrGcJVMU4UKMoyMwHtl
sEK38Zid+qCBCKfYt3VVqNFKhr+TnL6M7EG7ATWe+mGugPdkwTXKQR8bYgMuX8V4gbuE74zBB5CD
Tw6iFckVTK8qAXGxL7Encv1oXt5adA+PFJ4Ud2DLOJl3AkbUmEq4OdimNdh17qsLEdSqEQiCC4Jy
tSQjbrOInz+RZ8mNmEpN181Ux9l5LiR96+PHuoLzG3FIPK6cEljfFeMV1p4ax8i7GqZS0Kt2/cGu
AUaCnQklwTY3WSIKkWOm0ob/ejILMARnm3XJ9LmCe3NgJ4ZKgqIzHNTM6XdV+GkmkeQJaXbNkZhR
v5esi5OUrelQS1GZqGGjdqheDm4nBhd+y7SqZgg4UntH9/xUQA+lEZG9+SxauY3/SA2VXnFkIbTM
7PENEFtHJO6olPQJbq5NFoY8rWc9f68cLOfqmXsjGLhOCkw4jUsPSHwaEafl2N/WYPk6Z5FNg/6F
tMgBd4iU4pA7j3h8ELdIsID0dBtKJZAL5t3HZc8wB3t4CuIPXZ08SpnZ1A57t6BH9t+S4DhhVLxE
2AQZFF0P8gdd5fHZMb/Zp/eGMDc0gN+VaAZq6C2TBMdBIGg99XjFRSpELhsJ0ICRuv+iEFWvrd4+
zZIpo359BhFywPLoUxxvZGcsQ8HORIfZdWqgOGtC3xqwWtnOJeAW43lQh+CBWXVyakzWaZ7/5CPG
P4F+35fmVEuBDac/03YPHRB5BUtlGBtc/wAqKW1YFL8iiS6C/8HEaVUNwr3wnwR3ovEK/ptPddB5
xJZRw0Oqj4TS6LdRKH0w1ZNJsrDEefFWQ504kivWoWC5PMa2cwsJ13cLUKYu/cBFjV7aYGMeE6VI
OoLsJe9zNHnkh0gJlcg15sGQKJtuojWsz3T3976FJU8qHBp1jYbAfz/wXwKC7a51VrsV0rHZPW36
TUzO/50VhB4ldFSq5AEF+5qT1y3NmDRWsNOHV1w77oxGWgU5Q40pKftTUi65qB2KpHZ/3BeydnyT
49oPFIhF5sUs32v64kjSPSqYtwWRDuCO1cYxjCr6Go7xgZkt4lPaUWhyAsE9DcnHkSCuOaPi8c4k
XwCLp5QwtTOkB+OWmBqzVxmn4sa88t2Tl2RB2ZgU03LHEnZ7um7K+8Zk8zTgq7GQo9Rlc6uxkqsp
TG277GrlZEH++Z95/OwWUuiB3NJI36/MfobvdZ5SsfGUBsN6NHee5PZdtar3uVLjLsrWVFg9BlCj
TiYziSbUVOpNdiV+ZE5lTcOYao0JB1+RZD73n6WlwjChJf27J0QGWwe9OMfA6RGHATrUh2DS88Va
jnoJyISR3OCDqtfFyVMNarnrMZVBj4RJuyJZIgQQbRXyEVA/aCz4XZYT7CwKcoEhNdwlfmTj7gOV
BdNUA33Kr4dc54QwOdM4XXgO8Xfkjq8tyiIwwiMHGdBQ2XCCbkgSWWGtJUb9Mq7yUc0kmogkF+eh
pRbR9TXzzS+7ZO8+62Z/pKPx5OVv1CmqJsur2Bf6AH9dUB/ILptBzVaIVRGcKO/URbK5NsD6mjvk
vyEmHOsFUmC7vaFM/GE+pE2nIGeyAYoBdoyGaB3Gntbe1VB9pZsWp7F5MlcqdCyogW3xGwuZ/Ky7
gqqQn4SpAYyEfUN6MBjYbugmErbVHG3n8D+b6mMfm/weH5B7bZ9/poxy5XYWn46eXAjyMxeyf4fX
lD1ttca0EXasmu8Qx+s1k9yjhCFuRYI5+6Qmfu1GPVHuKvvKSejey+j6hUZgPNkY8fbmmXk9Uq9W
kQV+a3XZOhKznrYtqiMeUnD+x/Wy2fjCSxxNln3YPEHDDPT7ufRKV7MvO6h7dkkla2/iEAkXeJzI
BvgEY7M/rPK62I9pGjpb0GqkR8lNPVBLUuv2mp/vRhld+GjWaOB01+1+Sark7qxz6lJ8M6xaWN4H
wSPAirpqLbwkaqRUpKm66y+IFOhOZ41VBNDoMWaxciPrHybPsx1xj3QzLnpmzEyqccIya0+4k9oH
UGRv5mZsGxHkAJ0effmIS8VTuXtQ5w3aVAIlv2j3y+1fO82rnJS4ejj1kXv5oAN4xCqRy0+6nRx1
a1Ytbk8aq3bJemqBjMwI/N3hZovd2W3co7gQ47H6mAiYuoD05rOCRDilGyQwaL1JZGUkAJmKP+2I
FYsHksQVnhDx0zqqbT4/49LJVCGXkhFyE/Oyu2VTk8iLOFLiQHBWqRnOl3wONrltEJza6dt5mHhc
bAkemZdwgHERlVvNP74eoGOJyXdp4bYk8dqTpllL3B2O/p/wCji4RKU9PxnQFUe/3AnukyGw1wi5
I/KFUvaDwr1AE/X9xV4m8vEqDFPvMa49ljyI4Rs9OywbPnjr/1nYLqtGiRfIc76dwiPoqNas7564
8DmyCYKOg3uVt1mszja5CNU5CsNoe6/eeg1WupEOy8hksHWJ5XjKok8bhUZjW0bvfiEpenFIYHFb
7AMXbbApBAayQW5llbKVMvBTWv0+KIj+xh4bDJjXeY4gG200Fxu2deIgVxgUyzrZVUUTk/6aJURW
tSPhCLN1emesRAQGiBqHhNBCIjadiUBW/BuRMpeYyihxjoejuju1cxbqwWOuqmuouN1XIoztSod/
u8XzecoB9ZppFpJVtnvlL2YuZ/5Ys80/U4IflE/ov565OWzv2MVGURUR6mKgZaBcxc6k6jWosUms
Skxbgy52Q9KwaBnWq5fW46dmo4wJaBivF3jQ2MOAaFlxGDWkMEYNBfziiqJssGXfg29uRbQ7fFJI
v8gjBDqaDLMu1d7EZD58LufCz8KQ5pjGWmIxEgKl+0r4ujggkKPBMjTefdOEVt6DCiJeCs2a7GJl
M/Ypg7T712aB8pz+1URfKOEzpizl1sk4FOqvQnJNKZUMphscMy6dR0j530ptNSNb1HjkJTIbuUOF
H85erCfWM/qnnwt+v1OB9GVqy+Y2HXx7GCtNDl2Orht2WPWAhdRs7FuTyIdBntVnTip27eRX4WTp
MRHnxsxpv8KiJu/4gVNm6lVnKeHk5qrYbb18uwk0/KZlFHDPO2kK2pLQP5LsUo2yD4g9jZSZUgPS
vziFCH8aGU0KloLNb278VoDg3O/KaQOjQnbhjv0RU8/+4QjkqZ14OVpf2RBugKXEB3x6yMlVj6z5
1bA7GLpCZx/oTLCIDorKjFW+ys9KivZxQ+CIyybtSBdoXqtJTNs9Sv6dSttJJzWGqzNyr0aoRPaj
BkfXNOHEff6hirFirNBRN+eJ92HGhIUN7gBGn8/6NWhdEsRGcdmlP0vKP6lhhD8gwrB1HPSiPpdg
MBaL638Ao6Pqjz1mRR1fOKivGGODFzBzlQuOt3CwWgSG/Q73jOsIZNWHze5QAeXrPU5kb5XaRvEc
id4uWQvwW/aeSgy0eZ2kllrc+De3qGy628hpqRcNp+saKJ1PIjJqVu/ru4/L9GCfpVF6HQBhHHDz
oPo9X8fCyfFUTgky57TEDAP8MnVxs+/5GwSaLa1QZh+OfohxKDZKPPx/g1vrX7wrV+e0t9e1nrJp
yGD+Qs5aMNSOVuVXTs+/NAXC0qSWoaCdV0zN/Y1leI4SWFx8FE76VSpd6aTuxDwvLp9uXDcsUEXW
bU4tnK3lKmE7/+Uo/s92hRPfKtY33Q0MzMRIg1rtMtgx+2OkTHRBSCXMwy2/+LHcIsWwdYIAGGBL
sWy8TRmY5f+Pn8oQR6P/dD/FVk7+s3ep7/UWvP2qHOeucpaTDPVSHqOIghf5WEF4cFN5paRWc4a3
MESu9LuWnc17sAt1bRtsVmBO+6MyKxo9SJQT5ocW6kS7qkX/AvtZOfp9byayseALWiv2lTXOYpd0
xwH/Varhb9F0C+1nnqCqulI+OVZbSLWOvYIqzXIwv+HvF0trW3QLXT/ZMecAvnKV97MfEr+kj0ZR
Id0WRsU110I56lNsDTl+HplFgtyJd5TjlxDmicv1Agnjsjrqvh8QypZo2ZZNveHgD5jrlar+NbAi
NcUvPg0NPodiEjD2IkkRj5eSKLPTHsOEFXY0Y2TiJnWfTt6WuPFu+R0Z7Z10vE0xIpVZG6JiHmLT
O0KNXJgQy+n82TME0NUTqQ9VphptUui62GA50OwtwhhGwsHRCxAcCr0ZpRRFYSoqUfeyarCWZF0T
dkz69PCSIveRFOHuvgu2PG/KimuOtxrb0fkG3610TX8OL5ITIYbETJTK6Od/oQchdR2XADk/zk68
QKrtExeKMpxc0ne5iuRkFgO9tiP0z0eXxYWsAqRCNvYHi9snk/ypYG00R3RYn0H0cio64OvzIC4y
zE1hnGmD26UBhC378u3SOhxPESMQN0S1eHxNQ29eTmCATgka7umsIai8JnEosSJFVpdXrkBZ65eT
Bkt7su9VBpYwOsK7pANVohCSdpVOREHbvp9YzZfDjxe+LAuKNcfNXKanwXddbzBN0uYAdofcsirv
q1qHMGhJ47E+udtP6sZzyGefoDLL45h5mrUb8PP/CUtoEl0XVVbfXHA6b4PuML2PayTWQyBRsDbn
3GvaH8xqhZgwDHlYJzMufWouclpjOb6CBqbpmQjqqQYvmM3hPoEOBGlcvve9USADjTyGNHPvSvtp
0NLbxiowxMzGO1ittunVZODKKhSVrU/RAoIMoWPSHp54Ga5ZNoRq4W1kwKlM1/G53GnHYDOM/mLY
AngIFt7WZZOZVVEEq2In9PlTpad8OWHSLtE0UMmUW2GoZzQ8abXT9+XFQGdNvnJmCSjcgfDU0I0n
3Nvx1skMSont7HPFek/1iFiRJox3jCYIz44jYLfk3K130Zr3fDU1o1zbu3e2ECCvoVPKM7ELgMC0
MknH+jy9ti3XYA08U756dD9sIpafWJ7ULW+rgxN+m5V7lSts7vO99v475ckbA3ut+Hbsec1RpgoD
UnLdg5qj+2U7WgwLXP2D24SYHDCUTokz15W4+JspYWKsESjXYeJeSN9c1+ZMY2YFvPWAR7WP6Ozs
DOGAZJ1bSiLouZLZRSpaxh7xU2TSrVskQBhkMrU+cBo3qAxM8yGAdRGeMHVGcxm6A8AhAddHQiHB
jIKzbHD36P95vaqdUm5pa7j8T07TrmhbgCMGZFrDqz6+ZdpGkhpLL/UWVrFeEZMIdaQrUJtWYEse
7clVbz4n86OhlALCrZijsEZNroInkIK9BAis8F8c4VgsBjP7t0XP9ueAmxqUbqDn64rG3EyTQt+2
qR/gNZ93EyhJRAyJzF7SC74dyoOyhbQsF5DItGZQWQQjQo9IXYh88vCACvHPYtz3n0cax1um2ZWs
EFZ8Pv4cMD+bQ6OcX+o4cM+Ph6LpyW07TS+6tNnHhYOc60MTHSYSs9xDw0qmpwRSZjcIrhhXj/QR
/NY/lrdk0onmF5w79pQjR+tFXiEQShVMeQXLg6ElQed+KVLnd4G7Q2Q5sGOYk4Lg5xLh9Wm57Co5
/9QUpu0vIJ5fpWJIZ0Fw4Yxpa55FEXyjal0ooZlcGFvyP5QrhiJhXfN2R6VaQKEvBIjJS0dNoW2Q
jIXO4Z+L3x6wduFg7/bKxFTm+pp+14htl3Q/RIXEAwIInsvASBtk9UGmRfYCWvJLjktz5o6Kpo9t
JHJ9WFy8dG47aAQ9Q9wVN6Ku2dmMc0vg5Kek5da07RD5OZTzj4i64qWjKE5syhZU+rIS5GtJlvQv
lBl+K+Wv5Pc43VbQ/nEz/jenKdyeKV1CCAaP3ZFCOi3lTjK0/gz3x+2zoocvmkZQP6HlXVGsM0KL
92crELvT3fi9DBxi3N9doX5C/VaZLFKF/Q6rcLy/Tw8apaSMKgM8gJ6Fe/wieFoK4yBjJ/MvzHc0
8pkYB4o0oHVkk+tljJxpUcLMoSK0UUZPUo81t9UAfGJgrBFnRsZxBANUFRaw+MmZnVEcSMeNy0bZ
n1YkqW7VXqMcq1/mDrWfST45bVtzGKf8Jxi8xhQTFg2gLEh5jZkeDZcBbYtfNU+ELna+qit2UOAs
SO80MhnglThosZ8LLm3XSuWWICiQCGzdsArhwlf8J7r837BjS6WcnL5pglTXEk9ZY6wmCE+UJ/lC
4yXwLEpHNTcD+mcXQ3MEcrm8yNgaAYJ7NwQgyEFi5JQE2LjHG1GuR7L/A5CSUXLnv1c7mKYij+zT
/YQmedchLYaIrUj+xdi3HWJQT1JnUsADz/O13X/xJJC2nRpaBWsag+59kWrIa8WhqOpWu558/6c7
eGZBVEDSJPiCtJczlyzprc+vsbbuG9JdYz/yWOPMMxTArV1+ykdYWSP9o2gB3Bjbw1+MFz0VLOAk
RnL7dh/K8BMfa45QyfqlHD278H0iIQxtdVHhX+0na6o+FNmQEYATJsdPyMCADYqf2tfiuCYICTDU
nDw9Ixh+KAF5KVGaGwhL3vKzX0DyrAoGE/Vyr/mrTbuo5WLNqbBTAPejjNG8XKmkie/WYd6Gamds
z/EpiFCq90pkWmOyCQdRfTzz516LRFkqGw0tcRd69B+KFSIs/6W4pcV9IZIHQz8auKtrki/5sfRI
5n8YCwWR3e9ugaI29owfhncP2U4K0G0DQYzydBGSrdAwVkJb2YiPUJcERrFkqG09SEv/IJBoK0tW
XUendpRhHrd7TPwtcdnfoPe48WOvYR2XqfJAMbvLuKZL5wkrZCo+bHsCs3olt3t54/vwWrbfg2Yu
OOUHqAN81MEBzfFek/HFSFEjtw07R+GbjBUMtD7f9PZjf6UZpR/GOof6Jed521D1l9Ii41Y6Rfti
ivend9FQ8jzjBXn/UX0yI9BXRiV40U5eJYT1QvCcBmxx5ciiDpDNo/Yk6jV3E80GF4l/Y9FM9MQJ
jjrZjLa+ziFjxultjPBsMZZusDA+74AxmTm7AiN6IvhcXgOJgNbUifCHWGtsMJkncSIZvtMGgKiQ
oHefiZVG8JUh68KKPP1bD9gOp/nnHROu/eE+Fz4h/hqfp9FMM92g4NFA25EMMgqOnUxLczPgMuQx
amEzWsSLPL3Qr7gP6IGJWAB5gVgs+RBwYdLx+p5ZUpxcWLt/L/wKWkFtEpbOf0tpss7Z5OReYHBK
wAyIgPANW9RpU9ABZhlzR6cCsyEo+a97zhkXpkzjJJV2DQNbUAuPsJDiO/dVW4t03u5WybbQsHmm
K/O7fhQ1CoJeA6SkYv/anm2LkqIPuMRzj44xBeY7aPKGdKCdDi3ZIgGG/KlDzqd3KhsCbIwaHozz
w/uRE94OeCdheRndG3eaXJoVwPSiHBwq+VJo9R7iFVVYBGC8tsFJbuwrBWG9ztBjT8x5qn00DDqG
s83+ysqBO9Vby3r+OgQ+H3GTxNVVK4hkmhn9hyE90HpNtQPyklZR7weYZ0QB5sbLFGZES/kOwI+E
fAeQzr/Itl5Q1HhzaDa2N5XCLsLRH+OPFrfOOZ3/o+0Mdmb7sh9VP3ZLB1/LPWVXvLYGo58UjyPl
lSXcEerUDrJD6m8ZeNcWSMHF09n5ZeKK8RkZYO1SfD3B5lYBVJFxIBiusuXG8oNR6IMAPL88fp+U
tQeccmDi2hbHmPzx6InTMtSQVlJWzp2xJcXMbFMEwOrfgsniskfKVPNeXR/xQTWGydbJnKGKvcy9
YU81AdZRIoiQcRsEvVNY3tZ4K+5Sn38CJqROZyMh+JMfcXOFw4TeGeaYX1b6R60QBW1fUvEKENGZ
wGfAxbj0naO7NkBdsYXjBj44Q6D5fxkcvXOqfTAN1BWrmTEdRNBMILkvgZmI2j0YvAwDu1gwRqvA
WX9JGKBwi2F4uE5lh+jWPKHu7Pl6zTRtG0A3pA0BqwQDOjJrvhNisnVnC4yWGeM8kdEwNur5/pCq
QWv8kJrRK5pKcN+J9MI3j1U8wdrZzOGTImAZyTsMC2qZa+9qUd2EpP4LZesUrLYVZiTTVUVoHLqL
DroQWbLWiDMrhQ+J4IDPjJ/EwIRQiavMW55meU/H5ZwB9S4jO/bvB0V30VhD4afWnuz1YkVeD9Zf
qDsRH8B/qTF5wu4u+8QIb7eQcEoGeeBo2Exp7k1j9RLt4R4sSB2P8KGd/zGilhnvVH+B/fbHT9C/
De/OaVAsWdcGd8bpLoNJjc9Pm6WPZUE2BdTTKSuBEyR5gkF0ZRh+tlOT+J3SxEyQ0IzXhp3rTjj5
gcNe9iBYe9oxZbP+CPIkbxmbC7DWC3gsF5l4MpGMwGzT8Ehwuj8vLFwAuAw5377M72iSTUd7CWsK
E3cObwjHVcDgikGWbjPbaVjLgMJZADeMz5jFSInETomC+DZY7QHqRwViVEVjKKWogz7TbwHZ/kvA
t2yPSbZH6gIJRYazg7nwOUXiTrdpC3Nd6xCHS2MAoNDjclaZMkvn/5AmHdSTEIpUqb9mkIwgK2t9
8Teq/E2pOQFDE+g083IGto+RPNpHXKwqIhDcB3Mjn526KSWJKaseyG80gp4v9Gb5SBZs1d+amenj
oZTFTT7nrejvrRe9Rq9meRcG3p6ozsUpRvHpNbq1hNqxaYpLF4+1eQdbdm7LwyGPvY4X9PEMoKSm
4tm5/QUwGn0Qm+XU9i9uLpkRPZOyM4wpiXQlKTyrB+YnQp6lJ89iKXdWpQm3BNF5LNIBLlz5EKS3
sx6fDo/vlkj5p2fm+Eg7i1eLsFzjeMTLzF8hVjP9XRZVyAhO1NmyMcZJiJo1Rw1pMRwerfVquj/b
0QqhvWlaIQj+lEw8eqtxmC3jNDzeRCOJrUsrCNvm77B0o72Zw0katuIgLspZj/Qh/Rhn+2jvYwXR
bXjkwlnNQuYcDEDaIJwP4g5yy0Yz5vRdyIOwd727XTC1gNWeRKtGHWCiw0qdO485YKRLdcWG9bU4
wUEGQn4xQc7WBfNEAeSZctuYUTzKfj9f59fMJwIZg2AMKom7psO1pC24WcK3Zy6Nbo6iyaAT+KiN
zQnDHsPdkGy1KO59Iu1zBccLjWUi+3/NvxpuelX9dJ2Kx4jq/+ibGFFzI6N903DodRZdRU3+niGq
CDEkW1MFUcbnP8cbmAJtNHCBwaoej3hmaVukdg0Zy+cxqnM70NNCxT/zkSAYepFo0MdpSA6KaZNJ
iNmCSncHiUj2uqV1oZQwKQzFSLG0MRUUgNX6m4dahSTQlSXSCfEKpppXw4BQEHkVfcKtPt2pb+V6
jVmhqJB7vmUk6mqVpYPc20bVrK4nnSnkEtR3e5EPged91X6gTY+O7UF3x5qP7ND3XKB47EwByan6
YmK0clzGcuPaNn9HLkz5Eedc0UaF4L59ERJPR/+SUXLKWTrNRi5f6uKxgobrATZJH3JsWJckgXfT
YF7Dyf/K9I6gnMp6iMBX1aW4LHvYm7S7DDLdAxycytjo4tbNFbEyyGvbkF6jtK6NuXaZ2ir6nixV
ZW/erZAIuP4iDut4+6yhCHs1vuDcCIU1E/cpEH8nwUpbCG0K31a4c6nhG7raNZnVuux0kj6dsHKL
ulJi2Rz0yLoGDZXFUbZ3/H9OayIMN0u1ECjxGtTNaGZ6fQYsPpvUX1Mgb0Sxn3pcIfxeaeL9M/Bf
qnsO8CNKqwocUVcKiWB0t8p/uW89buL7Z0GFdh3R8HzXNcs85PJPFh7PzoOuNm59oT08NpVwGttN
5pXoN0e/dDNmWNsfSS+y9nvVtWjh8p2vFKpwrONElGbK3dM5VQJlI59nZShmn07KnqvLfSo+VbO/
qNwRt0EL4/AJVHGlbuxPMYKwYkgMk7IX5DyE6I6GgwN5lUuz03+ex6jTPv56KAqaioX+5uMEZS0n
aOn0gBaSGbKBefUtc5X1dFO5gAid9WMjdbs4ALKAwgwSYdFD13OJ2PW42y4hy4OVUNz+znVHUTVi
X+k/Us0MMgkR8D1UAP5dC8x1+w0dvd361vLs1LTnzHLdztLfSsljKsCWz7Oxjlc6Vb/GdrhGJl44
4uIGYIrXFE8gSmhsKL6RH3qtmXEV6KBiTeWIqr0Gkg8BDkA6H9aCNN+4/XMWujjjd6KijaNSWQhe
zz7QTuWYrz6Nd5+/maQGpXj2RJgY9KU+kKQpn2KkI654Pumw2YalXaFqyiOMjVGEV9h7Yy5EGgFf
X0anXUM93dvQlNU5M4v/SiFndo2r9Wdf7wp2xpPRGaA3kYQJAyYCjV3cIvNQlxfiJCGhZR/5oBVD
lKcs5VWujgN7BFcrjWSclA5WVlEbSlxBclMtyfXflhj+x/Cak67WM9yJsVotxfnWoISQJUnegYJl
jSuBRpjgdJnp5tcCYmE1ywnLpRLn3G6sHM4bZhPD6eduEZhvQ4605AhIY3ZUBI3bAbEKJh1D2xI7
3ZBPBGdkdmWY81uxdeVTMxqvmNp/ng47BBP7caCQO8nswE5A/xy5YumFZbAD/0AiGmNFBkD06Eyv
9xdDOHdMmRxGcbSC1AZZDEmzlOJSs+mpPI4QnG+s7mQ/IgaanscU/xl4MA/tXwWFkgCVgxOuNvhz
5pyVXZ5vfzM6XK5GKZFV8QK6ErcEW2K3YIJHpvewX2xeglYuelZNWmjgGP+sJTUWaEAoKmdUO3iH
abJyFbUfbu+ATXu9nfhUp5fPPzrB8Vm8haQ0FN4LPhcWerYcYMcUmtiCkaU1EKThl8OyxG/CWtxJ
NVSXmg/v1TZa4sE9YS8DCyDY9myLKds8+gUtlP/EoOLA0W0b7ju4aFf40kg+v8IL1w4woILuSvBz
P+TPUhFzAvdcHfsI4+wJi7DMuRika+YLfAIg+B+ArJWajRTEwm91zgV+Tim66udGnZmhU5bCKE29
CkKfs2d7bz162nISabtfm8DB5laHZwhrdboQEKrMhNgAEBL6IJO3/8K3yyvspR/P8JRWSdeBBF2q
d/vyVGK+JTg4VkRFjxKlcMlgnfSKx90gCL3Mu82JjdJMXP/664WECmWK+TwomTFtk9ORJRGOJ51p
fiFKREa8Y4XQt/qtBnSiP8tlk+OieYlH+f3dyvFWIn65F6F+Au5QgVHxvAMoh61yTUZvWeAVzdcN
FjBQBPJGeg9RD8qv+jEU35cUSXudj7v2D0RiW9XYH5daXVRERjc8PeRgcb7XRr1hoV3uwr/fyAAw
t/Lj5c6T1jeK0J1kdnKOTlln1NGX83Ow1o8wsGJJc+DczLCeA+czqQQWS3ADvy6hkPAz+i5v9O8G
cp27NS5JY77Z+jsQSTpKs87SBwkeCP5+XqnfroAUMWwFNUT8YxDklNilCAsuSk7y2Joj+78TlR88
yqX6Z+h2DQ7yUg0qppQ8+ScXY/sX25uilmvmK+E8L/SSXFVhw9qnNFFY0GQTlNwYLC9qwa1Iqa4q
5jKrehH2Q6oDINV1FU3D4pdaJ3VD8LcIBFgls4JwId9n3iq5OM0UftoaoTwJOUDO21Z8B2nbVd3y
7DGCRl39g14Ig/qK1ISpwnHblpJQeDbC09SYrI4smIAakuFiDfZPgptNuZo0I+RjnFFUAG1ur5kQ
aD2W/WNfTxBOu772TG0P1HQ6RjvFAJITOxT3g3yhDDYwW9pvrEGGZgZzEXY+dbPT+345zLQBuGb6
PadfnjiZ3VdhJxGPu8nUh1kX1hJ1Dfi7ezBbdOftHFf0qMuUu/TPsjLBdkUFJ1vzFBNTv0mn4fXv
JijvqlZ9Al8QJwzR1yfukW9Ao/73CiUzWaXWkATSnVTd6HwCWCNP8vsjTi2Kkldbtobz4ALf+bOC
NsgGJXB+8eVirrTCEoo1UL4KCP+3NlJ4NFqSfsxe+zEdj8lSfPZsPrRzYYaTC16AnxEXzuwVjHLi
6Fabv/P/wwt6YDgtVk5xdLz8v5XSkfJqT31qGmZGLaAqh5fGEiyDS3iF3hGB3wm4io7crscyIpQj
9hA2SooyNlid4VXJLuMwCSqNJ4YTLr/xl1NIjGr5k0CbIwing1vMzV3SgQ/UHtUPiG7hzD0lZ1Rd
6nv15lMoFkREEg/pv19dE23HBAyQvcYYnFhlO6qXSL2ySvRK8LxHnZ2uVCXTUraJ0sblwCaSKBDp
VjT/o6AXcKjARl/qI8R3Owi6V2EFgMdh4IYkR5Aq5qsQ8VO9fvszvwnXZEJSaAXlujNCC3vHKxT5
6Oct9gRNirXTNzLbku6k8/3kGco6gJ2jFsOWpv9OAIgiHhMy2gHVvBVh4nAtYPkNBBGpJSDFzYbg
f27RxwJ/L1mfm9Ec08cyQ29DGHgxhgovV2DyjFNPGcSD3ewu21kDEuSTGj4qDZf2HbgmHqQsO+XX
imgvvg6BS8nQ6/n9GOfV5xujnuWKocTjjNVqjK7TxruARdSz7rbPn0CmQVHiKnRBSg46aipprMJR
94hlPPRwbKGT5vX/Iz1yCsK04aEBLu73SZvT+UzPUFROi/Ju8Fby8EbQHXeIWrmYD1sQ7H1AVea0
qGa9F6sBW6o9T9kFylDBkdPIbfVleDx0dQeBxHI7LDjMSwvzeeIybNe17y4V+GreDtCkBh98ymEd
zSP6clf9lR3ql3QYdeMjRbK0+s+3wMOXtz2mN0XE1dHDTeMxeRNQHW+brm3MpSnnJDM613E/WIa+
ylttOC8/lTzuIOOdY8WTd9PwJrpCKsFOf9Pc75GMzQW+7VpMOuxRoQV9srIH9NcnqrEVxFZ9Cfn6
YU7CA2uz8YPa40pvmfXFl8oemoGDe+9uG5+0nRJDeynOBDHu7/eCmYa0li3/XbFqQ6vdy6IYiBl3
95iWDHawsBNnQFLvBMj4+lr3CMWRhe42RH1pL7NhkV8k1wOGOuGsj4rJ/kiYUa+2Zn0J2xH8xL2A
aHZSaBkmzwZCSGPfc50CDUdOpPy4bOWAINp+BNLlhbYa0dZJ0Gg6yjhDYWq+Wkz65o2NDkg9EuYP
Ss1+BEJEauCjcw+i0KAGoEOOtz6B4rRfpvACyO5PIOp5MN2lyT5CxF+UIyyIQ1wBYGaSvC8DR+vN
nt7jXBw5oDRL3GDtO5WPqBvhm1tWReu+7AV1tMDE6lug1RuMVpt7LYXpxMBdA4OAt3R78Vk/529N
QkiSR2W0FAk5ZSXHlYcnCo1qf8xw0K2cHnWkPKwhOfddPAPvvyjXj5gXe2l0cQ++LFBFWdoLcsZZ
5ca30jQoBnbliK7OL7CbX4pq0NYE/R1HGhPvdqK6w3EPjeO6BWdg4xn7CDZZa/bgHK2xZddyDTbC
D6F9H+EVtHoMurPVhDmXeHylOrCCygtnH0wRXCTFkRY7EIva4l0MHK7ktSRNMHxPA5ZYlOdcfcNK
8qkSDCOEH8W8SCjPCqY0YhVE7z9gMg72OHaT15eO35Yvj1m7R+g5GTEYPp+1iJ5rVuunjfTX5Gpm
oqcaFuJry5ceTOaTV2Rq+9+71o/ZsuXnqgAh6SDUATNgemAhP/OEx1qIJAc/eP1hL7qY/Z9DIheN
/t7V+yt/2e77igYAr51s5qYTuEFiRPVQ9HkvLveaviqslWlCdOMGZWfejBaXMhy2gXFFI6VW6kwT
Moh/vjFzHbN4HG0byomY2bhsRGpMOUI44BQI3GElpycUyAC3I4truenUT2F66wpE0/lkAcVGeoMr
lUAF9nkg7wDvK8TPMWjvlqXmXiqZp6pr81/0J3CZM3Bu6OU82uUCzUlnDeGUt95y9ZDzWq6Amepg
1o18JGrD1+Yoo6t5/24TKfqHY+HEGqFpNWTiE7435YbpP3MUni3x3VM6NZj5WBLC/LB8SKKhgTcK
lwCZ3qaGaeVLak+S++7qJ4zdpDA0YTWlu8Luk25DcPbiXd7j9Cta5gKS08ZEFzCKvfqUrOk0UW+J
srlpM0U2zZxhhpfzVs1aIjMhunr9CytrbgtSiox4zHozd6eyrTKhfyK42nc5hXV0V2ARRIr/2YYw
K/ZopVFQj+xQq0N7YGNYsvIcSxvlTvYv1GFMA34PBvsC3IaqHO/Y4PtM7haPaeWDrPMHlMKrg4gO
JT2TGP78xVwErH7lv0dv7b4ppAnkhbQBjdSuOK4h9GumUoCBBJOheJ8LNvXm/xFbhJ/8zuiSmLAa
5UQ1OJsNfw9YhDReGfnMYU9XA8mhGvEa0LrkhDzQ9YPzNz7rhUOHUnPzzsnAE4ZRm1AIL3smZk5V
/Qk/9Ue0BWY68PuijOrNLAjiHtUHYSB288JySFg54Adf1FNNazwol8cajaZFPc+5CJYlu0WPT/eY
2lzxI0YWPt9gheiA+SE0//+eeh/N/V0cWK/K2/V6qX8XkaWenpU0YOmXL0Caoaq+HQNAyWOSpIQM
WzZEUQKpSHSDwNudt9UTtBeQZQgaMosjvlWc/jwzZ/7lFNu/DgoctERE/rkrluxQj1SxzrpmhR0x
8LNo7qwtfmjraJLObP4b9Tr/uk0ke8sNUf/QBiG9ugsgFP2Y1LALwYsXWmc3NcMgVTLY5Q3JChF5
nNE+AyhSD6n6qcuhO111qi4uvYn2MKPohyAhlK/MMxIiuJNIfXI7lltawHdSO4KAheei7pIQ2KYA
BO0ADsuX5mQMrR3Fw85XcEh2cap3mCy9F+tlUl0IgXoYlC0utBuXRqdx9sxBrxDaNJSVDxnd/JGC
gqovPNrwdWps+3ZvgYv8PhNVPcjSlkCW0pEKsk5X8Oh+EWQj3gaTUOrmmtRDBFEPXCmGqJqvJkY/
69grWL+HFPxyPuWshtz71vOP/J3bJg3bmNSNqTBbwvnbHEAPB171vYY6OPENyb1sZ3HoPRlhw40k
1iD1H01GNhdzrCVxf9D5EU1YwqJ7NOB7wxg2S2z0ebgwyx3U5fIegFidgnOcaqdyFYBEmA6ZQTtN
QAYZLmCXj9qS0C+f7S5X8CrOC9PgjtD4g6LuExDFz5FR/Om0+q6Z8ql2/+XMZLAG6L36JDb8BgEo
cFhMMTywvyQXB/6IH8NBDCzE0XF3y03hPl5JanPMPPPrz/yPuY4Nze3LRMIsZT1VEmqmNyH5cp8u
WoSO//ufY0CsIcBkwPOOwwa+ix1aXnvxAfGKdTSpCFYvGAj2Y8cvBDOJzEZPGAnUfkXJ3yIQiGHx
FZl0YNZ8YIIdIB7KdRvHI08UeLyfg3QFID32F7tIsjooUEoyIUI0a5gnAi39PqUKuavNL8AYVSl5
bax2YL7BcxWGl+Vwi4RGxlReiYGyRP43mjUUxQ1p2UIeLQ4byYS2qQeGsnEAkWfxn2RCM8Kl2vh9
fhRXjSUa1PWLxTRPtzJ7G3ImYMSpklklV2PB9Xy3yISkQGG8h5k4pu59VCcX0DN7w8DTGqSTEdVP
9c6AQq/28etlmGjV5+X5sL60X6DIfSDMX3DnHf5hAOETzdgAhDDaOG1Oapdhwqgd4MN6ipV9hzEv
6y3gaw8GllcBzuNjMlZ+Et774lOP38qdyBqhJuQu1ZP8r4VpEBCin+KQKlpRDrjfLb428MqvtshZ
+ErTZEBexdNukZmo4NwqaZSofL1RdcKaFEInTGLX+zAAk7o26hD+aPeht31k2zbvfHOJHTRU64TP
dq/vZtozJKw02gB5jNqFV9BBQheiUKJQQ7mojUOgdOzTA/VMISp/+XndYEJxOkgfsEZYnTNEIzJy
93y+5+ZYEcTFo9+gXINSYjhktd1DKK6zic4jm9P0jMrDR2DvhLfy1kPvzdBDxjMZMoCswp7OaRu4
Q9f7u+f3jb1BLSm8AU/gtZcf1pPnQBo8B+xO/0cly55DNfRQfeMojMuIETxOfIhxdL7nW0M4Y5fN
vzp6OU3JcXqO1ihYrBgFUTEy6XiZMHt1WFQsyBt7kqw9XrjFpseRP+aH/YpJd0jdNqBrJu0lHSpi
hiHWNYzTv5gZOWXwN4WB3ZvXYmLIR0KrXe82FaBTB09N8GaH2pSN9C+1e3ajTNLkz69y8jJG0FJW
FtODP67ecMxFh+A0OnLEw+57txXBk3xcXFFMNAEdpiUBF4MqTjr9NMx9fNHEdsBqME4l6oshq4da
i1dPdBlOfUDI1UDc1APfqb/CX3q8zDL4PHN6V4hs0ZWaNFK8IGJoXwXZzIQhTwm2Yu34G+FI99ks
6RH5qW5bJKNEVU2pZvp3VLDBoZwcblmcb6yj1AjVdWsKyIYEKagyB6U0hxDGsdEI5VUAnVuHzfBg
07PDaxvu/mKKguvKDDWU/XRFdX1vkxz4PlfnfUtdtRVYGggZmR7OimBARneoCeKKDLJJkPGYdRgK
YK/Ev2YNjgYoEAuL8NBIJUAcfRTVlcBHBdgK9CG+WPxaSwx0nSnT+MUWDU6G6yxq8X+WQiZEK/db
5o/Z8iDAageCFfWYvMLgx33vebtZTvSpFQ2rmOMRtI09kZfqAudz6z/qhzuq/YajwEU45MibFD/g
0jLSO1HaT5bf/TI90V7QhJX++fq4T22xDGjZEz68wyUjeRZF6yEBkz73AY03qFfJtESeAbErQ0fN
Q5qRpe00+OK3Ll2UvtAJF4IvUp+6fjGiK1LLihFrLCvN9KOd5oiBH3ryPJpizoHAFeqMdQ1JY4PE
/0gjZ/R9QhyBmCrf9rVJ0flbRYEIAQOaSw6LoiMjH5Lb7iWYXLYpIXlzFLo2x1l5fyIwRU9wXxo/
QC6+na9HSnGiEONJbgOY6PfuIOxGcltXz82MNFjnWpwSHrUyomaQg9A0AtbGBj7pjQxg8CmtDPt0
ios6sZn185cJFMaKxgurJFpgr1tGxxHDIkzdEWu+AHanTNMZ2jT824e/N4hfvgtWOGkDfVq3eWVS
nNzjFq6JBYiVsx5LtrNZSyEzxqwXN3Ws8ei60CIKNoJf+GedV5NJRxnnlzVITcYhspQywi8QwHqm
1qQDk6XNQ8gOy03+7Kk3qKxIjwSro0U5mbSDI9r/XWqZmIozZJXYKDHOR8mT1Xv6TnqGwhZPwkxn
bUzDMxYCPtSHnlSeOtqMt10rFRle+1MrdKmTwTkq8i7ZmP5M2q0wK9yGZ11dpVpv+zE8z1KWQfoO
iEslD3y5QP/67QLbqkDfUFhCLgNh3u937Izola6EJy+6vBY6txj0bWqJ1o2nf062suji0ZTnVEUp
tsvV4o/S4KjLiFl26nTqy8k2MpO40gKgf95tslysFJX8Z0ddlbSedEY0uRJCFfRDYkd4DLUOFxYl
+kyprY4T+Eyg6HoM6Ib1bxsY80u3xr3JIJ3SCxuvpLnDLUTyPSqEJ/Nc9YOYcSu199GlGJICy7/O
tyR1QcoVbo4s0srKaFBl8kIT/arNII1vH3vIhWlCfsANiPg6jOdSeFfiLip20xnliA3S9MMj3gLd
nG+ZBZ/g2QfPSGysAFteyjkHIOsCsu4z79vS7Grkl6jPbVVW85MMBRXyYOAztmffemg6UDubUrlt
hQIgsvDdqIDhONSi4YvBfxmn14Zjgl8kw+xrOh1kwtwUsiszF0EsGNIjRLjGo23fK5SD1B0etRHG
keL3zz5ct75MSOZ0/eXGsh6VjAFXsrZVcdbpwqvxYJ3x1hyEi+/0Ast1MxJFkh6xv/4Q6jL43syf
KtcA/cqI+HtZ0DTmRlldZ6QKGe3Vd4cnGX5E8O8+f5bSA8ReO77fwX1lDhh83oxCzmpHV2V9It5a
YbsstOOsgCL6NGuc/ub6z7eBvQK8xgoIZLUwtiT7wOp4Mw4KlLt2Y9KnT9xEbHDgxEuSRGdkVWYV
DnDNk3wH6jDWOWiGaWN7YKJdT1uZn7KZL6pRP8Yfa/lcf/uQ5cSu0dWWUabOLB3vM6KZN2AAsZsH
8QZHR2UQMr1W0XnOXHG5nRuhy1/u4Zy7QsizWbJ9w/zRoQzywRkGLl4BGqYSTjMzs18beGIl7Ni3
FrShOl+dV+FAC6UW+ptrPonW2++GsBTP8OMeqX/FJ/ZIH5krFrn8D4NrWNcSPvDCM0ItAHVRNyDR
A2rg82mkH+at5V1NWBp/tEAAiWkGbcSf3zdGWYV4JQIrcxfn/3By+iEkYY7F/W99492suqMJVHpI
Rtdy42TqaUwG3jquxHumFqBrFgPdzYs5MOsUox4ay3W17FF0D2QBrR03mNyYy30tvfKY4tM9vQjm
fySNe7AFsb6A8wX9vTtheM7sdEIKEHroBysruB9OiM38Ss/yJDG0OlSM8q8ykYAqEZ1NN4eMYi1V
BhkHajQzetX7q8+2dluOLZBKwURSv9gVXMSUpcW/kdy8gqikIF7HKSAF/jf+MGSKHHFVt+YwWBy1
WxGzoGHsDUv6/u77MYLqtQOWzYvOz2l0UxvOUJLlTroH6NixT20OW5fSuE5yxOPLmrMwFa6iJxVe
R51Lova4tMq/UTU8SU/IlmpUbHhRYiBXsBG/3KknvPRy/nzT9lxWIzRzOdAct4J3NR4oQ7VztDuF
ncPeYGT3zAyKyT+1Sfhkx7zwDLrhEQ3nw5Cm0cLVrbNR4XYUs+o8MNPoc+ZvphgvM/HILMWbr5p0
jXGarSd8ydk90+Ez8v0/o7Xm0D7+S9k2luyAoy16b6gKel7xUZuPmyk99Ea8uVH4zaYKmit5wMDZ
zQm/Jbxy6OLbOkIhFnQzQlrWY/ObhVp3sB5N86Thz7iAPn0KhtfSb32gJy6iEDVW37fWlgX8tgXD
wwn/zdPtkKcN1Pz6F4Q/GYqyhqQJeo+89NQEB5lcLmPi4fZhJfbHi2Wt/+WsWoD99Qfo0lVGx1UU
7L/rac6uvJyLjiVHc35W37d9zU7J3fMXZgs3Jn4iNRKQmwSZ+A4mSPMgMLUnDbZ5R/Iiv1FVTwM2
NFZ0oeNORfyv0VgxJXj4wkyd+b3KvC4D1QxQwYPUsa3yUU61Mxzu96I4HWTI0pfBZH6WtS8b2utg
diRXIx/WB+9qysvZssr0kc/KZLQiLQuP4wfnFetTtGKa7MiKpvBxwjwJuXimzHKXveuiFf8ijNHX
hCtydUqHeP1JC6ZZ+aGNaJ+Sf2Ud7lkUo+4J7jhtWS7Ei0R4PBwpvYcE3/dqFKEPzl/SR9CsmJ8w
8Ej9ECxDSQ5oX8x10xscN4Ztnjx2ultVBjnyI10RYwok4z77cEtYwG+Tbe6RhRbzwISMjs5umtqM
mF+E0ooA5VFKrvcI9EYubSUmoA9UTLH9W5PPywauhG0pMD9Yu+Q/mPT/2MxLQVMZrhl2m6djCppy
Qn8xjvXN9kNT7BaGUHJy6ublaUz94rgJ0WkvA+RH76m8ZGRBsATg/wHdM3/9P7l5RVeha5hUCStA
tDP27qCe5F/NEInbx9baMUg4jQnRepMjtloQz6GPfSwx9xIauKqxeRpKHG6pgT42OhdoUb3RoX9h
nLHz8KOXJSNP4SY5bTFauaMHRBni9OCEcG5KlDlJelhuyMCpKTVHudPwXGoyFqlkd3CswoLWdrv7
QRIelpvv1L+jIQDcedSNWoJXmBn2kjL7aMX7soCeOMQ/E2O4NsElM1FkFJKal7+so/hpVI11X5Cu
A3UBrB3x9RHKqQaQJNNm8N3z933IvJ6e33Qxp7xAv4H1gNXp1yFGdHkgP62L7/5N4RmWIrIZ4udz
KJYhBZRq1szy/pr9wQYD4nJtoOTJ6hnxKitS3YPJlk5vuUpxJRaS2PojiANxq5gabgg5BWx7f8uX
hiN9Pe3ADUhqNqd/pPBlSV4lRI+gpeQFQjaNniuaQzvi5O2W2S8EBTi5ltLaUKENDlLi3/Q5YhiW
sLnJwWIAZ1Kzp6B0D0JKRa9WfwHO0Fsnf5tI3eBU5097f+TTAGHQcR9Qc6m4igj9SUz7vNwJKG0e
e3pedQjlzob5fY8uY3yz3+kgpFcXkBTlSCaVd58T6ZbL2VygA6iqXZfoo+jc12MaKEbSwDOr7QuL
V4EIcI8wQGS45mjGU890tIzTdjG+n4Myv1n2JR4EKlRx66qpUcHEJN3yTaPmHf/73hUCc+Y/ednK
w1olCC76a5FCX+iH9DJoHrLGXtW2k74KX+UQlfmrif/pLOwSLb3vOI6jX2Mr90qwNUH7aBhweVG1
utK9XKFxLNclFzCuFIPO8Wgt3smZGDkqBx+NfMBFeCuBJ2TF/O+YypZ/IGTBq9R/TP/q55/zZWNb
CkPK6GhhdoKBa9vdY7d1+PJRUayAvnPV0d+wiBjoUKqUSvinr3j0ycM09osHsCRNIltSO0CLL9IR
/vMr6H9NG2KadsSpLFeY90d9u93s0i00Iyz1b7ABQsDBj4Evfzlm+NN1xoijlg8vUM8AlbDwAkqi
SSQ0oA5yftF7AC5lGziBQ5Wp2esekCI2dzAozOfymAyA1CVtwHNzz553OIb25qBDXtMmoQvI0f18
uKt++r98K8+KtU6N+ak1wSznxdBFacNT5YaXRhKuGXvUI/VNwQL8cO3G+1YysSN1pyJPJnKuuIgl
sdUtwrnz5d+i6uCbFdCDLrHvuS6/tEVBvIVwbYYW9EkaEOhHsTwv16bpnHoRrlpdNH5ncD6Ddja3
IRkcEsIZh2v+aYj7N0Pk0ybkpBgwFniqXSRlRUNZmleFwsi0DfWFEJiXoalQVV51JZANG1/hwDz0
RwzOa+3LiNCThyf48LstkbNlpDDQJYp7AS2112nKkB2aWrRYJo4qdDUtay41K/M9dKCXQ+8s4GTi
ls+304MyVwROyyPsreUeAuv7w5AIz+cx4Y9NV1u8ttS7XgOG8KiPF1bjC/3yBrOE/tt1NgEml8Jn
ewGIk5u7+1z74dVIb/scbtKhQ/4oHSLC3f5fjihRmypO0edaMU59oS3knal5GIk1JZOc7dyQOVcT
y5spzyGyjXOWQ7Z1Nbb1irm6Aw3Z6v0vyVyc8BnxR234BgN+asNrThbC/RoIVKmz5ms/OZerGlkd
oiCxJa6a9TO991lqSUZij0uJslHk/98sWfLik+9uQ7JZHrwnli91hhEkTdf6KkoR60uXexMYI3Zw
j7yMw8FXqVy+mqTn46DJ7jOupcc3q+FIu50w8lip7x/x2UhZlznGz4UIXzZr95USdS/f4FIYIjYm
gpAwjRDKkmMWbeZtgK7Z8yNsl69KbdQwXg+rt86aN5v7ZOIzwabQsW9nPw6qrYgL2JM2NV8t9jJI
NXWMGelujC3SWJQYZhwzPPsqIut8+Ex4P30HTKFmLtZl6uJaXXqeP3LyKNeKlrGm3XWYPT7sLiqT
P4/w8T6Ixvkfk3hjWg5wVIDrZTkeUU4IUi4qdrHGp2HIFElUjYyBWdoSTzUAKiXLJI0LPxBxyP2c
NqWkKXIMm/o6caP688PvOEQ6mDiGJiMH9DvoD9Zp2i6Q4cXEQgIrgeoOQAECvPUtmTB8kYqvmGYF
EShR5x3zl48uYbGVALNK1lOExJRhCX/Gpf/NFCt8T8AOpCySkaeXkqC60enlKKG7FTm7U3BxCBzX
i1VVCJgbNBR6nidBaEECAV7t1P4y2syrhXAHk5nQybGa0rJLaNaxllsneH03lqBV/5RAr3y5iE1J
A1vORl0YlzKEA8TkC76o5hRRUCk0snMlql8I64i0nvhVFi7SYV+259Shnx4JOLn51yBp/5dd1wZm
QJ98lYfYoYkvRXHlcXVhd0YQ+6WJdRz1fcqtQJ5cc6N0qLegh6Xdgaa9bzWzJ5bpNfhXPxnuALN6
hvec4/ADDr7OkGGsBUVGOFxWNK9SPpmcJgSi96Bm5ue3P+hRH2pjYg7SRHLBuGJ3ZxsaahQgpD3i
cefGIZkV9+PqOXnLsKlzDabAezoZuSnWOA9Wmj4Hpp7VdQ1Mduuhshgr4tbn3omPzJ/AZz3tJvme
FO+m9eULfS4yQltfiaIKACsG5YzzOzgPhlSL8/rCDsYUFF15Hzv/h2g6aBMTb1s36pKj9NpI68OF
xgSU9tQZMXennUQZrMuFKzqqY93esy1DIqU+DWoo4W+C0yx7sOpUgcMopamHC+2G/8/Z9TCbCE4J
wlLuVm37HAhmLE1J6O90AXNvyh4nUnDNhTxu6P4OtVfDSItoc9YqUGhdtaavu5PaidPmZSwdLjGD
MfIF4keAmA1WvHqBm0qCV/7VtmNw/fh44BOUPsqJDsgIpvCTh5zFarOO5gR+ANW7zx67wIjqSW+H
sWcYyuFJzugVJYvANl2LtzBSVkXeFiP7cjj+XsLFwY8knC0PnvFW8oU8nzGUVMaJWMCy7RtYvq53
eE/OLJYQq62eQbjvUJoWNcQV2KFCXq7c2N6dZhnRavcvtckJc6kgWUoOl2PYPBuQgLfkVdaUI6Xj
iUJJcwE7316XgxRm8Pxr6Xk0X809ZdGfQ1i18x6mkxreLh/YqHaD5L8lCZ4x8cv0c01I7RgGjH5D
sBnYDYkqwb/7ZUr5TuLUUMc0jrBm80Z+s/0Uy0pXzhRcrEtV3J3olSeUrR/vezjmyE5iE/V9+pxp
J9eioBBkDiIgq5pgOE3Jz8E7LCJqwhVMjtO0fbWvsZan6g1XqrCoq8hPqmUBbNWfY2VCpYHxBpRL
A6s9uZeMgL52x7cfYnCb9QV2dJPaogTVaBA05LB/OCX7FXsqJ/njaXZlYzMmYDw5bc2K9bmwIBvQ
79d72WjpGofokEcSbFBvxKWD4vtwM94SScIrFnuZ4XeDAHOYY2jMUejK+Cszy9lpm9VjCtPtZsQ2
67CH9tjurRark7VnztediewbmoqgVAOybm0TA3HLd1Q15kYg5AlB6lLGPkTJKsZjj1M8ybWTXraE
828nv/tkc8Jle47VroYHkAoTtBi282Wj1y26GPSA9TjVgdIcUjvGwR+B1ZFM67zu1z67m6lQA9FQ
Bo3HokIRYgDmKi0NiFmq9E+DSXMen+fXd4p5uKmPwbtuIlbSlRFhG15rQnNMaqyekOk1UZEcjA1P
AUlePe8SuwePssk++2UsO2S1qiPK3kFGQtsiC8/iyG5lJO1BzM2IeDKJP5DC0occY77kD5IYhQ1D
SBlB0DbmqYI7ABztIrh4dTA+uJjJhcEpdrpQcvhDzpmtDhJlA5Nkzz3E0G0tYSUOkRK3jNoRuhkf
rbE2UnriQKY0QbvSqn+hEX/LCY93tRJHINrCASsIdOui17n82DikaT/N5UEe7sWjuM8Igyt5uMSs
2HfI+clci5GWtp1wHHalkPW1RXUSuTk2R8lLR6URAWYZ2xmcX8m5MyZtp9SaVVbcn5MQiVkP0Buj
WpOfWvJfRvrHZU41amxLJns6ZFq9w97SmslSxiBWlUxHm2hr8dpNAQsbb0/CLSI+2UGl/EJQcl+G
Y/8sEwIiJXQjDkgE8R17/QRw4siu4WV4w7XLNwkLZbim7kGcw/VBROtqlNOQ9mQvFRmkbJA0/Zhe
z/7RI9V+73WNWhRdd1JMMk/0WjfUV/nEUIjke8yry37OR/901q0FxNNmzCrZqY4Uj/dmlKBo0u1X
CB2oPdzixWv1GIz+fTeR+IVCZSs4wd/wg3Uc9FdkhCgyjtBBvcgkWgrSLk/olol1U7bo9YJlyflS
lJbM2B4sQegiivnPKHCYZeO0S4TYPpJY+tgL4LwnSnYFJDMIyZJgloimXpo+IM0OZkSs5gzz/BJm
PIigKswkN4meRxDGMnCXLWUOiLFXEVMHUSiTOHB1dMez9ewbKEswlSViMDJMbOZpOACxmMrlDu+n
JxkDnXJ63Ok75HagfzOmIr6h6o5x20v/1zBk0Py4B4WXk1+wsY6GexSUTKc+vgP3LsBJ+OB1GEGg
TKFjyLdVNwaFS4M/s0S5Tm26JVjjtDBjeUjdSatA4lsyfQM8d6lzFAAVA9hDBkQyUiKUEvGI3s6D
I3DOH1WOXFXht7Ag3fqEjdy8QanDMnJPLbIgeaRi+evI/3JcrXFvzetI6xjuJ222gxpsmvhSa64F
1YfMUxW1/6kAym+c0xxN0oZjy/pu29rYohMqxZOkdxjpqpUT+qfSgMZsRPi9aE6k4wu43uUhKX8B
n/ymyQvE1hwKV2K5Tm30ZK3/hTMJIKwNqZzqGZepv3vXwsRLfWOQkbU/FVWxJp/pwLcl4Y6at+O5
wCw1vFRmEuuNAwq16TjnMpjRzfSUkjK7+KPk600GsDh9pN3BN/e9BcqNIB1Xt3oCX/N39PIdT9rt
Fh3y1U+P3tS96tRHr1YION09v5aoVbnzxNMyhpsgdPla3giJv+67plttEEUK5FxE5iUA2cSgzRod
QW6fYsKXVlLqRl5DK3y7s/fGL6abhVNBunRT/5DJdkiXAsWsSPojw0tt6cryn9utLTzjJKYS7vEF
P0bS1/eHIzE1n4ITwRr+K194rTDoql2pAqUmjxA2Lade1s6y2m+eCkF5cX+2i456EE8tZxStCUMC
ES4ZFeE1dgSq9yd441EidEmA9Dvj5rro7Cs/+vlsHAeItdl9UaNL7TM4ymY+2u3ocYQoleBAd6Ty
W1Xoo5ue09Bxzm717dT97XlvnnUf6GukPHSyT8wSQX7U29AMQ9jPd86C7NIVrQ8GdNjPozaxS7Q/
up+qip9rf57flB8neNdTZVsMWGGQZWlERnryyZnRGxSsBX8cu2VDtXdM1aMps7usIs+XA2A/w0TQ
g5DuouSTU4wqMkg1HqUynwPIWPDk5EMpN2pdBdQyWLzOKE+4HIKowclFL2VGmEK5FzXTcFb0zSH+
1KF+tbqGaI6jjPKIb+LUZPGyyPvOq5G+2QfdubzIuPZ3Fuzo+dTBXzJ9j/3PlZVibk9A//odAgIv
XAZGuSDuk9cWLIBYIKxdWtzv/RlAFwt2oLEnrOM+tP+mJ/PR1lu8amtO+aXmCvxSqsbt+gfUwDEW
hnqzaG0GEjgb0VMIYzDB2piEAYhzhJD9SK9NwIygARZvXeLdbOibAE5jcaDWLJ+0VGvtLym/vqae
JljrSBksKZf1Jc2nJHTlO6Y1ZO/mygtQxg79JvI/epFYbwsgIIJ9HLJFy9mxz+4Pw9tDssIHvhVP
GLldY7nQmXIauw9tw583MkugBFpF0LzrQgYMSXEjrCHGEuuMCf/TabpTjWnfgOEEcntdLMYflTuf
UC0mlezAMishr0x4B7rKGq3+96WPA00Gl4vdsd1BSHU1fo1v0mAzisDmWH3orXVi5qh5H6lCQH4+
tZd90o9siWd5wj2hHlJhoRJkC6UqgCTblxyyCbjtH5RLAi35SldGIyuTnvlGrsygwdQFE4ul3IVj
b46fGqBIk5+r0vQskIuMbl9FEEQEscRkklbbGATYB1qKaazJp65Iy3jFaRf5zipeXce7l2qISWij
e5RUuXx+T9QmXZxjCm8cfSuj1ghjeLqZkYldSPX3aTkFC+ajjucHt7JCllvfoAGjpil9P5NzKwHO
/dkslafRE64RtuXF69khkDoZwPv9TKcylH4qVHyubIWWf1wQ6R2QQMM/HKepm6um4S/oodHm1S8q
5x1mN0V9XulJ1Tdaw9rtHGcmx6OrWdn8vOuYZk6GMVIyDzpI3zBuDl5gxsW8ZP/OsDfXEsW4Mfwb
P6e/CDohjXe6GS9CcEOq7hZe5Rj2TuL1Vf6R1EfBUH/WAE13YsuHlAZFgL8/wX+R0QhlrIhJl2MT
5A34qnW2OMYkr81B5OkdcFJ3TZb3zekuheIMEDANIAGOwLrpwwAlH+dDSralXW6s3nf0n1A+xfGY
x8vORwWXQ3DotGzfz5S+ifyqysi1jOkIvRfEqqq6xFV4WlWDNlrf9QjV+kDdYTpe3gOotqmC1voI
5N8mdnO0L2ePTCOfAZWsQ0ggOJroGIM9EqPgghGig4KDeAP9DQqJXppO36cBEnU+aYWq+7cgKSJc
kPzGTnPSgXWENQSAYf8xbdBwMOuU9z68mc4MQuQhCQ2TpPsUc75aNoG4NNaYlQCpJAhXeqRiqpNI
VyQOy14BcqvaL/Jg9fnr68fUQOyFY/7n+hFmEeHfQTHCKpvl8l9q8J8QBe0yqGAPjbQVvv0dvpPF
lXXzQbEzKF2DXTFOnq96kj7qpxlIS9rtla1LH12bPb1RulDJ5dmlL7jCIRRL03EV8D+arrIYSH+K
6u8Yf+kL7ax85eteRCuwS0hwWPpdntiyLDC8Nlgi9aWoCUrXcAI8n7VAfKNUEdecsbx674u2kFgx
mHL9Rvsu+BKiisHjqs4S9lJpOUU35RgIYurbKMeZsyDphWSnK7oJm9qaxLuwUZ9puTJ0qLHVdSwS
BkXPpqtmCZWG5Kp/X0GQzKhFu9B686SBsUM+IqvKtICoN0nTbJF2MIzCd3xdpE1pIPg1aL6VUw0C
/JRBlQ0Lth25N4bBYncUlO1uWioJ8eQsILKjtD2FyvkQNo0owyM6YQPNu7VRWWXpD5CIWPk262e4
OVEHxJpQf1VOjrzL+Hp3yvGl389uX8qMkXXHZUoDg4cBxq9xcp9Dc8gzkVcuHqz21h6gohHZJ5+k
NbqyFiqHBYN+8tYTcmuB2kqQATTw8DOyEAYrnNFSbEFPBkmYUbtdld6mZt98X3/GH7p1j7YedXeF
P+qe+osvPF1yQQIAmLFszoN1TMsBfmygCKkt7ZQMh2FiFnA0PjFBp+a19kmhIPyixPO7icrFww0/
NCfDtM3qT0UAxRdjhjNzK8RcXg1UjJ6OMfLjpQdmcyP/VoboO8rbLJ16jkurqujuQUfkSHuIIULx
I4eobxcBrshAuczobw2O3dPrb97FzgOXbf9/2s/9lFd6fiGCpEZRq6S8VJiBM5GYgKE1l3qwRQT/
ZrNK/Mdf6AS/7YvXNbFA561ChbkhZr5U/rQxdwt3kqCNWeMPx65OV4GiKFdpb68ZAAWrjkyCv81q
jaCl18VGg+fAz0teIItY7fq1RidfxIltpiM/iEwQFqLkbQZoNqFFotVVy5cyYtv/kr3Qgp9F6pmU
mFpDRBbD1JPL/25eL9FkRQJBXSSMYZkjLZ4bqfRX022jFGzh3Gt4KlnwLa+QXdXfD7vaP90jmUPG
VhFAETy3BEmwNIt8obJW8pUw9zPdVPL22T/MJ2jhbQGrj/kKZYjVNuIBaPAvOe05r2K0buXSMbPB
7gjxxcMypOrokhe4viSo2YDTCjqume40xU3sC0uBJccN0gusFFo2lyAw5XtHloZwr179s+3V2WYk
tCaocRrOVJMTI5u6v7TAcsescpjm32cmC/bxtA601TFzm2Y0tpJWBJUQYBt4NFjGDPxFT9dYya6d
54OrOOn2VtRKdQH44OZxcaNFU2NfmhTSlk9CE4z8m8pdGIn1/lbp2cJuIU5uKQF/YQNWN7Jxx/TM
ClkkAo3TsWYHecutnpyYx8TPIrlwMLsVltCPeKpHzo4Gy3JMeCPNeauvL1bcW2z6MjL1HBtqDvGp
AUIGz8qh91XilBd4iY+xLFI+MKUHEqgigmNBA7+YXr1NZGi+4pgURkk7cYLnphSsgNagFKmzSjyT
SzO20lC9aDxFhWgTF/zkA2gT3VV+DAn6+EzPuGRPNgdWeEzP+h9k1gevpZifAdbw9AExaeha7nMw
YkjxDnapGJByBLeZNDcC3ALOufVEc6TLpVG276Aq9BBBuvY8uEoM/wy7KL1ICQz9+MS67/+pNU5O
XMhLQ5SaH+JkWOAsDmQXbSMIIv0kcCaoIqYk4I9JU4FX/+VxQeYvxab1B+itrN0s1OEk90/taxVR
bhDg7JF8WMRr6KiQNCi78U4vSF4GWjdYQ44AvZYS7m9Rymzmi6ZDE6q6k8LzBRbUgi4wLjmYtO/n
9SB4I3YoqwihjcwwnrrqeK+LdJ8EuQgWgxBnhApbeQ8PhlvYOfindJOXvxnJ5iyQLufU9uPYo+PA
VS/VlrundMp3gX0L4SQQRCNu6ltHN5ziSh8IsolCi9HmKIhG6AlL17boJoFpfXMUKH78gjKxIBnY
jRTvXhhJJ5zmpZApzEu91FQx5J6bGG6WhZfBIC+ACxYYyBml2T6tH+Wic0dOJvFhduVlAyfKdgqU
7JXwbCQwnIEFUtyR523a4isJDiNXkXyuVyXaxJ6ndyI0XOJS/r5nLni2B4sLM9Cjoh/XQv0k4Bd6
v3NEE7tMia+Sgrp4I99VhY8qVFR3+IsoukuznsNLmCHA6b5diNMW/akwQtatw7eesMADVOA8wgMS
z+VMel80mJLoFxKaDKmzxmxrYFO11n3FseJQ0cXnuT4J4VG+3wEhsxnqmT6IobvDel7cNneraEpB
4wpJADTf7mL//8+/E6m1Pigsa6JnfkJKQILRqY/dMqKYqyODvOAaLtDwYNb2ODWtVl+wSWQrnJY1
2rT9IB4mI6JN4futBXz8HWXHTFVqzgyv8y1Yj2dYvlto0DKKo7RjAlP1q7dnpHpA5BfcxWu2P3me
m8bve5V7yf0ayA1jDfu1jpwriBqZkCUdWBSA5vptNO9HpQUzKmh/sadDnW1G88NaUinZO7eXnjY0
2jz4dXRhzh0CksDCyf/wSqXQD2lkfI55wTslt0GJvSAR37pBVthZ9AAwwZBRAnNMngHWsmtiL9Ab
1i0Tvoc6hw+OP4/Ue83PtEJT60V6rK5ZodqYRrAV3OHayceprA+Tfr+3vDCroXKxqTSc0iK1JZmN
+69kS7AX87A/QEOo6HvvUmWE8K/r9tUrU7qlq6/TaKOgWoAzTzDJCEuQmE/SaZVUDwew5Np7ofsN
lt5wRMCo1IsKvzPBywoDOUhyCvEkX0AH3VYNbS78Bn7JsZk94yVDh33xswOIDwzpbQLpKwMDX2sb
WF48FHZrVPUAPzOZJNXCBW39JZlCPV25HbMzzJ8mtLiLroD4T7oAygjBH7gc7PJOWCXfxjUH4n5y
CbTdPNnJcL7lWHLd22+H9FJ5WiaWlJt7ahR+JrFgOm5RvvxWvMxk6efY6kZ2gOYFlr7wFdXZtZVK
Y6uV7DS/IxATcw10JSzaW02GrZ3YvW7Ff1PIUFS4DWclheheAYgazguwylxgWmUbaLw8+7FVnIZb
q3y/RydyAb0DC5GjRYTFhdKdsdO5rBbitfW9iVHMV5OvuEI2VQzacIsKQ1UNTvBYGglsuQeJ4wcH
oOl/FT48CX0DAi1KBEv0YBZXgrUPmuc9/7mHqannkBAWJSOVpzuD1h1EbRC/VpCKCaxTM8r/KCO1
XTTbSOXjomwLjJiQol2rArMaBsDeKrjVU/PGI6WmJXkHlpXSDyJef3YRUlwDgFPEI9z9eo4FQuyr
5u3g1VqbvPnKVsR5mGcUSKd2hNHoMfBWZ4PpS1FqfMq5AUfLFF0cLNfpRh23Bzi9iyvinamdBHql
QnKlJ+7cfrijNGozlBFrhVME08uvmeA6vIEK7YoqpbGsK/mfzB6LR+LcJ2mmAKBiT4aUxrR9pPZo
qPlrHK1PkBd5IuOIEI7JFyKVjOG87in/yNxDt/oa/5kkftqqDOlmkpdz8VcUFVEl8uT1aTWaq1EF
XPL6kWrYJYBah1EuUMpXMujqAdIcTYdxGC/tKo09KEa011CfRWnYR8AR2omGL3L2oITNG7xOi0e/
zngbsju8jY1BhIbzAvRLJNpf1tCGr2eJMBlp0e1azakdMaHOypyNZhW0zEmlXOZ2fQWHIv0qyAyh
1AeIqAKyafJmJsGJG2u+RwB4/UQJ/w+qp0SCnZf8B6zccumfsOMYJg5bFXnoydfHhe3U25QjaF89
jACBtmAFlp73Xkx7wXbsY1D5e9VJBWJ+tadcoAQYzzeSCUCY7RkadSkh0dVsxwha9kjctEX1n5t5
fWhXCfAHy8P/tHJ7CJv5o/KuSqiG5yvGp4O1FXxu5/E+YoYKuWz/XC3igVBKZoi4+h7bdx6ZZGRf
lXAuE8xPuQcQNxYLjUgrgP2iZqnwymEv5I5eReW9YBJHEzyCeCPqU50E2iHmsUV8zolWD+ZEbKK2
ydUZZOymGoTuDBLS8xrtm7NnhKyCbrp67fj8lAJXfh8zvSiPwd06VKH06yi3ld+h9Pj9MP288//i
leKNaQ0gVpDfvZgvNXkj26kljHYPgxF5xjnHJkgZHP7raG4LmcptUjOCwGol0O1kMlQwVHspZMRM
ns96dXViV9+KM1hEMGEHxLHlEwI79I20iE9PBOzvu3hnkOEsqlxhm0PXoTjQ6CLl651rUN/sXNRY
7pXNz33jQhZZrAMruKRjKbZF9ikcBxeW67YIyGiIRjv8R5FErtCHCcQ/LLckocfkSPr5Rs6hVXR5
FJUMzlKkSJQeZc8dED7c5MKP60Dks8eI40/jgtqikUNMINpRmV8PCIHwROsGzkTi5MiRXM3wnP3G
rIYiKW5XTX9B+58r+vXaMMcUc22kedYpL/enlcFLFnpm4EETxWTnepNKZeW35JJXbbBlbdmfO086
y2YUguNvequV58Z2naJSUWvePXWUzrflF/Ug6p8ZDiphJQ2qaA3z8CpUFWmCfdkDEmfXyxmWyIyW
AWBJelH+pBuE9qgHuaOXpjFIByvQlcSQCbmx4UekT65BJ5XCcrl6WW7qitzrRJAfLtewyImbwWOX
GBwQmyC43Kpa5+OoFO+qtodSl8em3QaiYqKQYITqLMDDZqo7Z28o8XfSCHIM1rWNp/rR8cKmubmH
4H1oonBwBgww9KsPJ3mrPaWP6Cn3arO/gh6QpkxIXaZK1fB8I6CYS4tNCNB27enTU8ZuswsrXDeO
yYaK9DwPQAn6qfg81/pXoxIQxnCW1z1ztCZrMgbluttw3ODXlEuMvIkJM2Kplzh30+DTxMWtS3kZ
aY6fSG852/5NG9yXAVnRhRfuumX4UaNnzMnSxcfQv1jD2v3nOyan2V+WpoZmf6at8AaUiLWqS2Hy
y4si7TjecZ3evs8FPp4mW5HC/+9ydO/gHU7K0btTMuGQOEg2fpWl58k11mlVif91nqC1oWzd0jQZ
O+cc7WG61XdXyLiGz+rgV0W6v2qARVCWYHBhRnkRyF2yhAh6exscMxS2bV0AChWVdzzMVrpYdHxv
7PPTG2GyGwRjGIUwUO30nmPr/3tGzMDq5Z3TjTvlXu5JZc3CeBfnsM0f92JHrItjB5vu9nlyHYka
m4iVwZK9H4KqMNEOLoByIvhoN/ghJpWfi/hlgLjhadER1vK1P+gBaAsgcbIXjjn/TXgExuxrm1M9
atf+CtJazU6kWV8WsfO7r/nhDl/OXMRX8bAa93j9ACmrwya+kBGtA0CWfLsub8EjAol8DKjQSlQl
cIylsUht3JDtd4uW/42Oq1zB1A8Dil5cNj+2M81IALLKSShMdwMt6EhWtJOAB9pFjfeQI3g4Jy2p
h72ccwvkf5jvj6LHSpny7Ym/CtXY7TasrXTRFkEjNPwYJE+6vVUZb2YMcwtFsp7ePafyV1PwWGNE
GOVtOGOXjzvEx9DbpeXbXydCq2zeAcoHf9twKViPgbmrh8QRzkpWfQwGbxxp/4peRQrXBQXISbXy
rzzMAK5+CVxBvvQ3jcyWeXrf9KDNLJDXATLNBvmvVkj2NnkSnPgo8QfiVZRypM04YYdYt9mZSm4i
UUtTCGV+yW5sgi+qXPcIwoYplkynuWhJzIR1e59NWmNwzJUefren3jIFtOL5F6WnlJ/WFjCAfasp
emDWcIJtKwjiGWsWXTBtpaZwPOVdXdzT0FHZU7zyL+LVfApXT1+SHrD9jUwsYkmsThuaW5u3rCsI
ylZouMXlaK/FR/eaiJpsh96IB6z9bM6zE+DMI1EgEWz6qGNFwfLWs7E93On28OduQ50ZdJFWDRY8
FXJioBbXh1Fm/ymMM6gnGFC1Op/gsDUCSLAiLzBMPhImaNIkBUygyNhgV5EKhle3SHC3HSFtMGpf
FO1Mk9eIvGaasO8goxwixkhmVlVl5wXY2tfFd6ZI9oIi//TNRmGxiG/SesQrziNDcjYvrnntSNL/
QUBk0jXdIkx38bvzlIrTNKuujJOVwzNXebkzxkSF50/lJwsX3YSw190mXTIRNvLjPV7+Os4bmxB/
ChqcqlFeiZAv7hWf3sgPk2W9W4TeKzmM6NwP8E06L5ky9W+18P+K4X35N8PpsIxn20MeTPga8LJf
zk4WVe3VP2fDKOZc9dLUyRxoEabYF2azW3OThAxjob76T4mTNNc2mSpbsamM6kqwH1taSMbB+Ki4
gJu0kbA02O1d6KQuDTYiBXYnEKWrkdbwotT2lSzQ+HK/hrmDdXqN6nzrTITUTZwNl39vXcbuU2cG
tGfxSj9k4eABKfT4u/q0suZUhEqdRyRNSpAX8f9NUUblerAtr3gS73I00s+3OWDmEV5EhYgo6yvF
GLa/5rpRoUKQjo1m5HzEioia1ar6SeZyeNPYEKgqK5Ap+wiQSaiif+IKvteiM7ZLc5vPAPCsYOnM
waTbI+/Ahco8eZiM6dL0qrZSKp6eW1fh4fpTTlW1aXwcQ6bDnjwXNE3LkWuwNmvu2CzAzVWJ+dw2
Be2spyCS4OANbhQ4uWkCbC+UZdXsklHT+POLOMSecK2K6M41fYYHFX2hTbGUsUwJHJYBALNR3k0g
iAsF1QvYRHht3C0W4ZZiz3poNJofW0JT+1DH3tOfjvFhq8ECjuOT9TEYOacTeRp4QgMqI68uuyDE
FET1ouXf7i2BLRFE4NeLmIAyCnDR/y17NIQXRPwF5fRx5Rh6rv48se6LMg3lM+3WnxVap4nBckz6
MtCuYH/1wdgBexz/yl/f8kE4BoKLPgrVfDVQvrOPRxvQLiEGC8pH+8jS8FSATW4jLYYAT36ivuTK
gw5yucH3d33Yu2cDtQ16YAmZ+crkwQ/4kW7f3xdDfkzlY5lKaZNVbyCRDMphWB3vwwexZ5SiA1OV
pGdgVb81wPZkxZZ8eXTUS2ijDMvOaT3abRwu8k38fstiGpPxCYtkq26zWvcJ6ECldIb6UCc217Ua
4C2tejtcwT58a4d45VehFkQupyt3UxKPK/YZJdQJM502zK+FR0aFX3UbLIb90kAPMhVuu7Ubd1+e
G/fgeFJOJOfOfDUHtZJK9wiKbKhpmxcUMbOUqjbXDwqTg78UGtYzLBGPCKqVtBO2hE0vcGinh0Ei
++mJJm/A5cpStjPGrsjmC9zNzi77OHXGSJe3zVyNFi230mzNSOLqzAg1h5wWmpb5hSRvgdvuVdGG
N6LOG42hW7D9Fik8lbeFwr2vYObjLgYoxP2eW1FYnP9k+gLKHEwHyPj5OZyaotksqwKwrNYKK5aO
fdQ2Xm0X6rMTKCcOSdo1LwDNpvxNapMn6+S+Wu8D8ONaGoU3tFSOB786fD8/JyUGQ/NmSwkdsa99
b7SHInhXTHxsOUDs0IYDOK8QZkBzzLyzw9W+CcCwT5iJMfDeNUsD1mW89Sgd3M/93XiuvnMi/PnS
zJ3zltb/HjLfk0FcJ8A7lBECNW2WDLbpI8UEWdgC9rzytyOLaxqMfsi/S80RieAPqCBA0XXiVZ0q
1xq7hmOsMHmjkrkWQAemCpIKYgLmVchYxs3SnGW8g6kIHtLIQ9rhQxAmA32s6aUVilmzrMsx0Gy+
MiGs1xYV9OymhIydtY07ggs47JF2Aq8cJAtsoOXfHJheuiZLE8FN/de/VHAQbitAHoZ56Up4c3qj
FUZHTuCbI3QLmDD00mpY6wdBlTlcszZIMyn7pa0FBf6Vlr8KaYbf4dJtev5lbySf43gd6NKHhICA
TKovXQQVAfnSkhzST7TT8j0HteQuL6zljmKI6EQQnqfqzQ52RyHWfS9HRXsRm7cMN1stNe63uhcA
v0Nip+sabgXmG8Jbx0hvKkbodq25ZJnwgfFopdfgamudwIrqFJdjPU6pMcf5vYv9tuitmaziHTlJ
YW079rPIqa89ZODi1/pLplbtsbwccCAUoJgAlflmxi4O6HdLVlouSOWDFUTItyFMIHPpy/yTFvBL
iUWu2X0WAQ05AC+0kxhKwoMqckr3rJhSgx1VT5EE/eLYN5puhlcJbfLlLiJYsV50LSlI4sKg2ZFR
lyYqxxi9Dd0CcQvPDimk4mWbDBGyMtTYp1R0KEkGQ0KoIov7Fq1r0ow4enN+hsgzzhW7m1M+QsDo
9BLc+xyFWhq6fPrVv+AYMpGbI81QzJHQAL8SRWR+zoNYqGdXpgaElWe8dxnMnDI50pS5jaQgvUHH
5dqRAU9jQuVNSOWBzwBij5d7sJaxqSrRUI+v3+GfyFR6hRm1+I3fY5fcU6DBv4c7kvpQoK9lq9CU
Jhgd1tq5kT5qWOvdxhCSqnTEarhgAtnpBrCm2gn6EXGCpm+KGDQ5bZHYPigXwPB7nvakX49K9dqW
I01S1sTv3S2rw3x1WhqIW74VmD1s4JnM5ce3Sto9EKWlc18ycyivfya5PbFhkVhhIbgTO0E/raNr
SOPKbPgof9iksWLJGogcxgTYaMJR1e2GmM5riEgkrv6eVogv5/h2JyA6y4BSz3VsHzwDxvH6x6x+
o1JtqsnAx8cZHpRQqCOx0IhL8kC2cwBBP/JAK93S4OvH5GBao0KBqV7eTyST9qeSeK33V2DGTC25
elcGW36QbInzmee4GPID03SCAZ+u3432DmVqtu9xmoiF29/4Tl8nxUPGzrJ/EFO2MsUxbAzQ+hsC
oqQqCVFXsnsobu/5WqRDAHcXndpPyzp/knS01xdUAjD5Uy5fTSO3R4VZYlFvkuDzG5gfwQcGrCCF
C2jR7SQixFShEJhkrLsWGsKiIuevqXxgSa3cduopbLRmVAGE3tv6USfzLgeNTzd8HzCcqEuezV+4
Gk12ZWbomjEXDwnhwH/JI/MMDNuWubdG96aSLQ+XqYOIw/yYoRvxl9ebrAIXc23p7AFGRmBpldO4
QLaXhyajGpUJ0BOM7/5XuLBHhXbr5FOviE4WnOutA6dGJTniFNChjYZfs1xizzsNJCqeAdGwQO22
SLAPLa4Jqad5oJgRwAs9huFc1Q77cXG8BmOsA2i9rcKmTfKO8pbPuppeJWYPwlRRG3gE1A4wtLXL
0WhVaFY94dtY2msLL8D8qLl41sz0+uuA+2innE/yJnPWIxMpFgkp5CrhHWt/uGYgRrpk9NNPR+Rz
y31iVKctYmMwkFY+fJ7fUDGsnrdOTmURN/LtnT4WVO5Xwm499Fy2FdelO8im9GXvtD7cdgEaF3PF
oLeL2pK9a6sg/oyRgYsS5zGVAMDpQ+/VhrPnngWzA9UQcthSf1tNCI+uDiM3nwO3qBX8umFJsKNl
X+/asyn0OA1ZvgY92rGisOGA3gXOp6MlhiOkDcWPF2o7W+iM6U4QlV4IcGhhu1FkPYtkRJA0K5tG
0fiauAFdJH1eMlRU23nfCOf8gxQ5FNX/biTL88Ry8I0sv08Qm3YHlPaAeP8tkTWj1XtCbp1aFts9
55dAYMYKTIrz4bd5or15exoukpAsNK0j9lIWE/JY6QT0ZfB3YSCnTEyYuKR0SXD4ENCkfOrK3O9/
jDUuh8lUyd2HeXxrAl0jFzLdyEN94t5/JX7LPVQMjDpmXbuRnSqhIDmUw7AOIa/jDMmpx2nQOcLJ
tFlnWPkeA7pMV6mbW45t1fJHDnEzWGBzOMeQWUn16Wqhc7m2BxDkHfJT06vexZLdajZC2dVnEWH3
zGc74nYgTGTLvC5Y2IBigkZqWwSPNj6kwdWtgw6BwVmuEl37WdLqYwwCYG09MHLytBnQfiAnm/su
XqldHJb4nyYN9u3ua3VJExYZhoXD/AelmIf9PROtjKHKivO9/pmNLgI3b/35Q+ZZn2CulJSk3ANm
QXm+btM1m70FtlCgZvhRcg/790pdr3qoTRUPzXRJG/VqipTu6xyRPCn6rZjohnNh/yMB/Ye/EX7K
mjkJ/6wbq5hMcIbiqeOd1vFt05a+tbv/Jdup9MljLkhobJ7xD05mwFujyNPEzw2eAihoFoH4HhNk
AU00O7CVVLmZlisKN3FEfxV8CaEPU2+pC5KQWFHgYj35tWr56E+3qzigcJG86hhRa/FWig5wLT7r
8519Sn+jFzMf6inKrNk7Kl/oDmNTKobTtrC7/GSO6x9US8ESoiPjaFxL+4xCe/xxa5VVYOBfakNQ
sPQ24f1NMf7K129NJiji3C20D+qfJL4nzAIV0eUZwX3BcHEA0Yenn6U4bgHsiEEG7ZQ0ogM/9Qby
9ocGKtjDT4BpUyZP/5EJpe0sVwyDxKwjqhy4Ui0+8F+lii81jk2KJc9gqckqQ7RiOpgP9H0/2vnI
qJRasPxkVmdvksNvjZGjxhjnmsuSQOo60d5BNXncyAcWJoWksjDJ3AFg2wiF2WFdYtWwKTX+kC4m
eXprS+vyOiMMpevtI8MbNFtR61n4xJCmCHHvHmAceVGCpkUMpnlgMjT4+7brmcxFc1wdWQJRHpyp
N0SSlxvpYaz+blFTVM/GU3ZVCUbFrlg8P5w08Wb64FsMfRbyZzkCrxcoz2wOijTNjEV7yM6vx7JK
t1nNn+A5gjpjF11oLRrtDRXL+B/6AygdmI52MHkBTJWGFCSNeKTEMyGCZKgGO3MVmLWdNAlIaE98
bLn6VCGDrhzA4naU/gNzx7bZDzt+VDSuEeUna+YKHqWAHSGicp7L6B7UFOtguBMGJbgIvP7pV5zU
l3xbxB3FQZIt5fyhjgprGXKdiaSih0arFA/7htZ/3WOOUAA8JU+maiC5WW5Bm5Zi34OenRDMOFps
DgoSq//9hT9xl1JFFMMlsDWx14gXVLDk56jAEa67/TQRwmioq52p+BEX7TbwhxBLoMwCEs2zqRvA
Ezjzc7Dm66t6O8Aq04ASMFJWKcCfI1AcRoQ32Q8Gl+hvV43uKUDkKHdK2+ePXwskTyEBQB29SHiM
kFil8oMvPvq5BRIOnnvGzRemvyuCXU8sHaIlO/dkN1g30M2oWZHyxB/0tYJ0AGDz9eKD7kufZh/G
p3Ku0BnWv2Ph2bzkMIMRYcqAvhDzdBfbN2hmIKJv0hamfyH32sTcj/DMq3+rBRoMZzw0nS07NIPT
2JiqvHn5aI4WFSVWZ7NzF0Rt0TY7azsxzHZqCGphVdlFJ3ssklOm34g2ETJImnHnKd+JT7kreSsc
CqvbxwCDVOUVqCaZPrk/400C6Jdm9US1KZmNXhZUhzAeWEL1VEaWhvmFdwjiTo5/VA+TShvYVpLP
CFSPRENijc4VnnxaDIENW1/5VVXBZ/ZJp+ZB6xFHzpZWOTDhjHX2wcCaVZzQ3cknmSIMpRTFD5b8
XcMDcJKHNtHCHbs4R6G4cVOdh8or8meT5hbwDbqmpbF6Cqe0l3+gyQQZWYjN3Z6Zu+WorGqTLTPs
5XBtGjDwwlvA1bhUCqdPuiLLKWgBdoUppNBPTSBylHF2yvtRDHPPqmN1HZE2vGCsSmcvbvqFGAGv
xDuW4JfFU1stLem6MJt/VN98PjrrzcKD9ceiTD6qGRy+zp3lsHgdAqHW+2mg6mOeOgBa2ENnyI8B
g7Vahj5yplIboy5+dCeR/Yf/Ww+o0ZZ549wp/MPafiRZUy13g3VrMhIVaGFUSyHbHVk6oEEuUzF9
ORaR33LscCZecoXetDBWxxlXz35Fwp3uYrNoMadwczI5yG7nm12gQAtP01J3X+XgInangWAJ3Net
LGl5a5j+A08i50jvD0F+j98dwV82AmEVV1HER/ZHN0q/RdQGVppoaLAAO0TaT7icc8pyn0hSs6nf
9dUhPnOwsGABQyxLm3YmS5YX9DyX8QCtAaax06O6dUGrv8C8kCKaTarVEQfmLy3biYZO0JGi9i59
2NrhnRME7K1I0ioVJrY8hD4a5QVKTnpY1ogoyarV26FqoBMzqG4/TTMSfDuBaqxGVMTBQ7TYQLGi
ek25NfiW7D7qLTblBnHuXdfNv56L6HPPwxp3LTtWjDzwf2QNcgS5Rd4M13BCAHQIggGYTexA/5g4
pd5u2LPNGRFOECN2Yf30sEBm1GDL99RpQY8CNefR6NmJs7IcQ8qnORoRLAA0tBks9ylnP2JwZ7N0
K+elj4WKdugkttI/vnmsR2eAo3+uTYOehPw4FA3uyb7eNvcFFgTosn1C+fe4TuXYaKwOoJPArVTs
I8NBkR7v8Liz8GxxGuyj15/aDq/VDc7C00ekTg0W61fy7uzLvTYmuaK4xR4yvsKeNvoPWKuYtKNV
aRWL8uYYabhn7k9t3fEl3JDUytukGcSKcOsX3BApehfb2WbNVJpmTj/zx6rH8xigGljV0takavvr
yN1T0oFwhEU1QgIMlzKevKdOCLYmNTKb4hHZrp0IQitzK3/Ld5ap2w/FNIk+LhMcHUDvoL+xfvb4
hcnD+jpUD35FDnw61KdhnidzGVylRtYukB+tWe0exuibV90e4TOR/mlHIfq46ZQo1JHuQYMDb1jb
GwaEo6nuS3PbFML4ZTUInFzg2qaBSg1batMza65+JyTWyW8hSjjx095oD9FqZRrq9u7ic0Z9b2Le
Qy1ClsX+6QPW+j8HVnGoyMpT2c3vDWILW4Pwp1FHLH3muD8xP7XF81oBX+jlDYekdw+yRLHq8kAq
r6hdnSReZQIAmajyGpaCeGTad+5IirvRgoHmcm10z83kl5o8q+39Aihks/KDwZpH7oQQk+exPM3W
d5bxHHnQGIjpZKnKXL1+dcOAoxM5OIzo5fZ2XOvJuGfjct4Y6kyFJ0bLyCQkClHxFKnYvZ+VfAbd
qZrEgCwmhbuzwBY7MWiLKGFvmgmfYWIf2DR+dp9ZBP6az138czXdkPxinowA1u10TQwVse+KoZyD
Fe4kZNaprm4ySNhtUN5G4Ujwgs4Kxc6oixFwncKx2p7GmosaXhXrjvl0CrwJtXZ7yOHQaECGrJYj
egCbccFX9lTtQFf3bETE55ZG0Kmu7p9T7vhh7Azshyh9s2AoQo/YcAh2LpIjHOYemgaeTVLbzT/D
hW3H9TV1v6GogvqE9Lf3cttD0VpCqXK+JTSEwaxqnpeFWngsD3x74bCoUBRwGDVxsSheqvSg3UKa
v6Zh2wJg7XxaAgh6XuO0cUUD6qwv7qITYqYMhqvYhnNFQSGGH2IL6/Tc+vBOj8MvGqwPl0YBAUZD
JwIUvDAn6vE0u5jBqNcj+wdYX4ZZyi5CufHeiibs8qWgvEpFBpvzJwarG4kXrSP+lj1f3udOCRXr
vJ35rtjWqJdL82IrChs7trxjH3+DHvqzInCMPz9PXq/heFd/PzRJQFZvsGKIWW2zI+3x//ez4acd
goH/DKYjTxeAAW4+hAI6x5JTEtScQFQai32BHjps+rht1YQBnEVGiAdlBEe3ryRQqJrnZxJsDVnF
ypf9vwXAD5XhLbE7EN2x5w8jEXL+BHQ5AV4Ijz6ziPcgXCqxAZrjwYH6vpM1bTjVUkE1OkDxtPO1
KQ7iWVbWZYrTiOkbIEuzJ6SCMUlhJg2nFC9sTC57hUQAefBsELYEFtvzSpxaLYVfHmg4SClA5Vhd
NRsWnlHCVl6kLhRXLDSOyxrYLOU1zDFd/rvtv30AVVsI3/lIfeBZpgxTddAcI/hDCTuI9rtOt2LN
5Q7/TptbpErnkzbKspDG68DjWoWVnZuHjsXZUt1sRtfdTVl22FFZIXr28FXLPrYBmjxcEmqFWevf
wgUVFKTDF+yIjhWDmpbZibA7iswvwTCx7Tfd8lRCyO6+YcoPeI4wmRhe2wwRaeufXyqi6VSvUE8E
9iLDQx0dMYzIazOMbmjNvyWZrarPz5qUUbagUMPEAFXxsZcti7xZU5/qqB/v+DgYPOUBnsvrluUj
bFDj+xZgfGVEQxwGZ1EDhf5wQgvuJQ1qvaHh0HPrfCEfB/cgrXPLt2RrTAdfc1UO+AT8Lif6+LLq
7Ye2Qrbxrh6ho++T0YU6XkekW+r7ho1YxdmpC497BL7PYxAT76AZs2RaijpgE8RxQXzkAVCxOkOe
RWrUcI43FPXW+v15z3wjQ7cjiKz+ic9HAkD+M0sj7KECaNDhZDoX9q6fzM9FkDHU3UKOKUAc4qqP
lxC8B/zRzaHJincXbXlhLi9E1V5FD1owPzbst/PlVIjOdgK7Dsvmt8RFpZQib6OqGm/iqTokYC6t
UladnK+WmaqHgCuAt7BeGb3TWmawREemNfxGVuKwO4o2Al+cQS6obhDg8yLazZdwGDOLw1PJVHZY
/SZWxdTAPDywSuohQSsp/MBCSfAc/TcznwM6KhRASmxVIWIecd3IrMOtKAOeNqlb66RRMXCWFD3v
knhDOTujcTTIoCsCfkdd0baGqH5scwgplWcEdALLWn6yeYvFmlJ23bf0WRATJsskIs236LJs+UPt
EaBcBptBzuPeupIxEwnXZM5sOGBQbmghoZvjihKuYcFlMy/15bFpRXHg8QHpgMeBxFtaOcexFrMl
3BLLVFREt4CYlocRU5u7PNemfotaSG5kY7UlndBGHnsBq2K06wms1QwMZVLJjRQDOMZkymK3rIe1
ZKRxPy3+kabtreJVMsSw70+IcjNjDqtiKzH2wTr6crKvwgSiYzbAxOBF0qASBOF+VBDCgXzRPFzV
08GKDBrEmREuoffrUPQrBDflwvkoeDLnaKg/uy1FvJLytiPa9jcapDgNU+8qEB9CThuP2yOZrB7k
zJTZFbQUhj9akqNK1YdQzn53w1A11fh4NqXMxgTSUYbGVXmWprO0VOuHArN71wNwmGJTLQQreEV6
OL3sXe8thXoacPzdwYenaUdzRTw+8G5d6zRxOqe0h2u9w82Rto7ohHyy3cb5pmdJLcQPre5RlJed
MPL1Nk5t1DZtnMqbET2Y0dwbi2cjTDgpBgp4RpnQTbXXWl4X4ECWR8qqhw5N9NmCyb/UCbUvaA7G
WrOz5N8LOhWehMU0i4fXiVc9JDc8lfE351HIwy+iOe1Kue4/mo6iphnhsMt5YPSYsBuMJ4atKMIc
Wi6hsjIEjyvwXkkNouK0aESSIVBotZxmzuudeAE7muI9V0tqi5Q4mLeJnlxnU/bMgCNCUM/c8UL9
1/1tsnyEf7S7h0aVgvDIzT3HrOw79Xt4wM3lA2fdVvO6zOoDWzu9K4VONHu1SImnCGSnAf1ORmTq
78RdBhjzr2++3VZbd6DdSZoVzEZ4BZruTVyLypn49E/m28zN7yHmwwRoI5t+Ef0b0DGYc6/nA4Lk
u3kSgzcoVW+9FPTUQMB3Hl0WTjahMcYOUNxNLr90QVbfNPBkVSi2GlzkkvvwMn+UNC54xhj3bzE1
opkcMOkR/NX5nsObVZc8nFMHwZqvWVZeh2sPTwhae5sxixO6XovoGOXCEYD8erDLjEj5G/FbCX9k
R9PmO13ua3YRKq8qjSe5l+Wf6N2JdeStippVa0+HTMmfQwjuUOCIXfuLK9atsQECUCM3gMpY9Zwg
Z6sUOrUUufELojg+iBSv3q2CEGptgJ3H+vfb2kkyqSPNW3hzXqqy9NN0VAjTtK06rPZLbwRYXtMo
RmAG8iVsMEV0R9Njbq+2FESGoRIC8K9smVreIj3fFp3g4x5Yu7BCp3FDMfrkql+t+EqMlUDLmdeB
dMFrVnlSzbhth1/HA8sAPe+MgpoISn+RH30H+jToF7ViAjG+M9u81amFs8Sbt+Bk7JM2kgf+fjBb
rHwQlsPfVlHHOWyxq2d8D41NYeMTly/h5voqorCrx3cCmGlsDD7FOzfFuLdEXc0TCrCs4itUINzY
vkHvVqdN6FDGZMGeMCvOPYEmtXGn7po2+kOuIudKDD0RPvtiNhoAq2emq2RobilL4miFn7jcFHMm
aqtskJczXLOxz+eKPXr1XBV4yJw647L3N47t1L3kqoyCK3r4q3L8C/uRkllVIn0ar6m6VIAD9mAB
wj+YN1YohDK/cYJc1G18LcN37G/qjTk8TVlSu49B+xRYbVV/C4KJYOGPDJb8CMYODtFJ2nh5Ukky
kRRvYwPNv8tWEw9V93ahDfET0KGO37g0vTRV3qKnfL+9uJcNm+H/nILrwTRiUVSqMBz2Oct/8f3g
JdbjimlPrMD16WMQXD5O/sfBMCSKsb6bjFJRftv/FgHSyTExDBatzHj7qE4hkwsp4grTOj8aRNMQ
BxQzbVx04g9otvV7BruNtOhtEE9AYWUdW5nnc3Dgj+KDOPWTgamx5zT7/35l7r+KHwBvw3FPruRY
3aZ55bAxj0bDz+XOyd1JXairBnxbLJMYALLqvhdWX14f2EJN4jlSFsXiVXiEhxQRDh4BbP0nk0+9
oVJtWC6gXcwzWBdsmFtmfVaE+xf3uHfrHk8MjymtkRT3i3AUhHhf8Qj4g2W1iA+hk4rskzfZRkeC
ndhLucpoWWoz/bGfo83HYxydcgRIglwooIpKsdJN1WZUNR27tJ6kDkov2C/0lr0NTg37p9MT8Uzb
X8siwCvZEQ2rATmcBLjTqlM6JVbyvmAcTbw+OLRTv0yu86aVbcwDatPZjBV8gR9Vvdha1oEZITFw
H2b5/AALMRL96NAsADgU5Jh5yvw+Jd3N88Z7/Nbu0rHR43c5wPCo7Jh1E04IIaJXKttUSjCIr7M+
EAUlB6jtp8GM0IpGZGmQdiHKnTi8fkki/CFOxqKp/lGTyjW8dUWuMTEz4/ZZLoPl9YSY8Kb3aZcE
5TfoV6UV3mJVl2y9TJvuejXOw81/JxjKqhoJg3RmXeVli+yBL0239fq+w2pqTb/Ttb/5dh5AmXhg
oklFaEBhaviE33+MubIArrp5z2EatZ8r/Do1mRIxUKOYBKGSKIUre+hEvOl4QLFPbjmQw1mvVc1K
Bh/lpsOyiIISOJl4hMI6wal8Qw3x3ySUNrfJQu0/amOxieOzaX/pcxALXYMCgA6+vbseK2++Gmw9
4GNRRZ8wkNdXgoPPnv5wgsuA6uLmbnmNE3VO/PIbjnpDSvXg8zp4TTN6/G1XFsrUOMFjb+joZ/nH
SkAid1Uy/pzfB2lTWUg0netp+N6wzgSClDhV3dHMVKagMNATZN5lLY89E3BzJi6V4YgfH3hf9gzG
YHDX/if4wcXprwQhF2t67YcUAVp94KVIgb7WPVk29Db7VW6CaujvMdZw7ONk7VqfQw7FREWsF2Zc
hXYpuIbJWwZqdmP+9eQq9VCstR2LqKegABrSo37CtuvDJJ4lEmH+HZQOlWSJ+nTxW8JKane/a3Gd
g5OhJzo3DV3SR7y0PhKxOCoFWbQ6GeH98qo2QS5FZaoZv5pZJhekABp7m5LfcWJUwUTr/hPP2re1
d8CxdEHj2QjWunbrA5r1r4mLjDsfFA9Zt+xrhIJd8hvFr3wmQq0rWP/4MxHYZx2AORR7LFl6GCy3
R8cgIekgPK/3SQYJhdQMjK3kiy+K30Q5ITjmlxbAjxhOu3YuZXEa87lOlfhCgba6/c07tmGKCLte
X5AxIxfIt7MR3OjTHKCCoabAYy/qG40GeRZEyOvXq8/H9AL5/ZoxnOfdVaOm169gtZig6XRdrXSg
IJna29Kmloi+4P5NtmXkHrnJEtHJPaQUAZjMzHNIw7tIwCx6OKS6mXusd123tQ8J0J/Uj/vibzcW
RTj1louKYAttuD3BHnmGgLTF73JNgFeRWMN0O9wgS0+PHgpIOw03u8ZCDzO08/DD1haHffRNwos5
aBAC7LEY4vtGS1RS5TH7bKhyfPvEkICnB+f1G/k0UURm/qP/VpWOcUvM4jQuyibfOgznNLxOMhaM
PEqDAc63J0k++JoUbogS3DFNoti/BFPeLejs3/PJBFfZCoaAwkNhLRpAC+Jfoankwg2FIP6YlLRp
AGmca2UMrP4336//wk2j7ewa6gQwrka9lUVX379BNsTEIDVJe6snl73ilDJOuJLYvL1gVY8wDwvo
6iNsdAzSFmFCs9/lbeO4xmHYetSABVgNP9sNYDamPH6gkXyJjdMoM4PrVWGxin53ztEryI4mTnDT
iy20KQxAQOruNrVXXhI9wTY7P9qBVqJ+9nat2LY4luBs93B4PrfGIlqlI0lSuYgUxNXuvOyMLBb6
Wm9lQ3aWKj/875mPr+NNmJWFQDAxTZq82A8MYq4aaufmGFaKWZN7vDks87XZA2Q7HJfM4bCEdWKN
uNMZljVuZT8cJir3epGAeVLBJyyHNpI2p2ZHz8fguuN5IZuacti4SAI3SlfmTLLY/8MrIdcU7QJy
xmhWjWoLNaeEanTu9csWOz2rPeX4iDHHLkjs1gNYF8WBgPCg+xe+TpmIoRMROFikB+xdig9/johb
LE8zbXWRgCOJ5LtgalgBcEDAaYKT4kiCpS2HqlC+v7gTzgdO5/T3SbZbXKjMSwnxv7jqGoPt49K0
Vpv+SfgSP89epuKU4/6J2yf9UBmX1kLALylby/lqwcz4Od3rbEbWbtWstwMS6XfjlZK7cLCHD779
XH2uodMepWg62lWXu6UK77OTlOjlV5qVsmBrU/aUeC3qoCctV+la3BFc86Rm7qRa6ZxjDbUW6Qvr
ylqdKVPbZFHX7Cc37rL1Kzlm6NRJ8Npal/MpEp2lfAyNuDnyLRJ1aDqg2ar9ZFAx1Gv8ZVQ0lApx
h2oI4TGlTP5rIRlpDdrto++fmulc3w7D4gzoqQrFr+2KYl5MYvBfiNI3QBg0nmCb0IfXoMV+ETDW
LrFFnIOB4YZSfYhhkYVMA0umGX/dgN00MFqgi9rDR2/ua42dY6DFyQmXs1PsVRns461etwrEGOO4
YulEJO2CWZplhKbXht2WFnpCu8hIIoVi55JUG0d7F1PYUz5qgkboWlfFZ+JtVBow/dHDNsQc/5iK
AtDjNrjFRmBt+/Hu6512ogNHZE//h7pxyrjQJ9Y6rhL1Hp9MNB4abo1mIDEsUd5hMl+CbqPVYDhN
qG/zoUtZW1S20qGdcKHojrQ70iYLB++VhHSH8tU6SR8JoRcL8T9ptNom0omT1vm3Tj2K0/LdK3sV
C6ajJZaWD06vv3qWsMNhzkTpKTh0RlX1O23WekptAka+IjXdRzXq0gme8Ju3svTSjCWU52RmmREl
i/svJK2+x9/5ct8g0uiAUw+qbmd14wEpg2Kek7eJgiSbYqL0EIG/3D22NkpuPFH42IGmNWYIIoX9
0Vx1B4Fjfjd9aYp+Qc6MZj07+tLvHFaIDWnDI7ld+6ROMvBiA0jB7OLpnI9wN66x9oV/RY3du+td
nl93DIzSbynefqsHM1hfLHeA+D/KPc+h1FvQ1vYgYdMK+TGaNU7hH6O7uRJ4WPB1/npWOwl6y/QK
quVzkqopZqbW1UfgnCOB72OLTu98CQayrReL4Yuz2hMgdRwrC57jXEHQf0hwqnmc2hd0oo70rElR
8GfaOuX4161sVjJ+KSQiSbNZhH97V15SwZtyB4kWh3QJiyivSsnKEg1n8mmR52kOkzuf74v3AbbF
CgQpSNWr7nhoQgjq+XPr9bL4Ki1vdpR7p5ERo48GRb4kvKFYW86JqhcET1lJEgtMHjX709GqyQl9
ADkGo3OTHAs5Kn43Cg+joaqmT75zt2tYD/Hg7AJc8troHDM8YM5eE5IVlj+eE+bO/8a29Dw/lUrd
7GSpd1TtgOzC6bLLxNFFRJRAZW4BGI0F9g2U4JdP6X+a2NRuuDFxbzKQep6MTrHYmbL5sVszJv17
9SVu6uJJMN8ywMf+X9Lk9dW5YU+cYLvEvVGgG7ig2sFwHHtQ+w0E3cty3YYoY3vqUMe2mon64/gz
/lV4fNj80lBn7Khrsa+KsexqoIpTwSYBoe+RjHOTqwhoCwBkdhgv/2tEZvWI7PQ2Ju6t/3DAL9ee
WRLN530nzJxr77YGa6g8FfX0bm+LipjZUxNz7fuHPKIdyAhxd0H4WNHfF8Veivh1Gv6nRKs8Vwps
oxpZOtFSTakAqd4InBgiJpBc9w7O6wzcLXDS7LPPtB5NVhsu8ps/jx+sy24LOmgPmz7OvCocwx4f
asht9B8FBqcGpMp9LI+4+l82QWicXLIwGmlrtAZXaIJG/fmnSDVSN2yZDkuQpeH5wMi/pwENniY0
hyBrzMira6WKAjGfyC6t4htlukjhjHCpJEcaAdGXowUzO26T5a+HlrD1XK4NxPaZAATiEU+Hjoaj
WiEL85cYzF/owHSCGBd6+1YRym2+hPGlZ9svfQtBCMK1cHuQGY6aHAtHSdfE/zUbQcdY67XoPVkQ
y8YFElmF62I/apHVa9ZE82XG87uWp6iuZBgjBeuXDZ57nFoIW/fZyJNOsNk7nQ5v0UcTnRw8EnB3
3NJM3XbuNhIbXQrpzzvNpv7Uk4O3LPSsLRdgbLTiA+h5BXt/gU5+X7bIA1fVRYih+I42ILEGgs0X
8Hr8U6TSDozdMv4uKslXO2wQA+0LyGf2C+97VO8Lgo6NlOKEwl2uLc3fdtn/Z+s7paO87sF0bLvw
i/+F7TORxzoFJBeDRBURCxsNxHroTR8FxcoZGTEqzTsd7Cy6vVlaF8FYu2ux/lU6zN3ctR0wzmeO
jgApMNMxv0wKXIjtTqQEXZSmp5Lj/hkXx8Mnzn55i40NMzT9K4cCernAlimimtdKaNEyZKAYIt1M
tKhvVZ3t8GSMDMDz9pFssfb0qrXufwCW+BKV++WMp4fKq7KUsjO6kJzJJ4075XJv8+zpwcduaP59
+vXt42yXOppCQ1pL7JYAZHpmabiGQHKME0OowmhHX8mhdWViBQkssGSjVwS2RCIzfx/WWKA56aIR
j4sk/CoC5QFm7nAior8tYHsUr+y84MbqeDkHe2a7ASA6jp1RrN9Ei737bmBnTU00Zh6hwFnI7Dda
mlD+dDz/akdISBRn77yJ7y7dIzg9j3peCGWs2H4M/FOUbX2pT717N4v+kwcwaTIcUw4VsuFlbmac
+zs1t42o+2yaw1zqTSnUFCv2bkS7HSZ6f10eLhLiwIdetrUqpx99+POUsNkQ7jZaiQRMjc3LWq0D
cNMdZZmfyMhajpw3YeJUBNd/UqQRzApHNqirA7VvSbkry7wP3dkkIrTGuI+BaqqoyxFAiL9wtW/f
oA9dnfb6qsHPYnl8ObcnuoAvJ5bGij2p/jHPjy9vwlR4EUhj2xgCACt0ZAAnc8ApSIfpGUNZyEja
nL9DQ5PquYNgs197VLH/XnPR2UX9ezMEjQtS96+66/x5gA5Ka6tgywrET2G5js3zJV6y5RtBWlzB
HYrfxUTNzkXkVurcwZ4IE/XZbj2JVLd1dlDZiN8TTWwX2qnXxttIV8xiDcnzj4DKkf3JRCI6wr9t
Ih2cAjrcPFmF7RoJ5lKYix9GnP8LO6xdt0lmwMpsYDnK69UeMQV3vwUyNw8XrL19/u1ngZWQR8sK
Ba+V6NmR7XbR+DNvedXzY/JXVGaQIM8WzS0dZYBZXRzYgBHUhRk2Jkv99X7Bd/FlwU9M50Nc+YjH
awz0PKRNOLycsXyD/CBq259vZ4xZZ8jlYcqnbqzTzF7MSO2iMfDm3hW7Sm0UB9RqhOXRcfPHNYMB
1obh/GYRgaYQ4AcgsWfDX4wVHex5zd1X3P5OxjyQr8upBvrkR0jz6VSAFxMidfVGLTTaB5FkYrkm
TKtJTCRvueXhOitQAFjW7x5PjqrwJx6jWao4gFCVdWHbTsoqihT/eEvz6Tighx4raVWHYqBLikqU
LYn+19cjRD6ei1EIrA4Qs5APVRMZibSzVqNg/7MpgdbxOcUafRlrSKZ2iZY93QCVw84nxDbPNvnD
6rj2yV9+g5eYyvz4KSkDyeAzj7sSmiQ8UpLC1zgHP7/visgWiAXXFwT8MqIOLyXmzXTkw8bZHaH0
pzF5oYJILvlgdS3v7TsKgwaRZ8vMHN+gF3bixxDPlG46gVCxagK/3+dXiXTazUeAF3WoHSvlcW6w
1c+wX6XxyLCSvfOwPLn3uch6it0R8GiKRunx/VQUajW78dCXqRVlVpfJJXVAh3VL90TsXDhgicm5
N9SaJVDUWpg8gExGUWUOA4bEGo2lGYi5FY1d5fvUwHs++vweI/6s5/ax0RgUc3s9J7As8/ZnTXOA
3B7YC/4A111vTx+hCKu1DZMEWMrnQPNmrG5/FfajKdGEwDUgxJhca1xHXKeDZlZDaxmH5RP8lQMr
FvvTo5c3Y+37wP/TFRuVjnpCDQjM/IV9GN/EhKoYyzJiq2LToY5i4RFiyE3YM4lNGIo72a5wi69h
HNJlMO4LcOXWZMp9+eyOJhzBpMGrLsysKgekypCk1SN7R6XvbFEyIDaguICSruAxX5GJpwGM/7jo
rJOu5vYPpSxBdEJRqrxC3/NGatGy3dCqdbe0GIEQkA8ZuW/nYagFa43chgvWAX63pQ2TMJOdS3kM
xbe8WAEWJV5tkdtyoBqKze11OcerC1RVs9Tr7KIV+i8a+9pfJRfjp9I+3zuFFbAj5oSLX0Mqi0Tz
FlZCxP0WZT5H9vaDcQqkh45giORBa7LdccxlkLk2CyC8EbO5k0oQE8+yGHfJuCDy0fj4aQdrNHUE
4qqqiLWu2w3hp/0A4gBuJsLJQFA27lzDgcxq3wRr4WrLjS8OQr2ZF8GWVunt5e9mARecCfa2Y1y+
xv57WA4pe+SH4Sxng5jddCM3hmlxdFSFvpOwmhwnHtitoGeUrBlVLskmgw9bingJUZVy8tVedB6L
UYydG3PIfl9xZO1o4fWhC2m+2ss/E2yVG63hOq1DZWPq9xYf2lW9eeyud9KegVnm28VPzq9uYlTo
eMKhtz+wieBTRDaE6JLj0Ci7r7i5TV7+MCtQ/vzbhxpmpQjhll962ugnIO8pvLjjJ93+a1lMP9fH
c/xB7oRzUqEXd9FX44uSjiU5OqSQpZMiqefxBlt9TN9qPKbo0jXiw3pYWEKR2ZCY4T9gKY86AFit
bITphMW6K5I0+VZmzEqSRm6Y3H4aTOcz+SSb8gcmlFlX6KUck7S+jJMW8NgwJiXKhUn9FSFXnn/K
af69H2IG9GHuGEa/h1deVGtOaK0xP+2jeX0m78UAEdiswUq8iZ6b2rw19+3CKBisRcJBiblPXnMs
ywQ4cc83uMFMPBlv+a48BxzNrJaHiRDolVQQ1uivQTXunwaUqc3CQcAAWXfP9dRrTObQj4OGaLEb
lm+dWaDmU4WyfdD8JHyaR75qZQp8mv2l7swPI9Y0xXEo8wsgn7xf+wTRcONNYwoBL07Qk6nDv1gA
dftKD2pxd1lS1TYp5m3QwzkdfqCdW87iR9aIHlSZtWko3Wlg016LC2VCRxXffN9d5cX5YuTje0bK
znwsZWMjy95LpqF6wvCUgCsUoPmPsk9HFOtt6qVZbVyH4FNsROeFeC9iCfE5x4jdOaDv8gJVu23J
86/LOnAZPfaCJ0Hs/SLXy4Rmzs0BirU5tZCxeh9uuSx81+omLbcgMJaljGXhi8Fa0rklmmUhbStH
kgAAsQlfAG+UFHvUJPAATEdakxv1jhnDB7g5OhaMBXGwzQtv9WooOMGFQpx2MY5ebkmEodbFoZSz
qYL5xWakTXAFHAigbikPeQ8nV/imfxaPR7e+olDNIKcI2wKNcAo5gz8OEa/1ErJAKB9N+CdaNlkg
3tu1/BL0CE90yiTyYV+uKuFYZUxwCzpUgTXgoP+QC59bl8rlZz9vqtJ5np2WTYrG5b/dEaKQcIKR
s2eBrtq08sezEp68mduWz34uB5poUrCQDIas+kCv44KZNuqDC03LS63of3V2Yas5qoQ/PqvsehGm
PHvEvQn4UYCUYc9LDju+Q6DyNqHBBmZEka1ziLjgDf3k6imOEFNXp9tSVqM7yB2f67FR/zj/VAim
7L/UA2lHwRaf1VwXlZrkhJlRUC/zziRxwL1H60esodBgQcpYM1jbUCGbOngMpVi7UTkJxzoqBBGd
sU+aYtxmuuVysdeN6z3q+jvRJDy11T3SN7ZDnWludZmiIHaTRpjY0j/LTIYdtOlAD/RskeXJ0ABI
Wkge0qJqyyGUW5aKOaeFQH6ljUIZN08t8w56YEbdoQH+N49J8K1G+SUUbzEBfr6KaNePafhfLFh4
S6ZZgSZ++0IE/iy/dhn8lYrE4m9koK14/2nyfKLy2JcLspSMGDhiPf+wAhISLMV/Oy1TQnyCxlvk
yKyx321srslr9S0oGsi3kUAsyqaNe+kb/WzOyff8jlVWDOwlQKgWQFgs+IBxqwwp8vSFuIpn7SIZ
A0RCtrhxJ1OiIIw2irxz19845MX0+fWRzIBHPGM9hXGPpVZs57u9AFe+oxereDds6Wldmm2n/Mhy
3kn//KdXJmHo+tAFtjObo7+QTnLsw+W5FOad5A5TGE8ENY229vhJonWLdt3Vo3462ZOs5B+Fiha7
gBRFjazoLdOP1IBf1IugewiTNkRBMt7cVk9vf67F/YI7hU1mxj4U0QHMLch+uS1GzfOoA4ujXQiy
W5Tc7Hg3+hT+6T6eoGdNVnMn7AaQOScZ5B1n+FsomSIPog4dlY1bIWLq1ftnoGn2ACujWiGiR78I
pGJxMxLEnMqCi5ukEKSerTcJDydeGnd0lWf7MF+a9pj5g3dZ1pso07bWTOZ3TQS9AE1f9cqs2CPw
IEAl4Wfq+gy89sy21ahQQIcUb+6AA2bwg5j7NklH9FMY++c5+Mw3wEnBVcXRwvAS+1trvJCh6PiX
iNoPVIII/AYCBYiYpTHSc0bIADT2JLcBWmOFBt/Ji6A9BxJqTde15RCyEWerrZUxfUvTv/ZgiyiR
t/BegQ9tMawoBU1WlN4QuAyJc9bxklge/E9ys4pmf4K1Hn66H2Ww426PZ3qnmnP3U+3QOi3O6dMv
YpOyi1BWxdhziIm8vTqsSdo7BfYbW/gDx+TscbjW6QNsie3BVq32iJkPZExlm+mTT8maW9mP9SJO
pyWAyRaD6l4g2OdEeVU2HKiQSTnEiJ5FQNgMX7rchjQL4AXbu13bNSuLM7dV243iVlAoGwnCmt9r
GJhUMpzwS3EJeIklFyLKcZFpeFs+U/BPKN9M82PZORewKKJBIniFo2L2rRHc0wWynLgHw7TcxoIb
STG+60hfAGUFhHUkWLLYKoxVbL3iFtJayq2HcyjtmFkDt10ltJG4oM0rorXO0mjLJMyyv0Y/mvm2
37oyZLcooRbfQzLE2G0sSSiIFf8aspCSVA4kYqMjnEfxfS364tHCMVICGCT8s8sK+M8iqj0BUWgs
U5g2ASt8QdruhZ3/Y4SRbbeY4mjndqsfaQrwib7TBGSUT3X57Azg8EgKQLu9POi31xHytm5v8SF2
Azlide7m47TdtSsEhg6/onR3UhEMTzP5yn6RkiZAFDhdbte5oamX++zoChnsJYXTNEMuJOE2lLgH
cgNqBOmtIHCVnfefUkYvJ/kZj+KsJuHUGVZViiG3hHD5g/ilGjecat8orhk99bRma/MzuZUL+HF4
/Ryi1fxsuEOw8zeydTdNvMRs91T8TR/77IV0Qhs03lOD6BygrkOm7cbcGuSq01LvJjw6uI5ZTNsZ
SKyz4/7I2fxjl+GqBelLXbv9kmB3QPXdv0i8R9jW29vRGybDutf13HA/0qtUVq67PCTmE87DtQJB
3WceIrMFXgjAiP9PRHxA/dQvSnI/UAuv1FQP4LOQUFukyNPASnQbYCwaMWKzIt/c6T0AW330N1XZ
a8mlqbgg9C0qrBAOX9aE9ujznPJCaWqBxchkT3V2twGWmWYmtKLxrjkVAi/n5n8Wx1LuqHOsN5hH
bJ6YrsyClkNyj6DG2OT2jQzw6zJ7jS6WhsI9mvnvz50OfQGyU789UY2Tj/OIa762EGfpqeGmFRrp
StGS2kghCDrxzusZBc0XbjCHoci8arvFmhbMR1aJMP3tsXAjYJ9Nzph6Dfz4+C1U8I0tH8Joxuaw
NRo0GUdtCm2z8+9YzNHEcckANXxUQ2o+HJ2B5KDkG17xXPRAo61/njoPPfhsbxwGOcsTPnRdKrvu
lIGOcp06wBLc9EXTpXa3qLBZDBsulwGhR1ygSW7hKeTR4HunX/cjSk721SdX0ue+lDvALT6je5Z4
2XE6J8SxiRc6xOIZApQRKkcKP8Zt2sBO/sx8w3WKv2nUa1pTV6UvbnhdzLo0/rmd5aa0C6v+2Gp9
99CFPfW4JkNzFSZ1UxE/zv+U6cF2BsaUypazMAoxCMhQAkMdUIzOu65fh4cVkDCak+smaqaKjPl1
OTYofWdjw2/tReQpJYk3ZDGUr7jLNsptTVGRXVQtvw/UGsciAhKpK1mfBbsuJXlLJKDKNXQDUYFp
RlqEWRKVGJvphy1SYpoDEm1SneOMJOMJ/1f1GPvlPiQ1lg46hFCLJzuVqRp8KNqejhgJqjCrSF4+
d5ySOlKmRPydADAb8QU3wZekv9RwmazhcBxHNcIGgQhp5rbj1TY34PTTFbgzbfEhV/vCs65sWsWk
hW35lbvNwtqtyMZlSnc0ctXQbagwumOYLjKPCKatIVxEXAR8PI56xW1+Ria6VIRCF94FAsoqO0xw
s5mwY9Qgy6FL2ukunpJjntS+ivUX2yU5xLBQnCpfY/W4ScoeUitY/6VLEtm2ScKCZ+WafAxdTcm2
LXiioBMLLd+DabDYvhchErxXa+wTjok1lRbDexSZBGOTDpr6auX2Bhu1c6P1LxOAr18IYFoYsdAQ
J3zWjDaXXMtSXDz2MhYoNaiEU3A5O3rYLZHUvoBuRIG1C5fljnVShCjpJ4J28cN5UV5R4hrgXebq
VeWEAK8VTt1EwIArAhFepWjkDn0tjgDXT7HwfTt/WKlDTKRLupHSeTdMGO4cruxA0hNCxehUMTOc
063oy0njYfvUjXt7h1QzEFs/JJuKFWy6iyv71UyMs9oVUAuWZ7zaBSoAAJiHMGObjc0ObeRCByHJ
7VSNsUQVyZ0Uwne91k/Gq4m7GYjdiK0Yi5pFanOvZcDXlFsT3lYw8hVWvc5kbVCEbZrOl5YxQZzU
ziSNhgkX0F6RUoYxELbdAV1qg1EUc2QoBMfjUklNUdYKona2YIbwS2eCl+/svqi5SwwDm1OQWt5Y
oL/hbvtJqhheGAZK6yzvs6qOC5voiFWCAyQPSsrI0y705WDCWaPEQlSdzq/RhaZxoTwKRGD6UATR
Sh1nGMu32UenV3+ncsOk4ImMmtf/gFObyP+aWAQSuxKIx/e9U7opDqXtTUyPwimSWs/Rlv2Vhscn
rl9ri/Y3QZh2BM7cv0WlfXd2lLO9bFWm3lM7PW7F2RSBao/vLh/IFAWI4BiQfnkdVljGUzhdvqP9
Eg4G1y7lAVfzkLeWo2XIy0wUvhYAsSpN0KiyMfqQunEiaoiB1camlQ71mIkWn5Pa5gjZb7wFnDSL
T0R1OJEc63stolAgsIybZZWH6oFKpi7klwyTRGiELF+57PXujrpU6vnQMLTbnk4HarqbWGCjavFP
G9XHfZVczSB5hRT1zAoG8rC4D9kncWqfArWlVIq1HpxtvHFAk2U/E94+gyJx32fDu7XjIQIQ9djf
QviGN2PLU0ivKewdCkIj7ZKZJRGA3ue2SfGcrBlA2u8kbtDBqQx+VLCKp1JpytuxR5WPTTMbVLga
ilv0V6WZzF8Ovlkv1NVU4CyhyEsGWifXwRjX54EtkSANvcLG+OxBpVflKfnLMQRao/qARWinzadA
yEesdUO3wyepODlPMrqeFkKojGMAc+8bJKXq0M07YhE5O4cOVn4FJXLEQIkpy7aZMnANrBCGun48
x2mbVG4B1f3J1QBr7zpZxoT5Qc/y9WM0xfnOFCN4n5kRqss8YGnvT01zGyVRkCn8PfuaLdlPJ9I8
KQB/J4+yp85BiRqwdRjMXFcadIUQ3g9nCY5+4ZV51f1bLzf4I3svfT2mWQKRD2ov0Sd5rVbZu4/3
oTa1FFt9mlQdZfriOejN6PO6gD+d+X5VfIH1Hwu7HKAvrsDklaupdRK8JR7Ijtz8Ybm2UYoD/MHs
6XzGtJgKDtCK6+Jr2sCeYjXqNMIT9FHW8gOCKeqOjLMFczCQ6BiJx/ugfDvp0RBtMk7aPT0P4Mmx
obIjS06G0dU0LocnOHd8q6hFzXmAb0/GmA859FjqjdCG1/Uj4XDCtacfj+SU40zZILHfczbxShyb
BVxJ+CzAGjIV2dygIT+V6In/b7nZmoEYxC7LM1Hao0q5fypF5s9c5AsTGPAa2oNpuc8re7Lc0Wh5
ReWkL3ytlnecGgGC3kR3EMkFY//SRp5OsoYoUsjJPJLc6+Ud/4S7YII8+kFkk0YWsmSdL8Xf/bi6
CI+bZ+3nLndZQMQ5M65ArDkOdijUZ6XIQRaUWSGG1EFWc8YkvayWlVXbY8KwlCzAm0/Xz90hkpsk
RpsNm2FM37IpHkWiDxFeU+bzkV4L/47PqMksEVmbqKr4stI6EaYrZByHdATvKdLbMn2a+G/fl3H2
cNRVWbc4UZFrGSNWSrEgyOwXxSrWOG5Xl3Fa+EmrVX71MH7LKOOykPT97LIFL3VQnCu7rwz+zB2c
f2D4WwBkuF4GGArGNdGy0dRUR5CgaLrUtC7pR0//3bNiW4O0pB1C/xWiXxBdLomVa2NPNvqSs8Jn
zlGxJbdF400RxrmD1rWXjUa3P6vpCdAdy5tQF5++k1JPcBP6TkJThSwbNkrfpl7mLh+Dx3qfXrWI
AO/MsP6xNqK96w7bH+EI3OJ7TgftMJ49tSTr3EF710NUQ1TNaajljfJ71Ek9SVpN8Tc5GHHY/GVG
Tp0vtmJ4f433P9T99HJIlyEs0vSULzP++u68OwYLxm3USnxxCpB1BVFK/05+R9veNO5ZgpN9LIcd
996ICxeRzvXJ3MSWWo7OeRPW6ZDUSMiIT2WWO72/6y478Tnk9P07RuuUqPsHAq2cjZikxbAGgvv0
02GtHenWJk8mlA0ets/KEjyzkb4Jo01ZYQ+Tll38G6WVsPqg03bmy1avaO6i6BHHfnm1Ax9KjJF7
Qy+EaDblMF8jH+17C+/fbFWkE8w4XpKp5SUUSNRFQwDlIeSMTmpwRqTjmZ2m33BKBqISTpG6MltW
Tl1jMKGCn96GcBwR/KSPjezHj2l1yKgFUE0n9qT3gqdBd6LwbJbNFsNaD3kJnzvAlgDOItKkFl2T
Bkcb32FOuoo2SAoyNVxpSsuLGv+GBF7/8j3h9tVXtN2H4wzBatRkUUQQHUUlduTQl0Hz8FuwEZuV
CTTKamufs0s6LIbEHNGeEVsZcLbkrkYOdPhaqnrzHvl48HdguP7B5zeu+rCbIJhbXENuZ1I1u8c1
efbfHpVQKp3KbDfd0SGWzUZ1dk/1PFz/o/NPAyXIhTYVARx5HD5hKGjY9LHIrjYWEPl5piS4MOY1
xY6sEOmi0U5BpsBmDnEzEOssKveDZNSyYU2PbZ54lOd+0AtnP0OJNQPEdgM5LXG53LkdDhlAL0Gs
ew7l7zLRBRuZzPvb6mVKWX/gNbhoh4hiPsuZt3vi6pSeMzHUPDEQvpvgyzl5KbfCLaLN29qgQdse
b61dIpM8BmuDKZqmF3VSX33FyhesH7hm1OaGDnZMLFcx6YpY4AFdV+JcuDZ8qrmoON1r+Yr6wd+w
cP5eFpcvoiYxRKuohZeTgW2SzDg7vgsuooFd2SubHZzag3NkXY5Odt5FqGyoFJkR3vKEWert7lf1
s1Tr7ZPDiK+XZt2SPofbouIpSlo1rzAz2r4qyUCF1LHZggi1/TQhC9p1AC9vUE5Wq2yAaffZsWyt
Ec2+qKTBjSjPwV0MueHtRcGdrD81Hiv2p71gGeddAyaJCN4LwKYncBhLfUmglSFSXWnEhVnNrATr
cRaWTx9uOBALwv0rLY8Nkeesw54fWoSumm0PrHb7v4Gqc1zTqSmV8aThtCgROEv0DlE60OXmrgiM
1C6JpSFPGmLVJOAvVQTc29YANM37i1Kolxx/JAPlkzAiaN4V/CeGdkbqWohXWT3AIewDj3M+FcwS
uGH4SmDJV618XQqK3mWKIr4TM/5DOV1RpBGlG02AO3AkZGaxBPJ9aVOq46As0iST68SVOrq3rxUw
dWWbK3/hrmA60nb+7hFuw2I6LbSEA7CQhToTZ8YMYKgnhZ7qkseN+/9P+WagakcVE+NurJksr43a
+zAD8Pzr5NjXgj6ikXJjHo7yV2OEg2qK7BScTJFKNaSZz9F9LYtqJoxuW9BSbI8p9AYLtkJkEy2h
SWnN7A53LAYTIX5mEQwUK9X3Rjt5y7FTyUcUzGRuHRQ+Ed7jLrWL7AbFqvTiyQklv+Fy3WPr0H3O
yIm1wxPdkHvguVLNQv4gWg8bB5ly+kFSmv3fqjtRO6j3cVBDKBdebBv8y77c5FcVSAneN0XTAzrc
T/MMcXZGTgVgxFyTYoNpnq/9G4TtvfcJMzw4y7O6IVIf8PcbY7mrFD0vEYlBFJU7Fc8gJ2mih/Wu
6PCRmXdVBgtIg+GtgyrYQgKmyzCxwSw6tFJ0n0/IM1fjtTPLlLp400vpbr9l6joWEKihZyG8y2i8
c9zmuNsTtzH8EMD92e1nRftv93rUIHlI/2yAeqR04C4h12dziHWQRpsKDMEEholpHhNOGo04Gxlb
8rg+fpuXr/lZdAJW9RyALmyZpL+klzFoKftDYLnzE/xIuhwYw2/xw4psoHQlJSLZP+u+Szve6AgJ
XSQwc6Y64lsPZzD8uIf3NxEyGJlCUWtoH9jQXLgOl87N/AoztM3h+AiMBgEkzpxVkgiX4fSvLvLQ
CSQiZmPadCFvKSyVJWnNRdjycA+Pno/iVr8lPoYQpSZ/ieoWSt+BNcshL/X34xHalmiAPAq64Jnd
+0PEPFZBzIY0UMKcFXoAIWe8DcqF2D0vSPLAZ3MN3l56F2gC1TXgypPpOisbIlkqnvtMM4p4Tx7e
nZ+qE3Htzs/6KhjaD0LnB2+li77GJV7doAhJiXf5mJ14O635HDyTxU5RL0N+bqOnowx418XhPJ3c
rYNNCztdkhBJUc1bED1PvDhhV0MuDbyUP7DHWCxgSL8wMmvYJr6F35+WN1x6D0lsU0Fxvyn8uJzL
YSdhp2yCjWHWwE9eDTfyhS1ooBrwxRk7fYW+28nFr59NfTnQdv+EwAcPFrORJtReywESc+I1NI5w
LVlpc2tYprgGVXInRceweWfQ4dZ+M+qC+aOsvXP9FpnYg34lv7y6J/oSxnHjEqEYrnmE6xVSb4ZH
9XkpjGl1ff+Pe45189BV3dY5gQUpica+GBuTipgKShZWtiqHJjqy6lBJITMc34BA4b0yPgqYyeAz
vccTY22IJSZnk1RZ+gCEK4DiyqqVfJG3UH4w3dWGpkzjMFN0y3O+8EWPoQ4WUAm9xhGk+drQBNXt
5LDg1RjG++y4uqExbFxfl2gz7/FFNbXkC247kC08pAGx18zROVMZbqA0qIgbQW0X4Ak0yexdqIrl
4ixuxh6p+gFn9LW3idyT0t+aw/v6uVEq/JSvZ6GHLI2lrZIxg6fWoZFMgAMFMlFu5wzZ2/eU2JdQ
wpvkVMQidLqb8yb+pSF9mSci4S4/6dy+RN6PwXwy8TC8s5aWl3sjjSbCJ2BYOPR1l+yHTgJlrr8g
4rSxygr20+ssrh8qZX0wqYDEftOwoyOCnmJTnods9KA8ehdlwekCsATEM/k3f2iczyR7m2gdQ5J4
9WTEXtDS8VoJ3fCrytU4SXFoHZ278vOivBNBxI0pvlOYS4LK05ul1OpS6Cxaou1yNXb95CX/FGH/
uJ7vJm8AEiCR+UNDjeaD3qnCv0waE9tNHvRP4L0d0UzFXFwtYftzG6MHTxqYvm5NQThrj1mzX4Nt
wm24mrTmFnPw04nbXpHLx2zzK6OmkhBqV+P/8o/LjXJtib9iGKlAbEYIEd+i43hhv2rRzCnSvfIo
EsCdUqQbNFGy8QmQj3HbEV3o2i8yaZ24O4FsOZeNavYR+XccO1v4xAHtpC/y8X5QIFXRleTnkfe5
oWAjW+Q/73VwNhjiBprp5p+b5FPnG63daV9fgHHZ8LdFZuV14WfC6RgQHUChjUKE4XL/JJ44fy2o
1BLoVKdx25oiMzhU1ZwCE0f/yGI314fGfVfNEcC3YZLl/C6UgrnlAUXoR8fow+T7j3vdjQ3/PC51
+kkg2j7570sF+QOnTtZ/YWFbMCd58k5I+/p0KJfRzgEVxmFow5SEV5Hb2LXjT9GuGrzPj/96+qiJ
drgCeJK/zurrYJM5jP5+CrNtfomhY3QuPpGKT5AaLXi9YaazMBdcwPDT9TbNqofD1ZVKii2YX+Tv
R6nqNrgT0HAukbeHtBGterihWS19yaMc7uExOA+vk6C9t1jukwvu8KJcIcHTn4heBujPu9bXlAMn
lY0K0/tfm90GWqkEvu5NwzZ3amKkjKq/EJdRNKegCfFGh3E/JMaqtoB2RE44haojBHGgTeUPo8qg
wcwyK9xkxYwWHjPKfSLHPqGUiVpDoSKKQVWdM8FVXhewCOcX16UyjEeZuleydkW9tdvwttD2yAG/
JOfI/tdmmS/dBJ4xPk2DyBKZSLe0OeCoPmOylRGTb1JBNPxo5canORIf0g3dIO0VZvyxZRDo0k5v
Zm+i00Xq7irX8zIrW9614SRiZlm/izE6EinHWR2R+vt4Gvag31244vJrykuyPgoYIMkpzBA8cmp7
UkMQXQX/vULzXB2NTEK6v5DDOHMuFkjRCsRBXVLqMEBabduMkMnDyNP9i8j+T05DGog3Ih2Nitqs
u5a82O+lilXUPzNz9qqvrMn4QgpbkiSazgYTlm/YeHq1DK1BHv6csqW9SNYT/ZUHBjmG2Kw5htk7
AmCCnWBREViPeUWy0FebfkgCxKjPVxcDaCvZ9E+e55bhxIveDOSCQb892KAnjfm/gOerihJFN9bZ
FDke9kdwmqU+KNzcTdPUkPcwm4TIkacRMdR3hkaCOAcLKm4WyGCua5vhmt+tGAAKPv1Cq2vGnFzu
KJkeSyNR2E5hs4Mv99l2oMOQWCbqgCScVK5PMupCt61b2k00LK+g2QaEcg1vdEVktVjU6TbvjOjW
Gzwn1SeZWwz+bSZTEigDCgb6x9QGRnOSb0YifztQDhKnDrftfksL75AMOnZakywMpjRbl7wIgFPX
0nMsjnPAc8UyCtGK3gioUgMpIBZ5NG8HG+JKiEfzOJaRrQnbkfEepKf3kyCfN9YXWioCKV0QQpGf
EcUkbc2e0vIE0KGPLqN9xT2+mSJId2Xd22mOmAbvc5LxHldrwUV5ZoFsw/7Bx2dcJHPhyDk0OPzx
hwZDocXhSEpiGsr4D5vzoGR4Z+/hlQnSBuIfJwCchW9UDYVsaOb/E0yNqaEbu7bg5GZXrxTwhCP8
rKNt+0BJbOdHzRPoby3zMSH02EIJMWEnSLKKIO9fd2vJEJhPlLQdC4jEQqzOKH96xiUabzAw9xqs
P+8UNfhxA5/GzLt3PauJ1GmkZECRdmmNyu7JOU+GqomKHOxk/f+qjB3ww9iwarJx4zXYwg3eL5qL
Jl6RQQtYZodSrCqyIiBIOi9feejI8HsO4O/S6MaLwZhPIn1cqWugvt5EzqKGcLfADwEPjkqsjqBT
rA34g1OO8XiWO6PFmDRYodNsjsLgorOwkx/rLzR89nucC5Skezi8zBJCbPG1MHCzCqWuyxAs35ZR
DgoAoWPJU88K2QFeIn8pPpvFynp+eKM+U8/LAUooviQBPZthNjzte+BYc0VWBxXsizsyrYiP9YH9
brFByceQBQ2waeCXrpDyGZh7cjw0hqI+WCsGoSPB1JVcsvig5QXBQJvyf29T+schvbhGorU59SGy
j3XAE4g9JTpH2NoCIWUhh5d3T4XFAS236zR+z3FvJi6hXcKIa5oSQAYbHKXAN4pcksmfAOuXqI9n
eAVgHFkZJBXXCUyxnP1eH6Ukr6F/5I0kvch8X7CASmQIoD6rMEtm//UFIag3/zgOJhYMUPhZ1340
8WZceket65G84WD3kpLWkn7vr4XQyqAblS1qLJaZRm9YGaPWwJMO4HR2KOkzX5eTr18moYB/iJu+
EsgV31EKybRdretF6OzqC32etbrFszjtMCl3yRZH51UMjJfuj8rXkW7Xx4q1TaHd0aox1jmKT7KW
j4Qm+rCd17FkcjhOA1W4NJUEnXcI9cfuT4SZIfq/VOpO1YLwZVSMuLrj+zOBex2ob1X1eHNF4gsr
Xqu1nolUJy9RBdszfo3wjyfE/2ob53CjjW5MylpGlipS4OScGlE6JbR4twyhcRzAWaStG0I7Jq6E
fOXH3F/ZwtJS4cJjdkzHqQs32oVCO9W6ahxXQn3SWEHzi91KYxO6bvqhfIT2ZvP4PsXIoM4ZdcOH
oSEplvkZu4Q950IXD3JDypOWb1TRqJKW/C1ABDA4lhug1x9961ZVc5RWL6MHDLUT6U89C9hXwRYb
r/dQqOixVm3vLk0MGNzWET50UqmXSlHhAshjaA38N1FI8AGI6h+iMGlDSS5CZu9pEhOEeQua9WLc
RvxCqDw0tqXkgyqtEhBvuKvy6IExvglGOu3m8zR8mLiXTk7xOS/cubtm6mhNdBodB0CLlxtsgNrm
X5bh0bBFm3G+yNCs1/DMfls2+XwuXkYm6rdlrIhbxk4Km+9Ie5/cvTyaBLx0T93Q1tOj3qrQCKnb
Oud4tXjj2odgrx+L5xBsGWHInzjwYq4H9wD/vah1rx26SHVDeevd5iuJwLsH2zycaRj/hY0uDW79
ApMFf1QutTNpZ0+vYWtrVIiBLbGs3bX9rIfVFmydmHTHI6j0t8SAER9lAkX15HPspqVExpCmkM7/
OREwD+dbsCA9lKoXzUgtJEvZghQsTPhbgNEweeUgCqoGNB5onBtK75RS6orRoCg+uHqUACsspjon
27VY5QJLgjp6At8lRLBjzdVAVfZjG1h5wr1iyNtnd1JUJrl4ye2H3CXWYLuwHM4yCJD7mBmsign/
WHngWTuuaiaWiZkZlQjN76TNOcEVzkthUbUvihMXYuC13HNHSu7+UiZA6UPcm3voaImCApY2VNxJ
ZfuN7J7owZrWFIuYwqCLI99iHswT0fyrhkOCvM+9nlTXEo+e/m8YamrAyHKsJAXMyTAxyBJaHpSQ
4eU3g9isGq1EPHcwwRxCyQSU+x5VAZM5MHQkgvXKH3xGLRAWfmTX3XDtyjcuhyMcLnkVO+DNZzaw
BiYagaBSHl98xQowqwsZB3wJ7t7Z73I5NFmHsZqluFRQmzBXrrKJJFj9BdOWSJGfUR3Fn08sU/LV
MMj3aXiwQ6M7k7cWLBQBdxfF3iEXKwShagWsBx2KaKNmEXFYwAxJELka/pD+4MlUBx1vbC+5zQI1
j+S75rv4Dew6GkjsIcvYtrCrN/A/WVl7A2WYPrR/y01Bo9JCQhAzcVjbru/yuPXAPGgw9U/RUe/5
j1PljXkRSryhi+NNeMefXzHhpZVwpzZidADe4BpfgQtr2UXdLlVR37OfSG3rQSch1CL41OedUP9h
KQ6/UESKNPPBQ46qO/wGOQEfVcqpn4mIGj8NSz/vuxr5MQhcuJhdGPRQSC8e6IZ4w6th89mB5qb8
jHgvqMhDUsE9NV0BJv4s2E3N6BnuAZLhImjARK955w/GfYmEPWN9WpJLSH5p9/Q6wkTZrOBqZVRO
HvBsxP7YnD7hh8EY4OXdEiPXGAW0EwdWq3usTbjoOHmAHHv4lBV9/uEYyzvMt/1vQtCz3B2OT0j3
4E68TD1U566Qk6M2isa9d/wx1+bfYpB6vaCK1OQR2BLEYBxi3pNPhNjt3rZLbA5WvPdUurwuLP5d
obvxatYlHuzzYwTomxopYJuVVx6LGIYX6DihjAseXWKwOdmQD+DTuLAwrqBRy+EsfsYp08Fm6uCB
kFqD3ezKIUACiYXnZzVwi4Q1DegoxKwnFl/50KcU1TgKk0jPvS6UF9M07Pcw3fT1k2WZRxKMgICc
Kpz0OKKBHt2WoZ50pWySYbDRfttrVXBoi5CLkRJj+6XV5VhOM6/gGxHJOnR+G/Q8sHZ7o3jAy77l
gx5f1nvZIu3ysl5/1XzPbPt5dh3+F0eRcNqmSOh2wcOfozNXMsz6YehvUH84cUcxXrStY2IcebAk
SdcOo8oJToO224YNTz3khh33JxxW5GKmN9OGttblNlFNQyuDTxo/IT5aylHf/TzRVyGstxN4KfuS
zz5IvY53AN7XPeryXy4cfpPnOA0n96Rsl1pb/1re7JbwHc7BkG+Fg1fRU1XewAWXJjKUqYE0j/o7
z7hCAZGV48SfXRLEHi0uvSWNpSlkFsNNNoh+RpQ+Ih3tq9FED6+F9JTZX7u7MsqoA5ZCV9W2GAOp
s+iQtjJvdwgvUS94hqfIPxwtGyAxSRdj+UEKM7KTIfCh7R286GOfnmWn2kHvZD3SLXk9PH3kRXBt
nrTfhvZ9vWhPt1P+0eDLsE1JfMdfTuUipgF5+q/g505IaLE2/T/kB7H51fhxau/DqM2VbecwEEo2
qXDivXcMUw3Fdn86eeL3g9t6tjFBLD2JLlj/HYEdFCtujeCIo/DUMtqtjHDK/SvgSGVGSeHA5QIt
WcHcBqOuf1Zombwyjr1r3/OhKA/BpoMqW3rS32cqGpYC047B/gakdaLv9JvzZOaYb5sdIcr2l9PF
mm6CYkeZnw+/AzeUNcu23TwpfwPYi4+JsayS3YDE6Z7flMP5PBeUuyNzrIn0SSpc3x8s7K2DYtfr
hCMrWJNRwoiO9tiJ1hNZdHGRgtERU5En8PlwHE5CAexgqFstsSbdr9VyXDEj0qULcvOfDyp4ZFIG
P8BKyn1IuNBNHNMX0IPMcBI+IDwHMzmO/p88NDTdQInIBysAS2qXDp3E/V+wJdo0tqxIyp8TiHDV
NU2PJx2FurOGa/077kIcgLWozS0id31PEjPVoUqap06WGV7JBnxymITOoW2mVM0FVxCpS6+nfKur
+VHwLhDmw9U/D/1uONqze2ZFX8uWgEyUmWEv5au+PVLX2iBDyrevJzqGZPreFvteW+ElG4RDxJL+
fEP/8C7vp3AX+6Nl9Eh89V6KzXc92xp+8s29d6a2ZEwsJnZhjoPdkj2t4FxYcAR9zONk290v7I4M
G/mdB5MXSXlsNYzuXFdcPTFkrJcxzUO0YrpDk6XbQxL69F/ALNVVE9LU942mD5GIMC7j+vPovcYy
AnVgHKKvW8D1bCScCtctHqVi1A8l6JcZ/G+oqAeqcLwrhgzFXVwo9k1EE0/LlUjPKgAydfT/lhIr
Q0BFRERXwI9u9pEG2Umk0PUEwBu7ZOCuUhVKiLi5xuWZ57IPM8CO38ogNtvGIQ3RL200g3UCQELX
Kb09TORakhf4fMI/X2VWFG8XQ4Bh653xwLB+NZejkcLlVjZmguapEhbu0JJ0VtX8c1UyXQsQ3sPX
vgorbQ27It3RtWg+7I/DPj+Q5oW1rvqyhWplDs9q7PIBgG9g6zxWDfNko1ugw4AbLrLAuKnFShj9
cU9f2ZHUQ75OT3KvAOq0CEqYzz3sr1pV0aF7lYUwtrbjaOIpE8H9aVU3xKuvMqEPOKSfPvwgmTff
9MIb2HGrRqKnFJ8vZW8yVPrhsfTjPW9Kro9PwaVGdw6xXcNViNI08O1IhUO2ykvvMtKLbYh/mCIe
Xktv1pf6+j43uyuDhprBYPf98A4zWu/YNXG8taykh8Vi7Y78hjP5uzkoHwVDryDxcW3Z0aSrd63T
Pa9d2H0qnNVrgquXWq7SHXDnZMOLMIROgr5YH1PQeXaFqmaS8errCfrCckYpL4wfkVuR0BRFqLu/
q3QzzAGicssQnl5mC1ceKrtcn+GFKFdniBzCqJCpX5NL9dc7XoLkFXgLzTNhcCRB+jRAPYPnnb4q
RYtOFGGz96/Kst/pOxPy6xUi/PwtLQLgSdH9slFdVOSKDQHJjfkHhYqckh9kQVlLTOHc1dZ8xS6A
tmYWA5b3ma6rEIz6RO7B7G/VIiOu+O6NBAy5bYDBbelFh0QldUvOVBw1dyIci8F6noryIDZcrUbz
iUw9TIBa2sD5ltzDB9AySQBYaoE+RQPojy8Tag9tGyS+oauWgV/wuDnfCRO6pPB19PUB3lcijkGt
JppYu6ecokN+XjrQJwmolt29MBBXOo8DKFhN692007C3FxSOaQtz7jLXrUrmC61RXKdtu3tY5fF1
3hICw0qd8ZFqOGi1YdyZ/GGnKT215iWQ6thwUMeBCP1uMpYKPDKxxjabaGygiBjFIswhtloJA9zD
aDPKvrOzP4AqthKwejXQi5Dq9NPORGyvwx58dK1IpR5bjp4ThqViTFiUcHt9G2CLpxLNBaId97He
lunBLkoMMzI9LAzUxX8oIeb6wIb5LthlDYClrGxrVNGZjxU4u3DihIQ7aX6v2skyY+Wi1lTn+R+s
mV+nvXEKCnr0AsubwRFAbchAZG6DHpRjPOvQMKMVxSl4IEbNGzgCQS8Njy79su3U65dHSqZuHZA1
BA3QkJ2Uv5tBT6kr4EKyHqcVpJS8BI/esPKPoB3x96V2B5Ofc15RirQWJPBT2iReUS/xHSwqF5u4
dz4regeE5dch7O/NH3mwlAeQhQ9ZsfMKx+RvbSwDnOtt6LzJ0vMCObickvOTf4trzrYm8O/8ATq0
LQ+oKI4rMQxFS6gj1fFwrnexGNHuYrT4MuurQLkS3LTnB6SoV+bWm7GDQNvsUXix8muZanxd0OiP
kVmzp+lFfVbr7VTE6nzxGMBDScUpRgSFqZAGdWVxAgKFttgT1UIjz2Sq/P6v8t5CAoyzfExfLrlV
b10ttw0LUUUa36zxTkHXjpsdDcvNAOBYlkTmvfuSXZ795q+HdJmZEHdF4rmA3vUrLrvvZiaFOyC9
qcE5idxL25tUxFIlKM72ekIdHZTq7gexZLZlxNByJ/5aRGkeQrz9XlPxfHhHhGbGncV/ideLXJim
qlAtTpbDJHwRss8REwGhddKY4n775ltoKFRjdaGZyq04NXXmk7hXj2jJkWkwqR7ThUUs8+m/0+N6
h3r/K8O6LzxViAI8wwTgU1T7c+TRK5JgQcgeWlU+cux/aTvK7CW28XBkVxY46aEmvHf0TlCMclTA
+r6HOp0nOxE2u0jcvNvkRai3dKfzqcbQArFKj1octi4XbWoiMZ75HZpQQ8/ZXxdXKVR5w6fUcVAN
cKwWNQaUFWqTP/QtNWqZ/bJJfWymydy2djE+LATm2kUrF5dmeD0l7SKnIfItjXrO1K/ybMVHCAQq
0ZjpU3w6Z3C79atiNaI3MdKEW3vMNw9H5Db5JB6Tf3SvG65GY6X6ek9xTWttxz4vi3ZbTqaN93DA
YScgVttMysyurWY+m9/Ssyy5FPZa7qgv3tl9uRyecx/CLngIfF2Jl6JXubDoJ3cVJKnEvc/ZAJRZ
FFe4BeeNVv1LjgEllS8jwwOMcqiwmzI+zdMyCAqkpUlivwKHTJ9dFueItSsh5X4j/biQqdqN4+aQ
WJZr2Sc7guWEw1C8Y8ZKmyLml3vXviijI3dklU1GuA/zpmiNTlJTHIxlt7Qd7qqC74JsVdcPOIrM
+Sc5HMU/yNXAHgbWhVts3E1P0X/73UhuAKQu46Ma3XGX9GgZfnFpvEz1SmTDRToTNbL05JFMHJWx
kO5TR4pllxKNAN22fymuUe0H8f4QLZBK3xEkQvNEPRyggeWJbl0B2y5UjAeIsQP5BE+dmdLtSbE+
9DiQdJWqy5JmM8O7WjtwHfwbVQzroRGeiRNQFmu0Bdm9knkTIL3mJauVPgh4KChm6rHiLYOQwXQx
Odxic1GlGzKrZHuqCG5C25x8oLI1ut/3yoaBpr+ilf39/w3uDe4ZOPKxJVu//OBqbsFj3qV3NaAn
EsWfTuwrPx5XPc6guM0o6hEbkIo/4vUpQvz6u2sPypCzg8bfnhEEOLEzjyiWRAJLqAD4wINWDoDb
wOhXIwnDAJKFTSKAAZw7+I2qpuxk0EjgKsC0tvGjXrUJP7cwUUdXvXyuVYCVUn31Cu+Lomdr6DAM
JYUE2WKdbxFPGYdSa25af4+SVNi7HT0dJkjiPa55kcPkfylHlrwx9eFLVDy9b26Nm/YhyaxeJtRN
buAz2soX3VEk8x6KX5qJAgGXliP+vFmADq12A3Ti6ZQHU1/Gs2VsTumyZ+rVAjmnpv1xD669amEq
EWZs8/X3luj2fhoBmT+H/QI+sWm1hc4LvgpjK1q8ZQMVdX2mxYJ3IqDqcRySf0JRqdLNZqEg9W1f
yRKLfjUUM5XHFyFBJyAH4Q4UMcF2yYycR/PJDnpLJTej2FSUHwn2TFzffWXdu+WA7YX1eEGiCBlO
PxbxWxbVisY50KZH8xQryvRo2KTX3T8OdmwdqRuFqm4lt5jeQMqK+2M5Chta1jt71319dzq1B+ys
9gkzLXNZMTBSNSLsYYt04kHhsCkhXMVTBv+YWZt3fw+AqvYLwLQ3BsWGVsDTYE6+ckEiCEetlcQu
cu6/NZywaxbFQeCasTq6LaHV82aCPFVHNtcRURV3zgzAfI1qXEeo/CY4lFJ7FFIXU0jeTQb+a542
ehASVArpEPskHwcaN/pb6n/1wEBy0SbECXiNBMB5a3laQ8i/AJRvBtWVVCXVTMlEuiiKpMY9JLWp
0dGNCfRMT8U7YvWPSfI4geF6YRfcYU8Gzpa5697NNocsPjEUxHEpGba0kpuZXa+MwxtbeUnQ/n+A
HdhPDDZVJYir9zWs/KMQbtuSHnkxiYRMwrumyOMkuGCrRlcEPAjDNHMImrasT7K4HZZuGHPW8spd
0kFMIQllct8lTAuZXkWGtjVQPJfEruFc0lduu2m0b4wRi0H+V3UQrMgVBVL3aq6xv1ChPFhAVm9j
l38F0SGxoIfehVZu+8jS+zmxDsiyULrF6cw93Ub/UgwOu7OESAMbcF+WxArmJkXVuLkO0mp0xRxi
PMvDMI031W2zPFXjT/rbrn/TWh9iEw4w454flIOe5NgH6ixhcX35SXieJT8/tDGexzM/ypjbiHvD
fJn9ZTqTbHWNDGfLw4N3MJgSWovDgIx0G3z3XpnndOYguR0pigXWokpliPiAJoAqyS3NlsU+TVjT
31hTPlbMZYZRWmvMD/L0OXGHjbXur4OROuB7qyOgnhhEG5ZQD0XH37rZq4CMXc+mqLR536leQuLf
2/GRRirFZbEzxUFkB6ul4idkP4btMb08TFi3AmX/fKTHhISBUM7QzmlpVIJ71E1/Kcc3IexehRRW
V4WbnizrIdjuzlsAadEacuA6OrNxr3zfRLNJxiXHfIgUHfLV2cMREMlL/KWQ1JBAPrsA9xlmR9nZ
C2SLr+GAgz/8Pv6Bst43AudbXGb/ST/8ziydIw7DH5HH95gf57k6tv4xg99KUohsxM8dD4s0Qm1z
Qo5Zq2jzfacVMQ8N7BW71tB6np4vXItVHPakm7j4oG7s/kK9/2JWBA/bJ53Co+Fw+OLnpiIBlROj
A3Fi8o/fxk573YePSgMiXFuF1NnYSRPi2vLIr7UBhwSX+SseLmIEL+YNcVj0ZyDg5M1R31u0PW3q
bkUgv43w63esc9dJMdj5TIA5ewj6izJU44LdZdSD5CWOJCV4mNVapPDwdp2bl78c0VdK/JKYDl4E
+b5A+IDAiCSOkB70cpvVqGz+cOBUue0bkuQjLMex2RVJ7c6N0QIJIFz4VB8bFPh7sjKPF7xkzNN2
aQ898fL/EVe78KzrQDS2winLAt/j7vLiKM7lle8XqdPN0MRYomZHQZfdn7GsAHTWc2uj4ylYcn4u
tqdxuYD84u8OZI2ZpNDG5sDU2MrUKLxG4qSTzmElwdYlabnJizL1ZH7LuT8D5Ghbao3VNJZw0iYh
z09NOD/cr92S5/g8W1Exl9bSJLizHL/xo+lpBSQjo2EH/Q5WpH/nATetmtSG7/sH9Sws2cZQvSS/
ap0vO2CMPLc4MLd1wQamZxlDPDyFvchnJeEnKj7jiTQ0GAyCKXq0tA0h+1PW43iYtkpthuQsBHoN
kyYOSuGPSuRaYK13IbX2L/jMO7Mw8vWAjiE1N3/ZeUod9rl6pbdUhdC5f+CxQElMa1EOT5KL6/jf
atZ7Ch0BFNM2VeG0C+e0fRsHvjclkWjJd0w9uHbK7SaZBxmBe5z0bc7nEFfT3f/+gUyVZnxOgtQg
1EI8ZT4Y1Wea4ks/8KjCUrAo9MivbMHcWBuyk1lC0GtxXYesk6LwqeuzNnmIeLkbSs/2CiZBbjX8
G8OnJjyD8vqaCwlvT8As7q/Orr5veOdSAdH2kGf5RKGgVe+mXuLD6uQYzPUCRZOM7F87eS4jvpHa
PEaDjegHoRo2IIHQjJ1wT7PsDn9Xv9V34Zmi/KZ3vQj1rl4Ixg4VIMoF2JZhZhwWh6D2ZS3nhIIe
++Es2W1oUszQNsWVsEF6WVEt4JBPmO7TJExM5hvWN+nEdLZGSpdhp87fDZuIwLzAKd77AJi8fwil
axBarqmgOpeeIOgMxEQ2QWYkLza2+n+RImb3N2yNkcUUBOA8kkPLe5OQN+Dm49FQGIcZjJm+ggZL
jCn/7HzTIXJ/SsPzDRsqDgjVQN+HOfTZ542s9VjqSnBt4VmiMMdfO6vvjVE1ujXe8/ygngR2eUWE
WijabdUHuTjsWLsK3oEqrxepvkOLLbXxZMsCeGwvPdDrvLqQdzVGzj5PT1nYnVS9tXJb2MoI1sfe
oH020JVJFQ3LpbO2yEcb/TFWi7XJbI0jD/T0c5R4Up709Fd3wXRYPrwEjGbWCRbuTBl46BhGvTp9
qbPZidnuVJaWC2wfhvEDE4GqhGFpgnNBNNAXEOyHzqxJop6G4NhmbJcWNQGmb1xVpA7sjrz7HmmV
zcBXxnGOPx98C7KqKeuiKcC8ZYndOh1Lr78IO9PyrfgqRpjC1EIl6nf2iLVA5JhiVwgajCz4AcB8
pUkPvZ8C71ZJtfaSreL6kLjlcLt/43LPI72H1VwGnUDoAayHpNt1EanLyEr/OoHj+jskaJsSOaVY
VuFAT+TIXNkCZd29Eu51ko0YBBuG3K/jxdvTiGKsuj1e4pEUu3b24unNpNYOEkTBvNGt2HLEo3fe
h+2N5R1zX3RVgoabiK77irOGa92Ne8r/YLcyUTzfLI52N8C48Ftc8iHMUT5QlrHdRCzU5CFwk4jk
SccnZzypxy/lDzSoWry2ZYqaAO3TB8Y2I0msIxc1TRKahuQ1b3NNzs8pzqxsTxz5nnpEgnkFS1Lt
j8deTFzMdtTbt0rY7hTe/gupLbFQoOiDU1/og5d+yK1xbGCjusKGBHBao/+mpYQ5a1To5/kNDTeG
0BZS6ohoxPv5MkPaV1K287Q6N92wviUti5ea4KDw01mRIt9zFZsQSN9986Vd/ut3E0+vaLfUwjZU
ybZTQofInizgn525mxUFmWZHi3hQDL3S8qJjdspI0HUDZuph+PCMaqo+TuuBJH6SCk9OLCuIW4b/
IfyD8APAJnmSDyVUb/ii32tYswmBl56ZZpg8vBAtD6QiDsKUGWHnV8FJ8AJE71vslYghZ7dTYU6s
MRb1DgiKnNVB5UtmYDh8HDqTVmYBExRnEW+wddbUAO+n8J+rsJR+KtTdDsK/on17WCACv/Fvnk4A
eWnlYf+OoQf93woOb0jh7SE1hE6K0JLi1lkQvz87dvKc9TTHKiRHOIhMwexc+ndy1567t3vkTmcy
SmeK3STrOcGqbIEq/hc+dt/gvoRQpevJeUaAWJB8WztKMwpqbf0zv5g4IsrRbgOIVG7QgpAksw8q
Yuv9jpSToR9xN+DL8kladnoR++sPZPiY7oH9dhSRltV8BSV9blZZrHaEsyidfv92qSSweM7Ie5Bi
0MIOgut+ZZtWC3EnqTt36mdkwrYqQbs0MQRsr2nJBFOPbBamdxZHXnnctN/6Au/aFziiLHK6PLnN
WZ71u5Wteahp8E4wO2XAfon/4qAqi4K4lFJ+sBm4BesVQJbEYVhcbIdzMWKcrct6H0qYJ19D6uDG
Ww+Wdpq215SpN3ufCTo8FxoWM44NXTr68w+YQ7WJj4+xNM3sOdTymu1KvXDQXCSJHz7P90DAyN6y
NJfF26H3dz4v3XvlcRy5FzMDVfm7x3qVscIIuP1mWxmLrj6b+pBHyaFsQjl4/vqf2j+IfupdSMU5
jR6R3j+pIUvc0g+OzrWwehg6+7mFoJp9egTvfYbTE66RjgOnOpuS238fVkGbGNhKnBGJqxDf4wPa
6g8H2M/z8icYhGUHU8yuyZvZdFV9W2PUORgkggMxx27NXbrhdm3eUAawmL/vduVaDfBkJDOZtoQ8
rd8I5BUkaR+/P52cFLu6e2qQ8uJ7HsS123xjKF8PacxKVpTMSvrPazXYAlPYC//4jH9CghtsMyIu
YMJdAFE+Oxj+lIt5QWHeSa8MG+s62N5otX2XtMLvYRa12mRl9tihi9dO3/OghDXdLdeWdGkNK+t3
yZ8BwuqB2/8dNWPVPWQ8kYw8+ZxxKr2K9AVtXpTZl/jZpDLoln1DJZlA6DrKk3Si4pCFlHwK+kca
R5Kva++PyQ/TCYzUihphJcNo6HV/710kOmB7hcZeeYR09uknIoAgIMZsPsrIbtR++X/beR2GFCua
8K4Ao835dXwA5CZpdUB3MdP8aa3mgQ4XRYwTQJait9mbyqTWTRoBVAP4ivxh+pwqMrowqXhzSEXB
c/82wNHdwlBh04ijYiN7qpQ/OjH6NDFrtbqHMV2cgTpTUvhqwo+jtVZ3z4H3MaX1rf6NeSCHtCAh
BLn8biS1NJaI69T729//9rm1AH4va7coFnOa2jYqM5yOsCKhsS9f4QrX65830uDG8P2U6r6jUcRl
NHQaDXQWHNKI94LU1hz5H/QeZkkfZLlkUX97u2/k389LrQx3e6uEntqVsw9BAXoFwiW4OxjH9UGx
QgRbo2AHShfeemzGNpyIjt2rPlQIQ5G6Nzb4CsHdwG+PMtkUHNVR7KdPeoEdWZp+LkFMwXnlbIyY
XV7uvnPZwZTn3mi4xnkTJB5/hLajmsxQ9FnY5YV4o+f5ChXwLOxnqTW9F0gYyBcADBMDUACuTUs0
Myt1VIwszmZjMHzl23bx8w8kz+lqyiUMFdzDrW0R4McmFUspgIYyLkYBaJIRmmFGwFB07z5X5Dj3
KejRdSbosYFoWlexFTFymRqMjt3mVu3sQkDE71/r3Uj6xP0vCtUbNJvFJyBgbdNod/trSTpcJ0ZJ
REFOXR1XfOI3O20CMl2QvK/1gxE2y/O05yKNUiJeZdkYqaT1vUSbEgS3RjtqeCuP0ej44G8vSBKa
hee4JRtBmrlF6jlmIzbK+VvWoYqw8w+5zPi72J9d0nmMrVEs2pUnjogOSqoDkyFnINphRFW+Gmf8
BdMZryzvVrdWA+ewsk11N7BUozewTWgCzNSS9jf+1fLrmo13yXaYg3aStwMC+RVTiMgaoxaC4ta8
E+0eK4HiG1bP2Bl3ionDnfe+lxbr7owwmvsSSXEavMAHw9g0KucPn6ms1941Yj++WYB/NYav2eP0
y4AdxaqZ9Ccw+IfyJX1zBecxvke//uaaqK73ejQFDZMec0+t/WXqvtnX5H4f16xP9uYdLkrt/lcP
Dm+GJfL0j7VUtkh0jug356avtLia9zBq+iWjLC3FHYHMEpZ1rWnIhiDODbloxvg0B4B3D6KSx7P5
P5NXhGbX0jCYT7D/SLDfdjLDTjwIC53lBjFPKN5GHrROZenxTjQ/gdopezpC4HoA146GvgLe/VwG
YF+WXdcbO2EJcJBMahWtuKLx9fIPiUn6t7AuG7LNzoLldXwIWVD+fV3t3mgi9fqeRD0T9Xvtpwe6
4yyV01iPEaQLJq84SZPI6MoeTXdJKIxmYBz/V5IS72xUOfUyG+0bk2lBbH3psa4eNFyx8jHNFK2+
bd1z5fHwihspZh4w1+Vt3i+fAGU8XP3Q07e+YPK/lfgMXhHoeBd4oOcLEhLF6AcnjmaB/GKuqoan
VZionz75q0C+oWJD1KgoTQgb8jC6n8+U4Zs5hnb0qAju9ahQiHnFC9Df3/iDz54PWrA7mFfZBrAN
UhuuioNOvhUr8XkIO1ieI2saFugyk5K1tREfSoGhPOziVJa01moe40+K5byT7eU5NIF/TeYJqh0Y
ZY7vwFh4k2+aYaX2ADW5RrewIbeN4QK8IvpuXGzS5ekduztRgmcmF55qFOuUHtqM6Zpd1gPs9E8p
u4afqmDnkOrWb8oROukfMWyjcvincrpY4Yw0Ry1fNudf2LsAZRtiPwXtzlk4C5s6eJ4W3Gu6TGqt
YJGPGnnRe8wHZehUiCGNWgW+4GFMAE+LhG8DrqQTEqOlRAzWdwTtBiQQAjv/DXa4+cgtD686WIh6
lvNT2U4WR/sBygOm+AioN3fzkgIps3tnzzaz8Ns4O5mRXXSNsYJFalSJekI4y1T9PkG8XgQvjMgU
xvUYSZFioJI0ohoghtiqdEAN+dNnF78CixKVYAHVDsild7HrVUiQgpOSvXbVywG0wSW8t6svAtqG
ssGy64b903VDN/l8imUpQk8keRRZWPSxQaKgnDgjLl4Ccw6RZsyBzhAU3uJItnjI6YLD/klfW2P/
KAuVcFkt+AKDFH4IAeUgOq8uIjkQllfG8ELWCCae4kaV4kOD92JNBKdhjWkc+dzcnplHPH2VRIi2
UruhmYXwBTlfXQnSYUuxpEawfohAhGi4RgcCRcSfZpds3Ziq/5XvSxMp9F0SRobfmGJeSEoykyAx
Hq6CSMn7IU53CHwhF2C18zW3+CfVguoJDsbbnq4OhdnNOtt2MQywVf4LD3pRuqGpVVbbhxmohD1W
n+gzmgri9dJrEsBXccbPGujl9EosKmjK1v7L0kS02IGQ2/CufBxm6p4bjr7Vka1nXHgZdWj6AMVb
yX+SXjaphVhPcfNac9/C92aFouH2hrGPozLAx70EXrqVuyYoT34r/SOgruy69uCGHHrBSAU8wvLk
jP/YyB/VXn1/jSVyVmkbjQPGWeGGdCwSofNxSi1AJjfC506aeV3wkTDSeHiibzZZ0kFz6+jWCU9/
vbK/ewje+9/lpELxIZlDxMqnH0ftqBnKmZcU+gVTJBS1Cd4eyzp7DZj8yZdr/5u+sMzkU89t03SU
phOSpDNR0Il5p/9NAyJndvEvurzbNN8mvyTYmRzTOUcdRuicAW3lt5KTHp8cfQqM2/hM2zp3fNZo
kWWcYQ4arMr3+UfoAxg/tKy9Z0XtKq3klkLH/jvFWT4bmB0p3e/CKRmY4KhgGei8CjHc1mbAh5gS
Ppemdxo/f5IwwKEcEc5gaE+fSe4W1ZgM1Snrmsult72s8ovRPnxSiEraCYGX4S8C7sjRBBHZbQyx
akcV9FmXaRukZu0CiEB3zFHJp42nYc1AKNBAGZFHXgFw6LqLmujqiYb/PKvfu56bqJBVH0/zPYD6
v8ogAhBpvigqjK2Asm1DmO4PuclM1gixf6xT8QWfboyge7o2RMw7FenKeVViU9SsMRscIfw8RqLY
+6WmI16g8iqHAAghG4jODMpdlGtppCtNEfBe3+BnBXe7Js4pDama8cNtq4pIMwK2UBXLJMafKHYs
D/ZUDPl2S8JeHAWgRPkVY/J+wY9Ovz6HUvCRGvG3xzHv5Fb59StmhvTvimyniOQy3Aj9UalNbvN9
ZU/RHqWvoXvwpO7MvaPKufp/EgRMxz8LvkRNpSWVFW0resl9mzxigbbQGVULZlWUff4mh4XoGrcJ
SAYBFgBM9Kna/FoFCmdjw86VM/75GGq+b50ZTNsXNCkD4IY1X20IfTPYQ12+qV7sd9l26m73MxbY
oNEl4LoIWzgCz7eXFUvEhpkyRx5PWfxUt5NHV2emiiR7DbvYiTS277vtWylws8w1uuL9u38SeFQy
oJoKHhSK17d3B+SRr9oZ/wRHnOB05fiCHKZY1aGqUOGCJMqN0mJKnW43p0djoNOn9Bbz2J6jb3YS
TKxHUjOUuX+OHsI1OQp54WRX7G2pQvL2SWPG6sKGAdDIk0iDehahSmyg5WRegjQLNYqPYA9vipVq
czGgC0WO6PtxJKDBcGXomi5N3+QBQKoVIPK1rilfqmTKeg4kYrduwVSZfdeavrw9Ooqzjh60fbBg
1NACuj1/bdwOa+8NvIBT7mlQ1lo1H9ytdIO/i5yV6Z5l3NYYwtcxvROfnen3RtceRup/HpMPpOUL
6jHVQMNMJXZrNpYBUAmi3honwldz15Sx1TPWglYDWpfk1cQtwcbiXc7MYf7dU7Pfx+kEmtsbQ/1v
KV/rgnC5wxVUf/Wd/nhqoF8o8pAIQXHGZIn6PW1mD2oz5wOWSCJCz+bnWO5ifxljsW3N8K61JdBF
XHkfQBaBWhbl/U+tmHymvSndWvAZApq+q3agGiQQCgmVe1UoiBttFt893qvY0nNbiG3u4PLmUEVk
a3d+cU+Pn9/0ZXcdbhL8GnfCCrvA5lAFG8RBMIjLhkcvHUbmSytwas1IlItSp63K3OaZhvH413TR
YbUKqzRyg88oVhgqS0nXQGILStN0+xAIggkp064IWX/+wIx/Fw7C+dcoq4sa4BuyHlyLF3I9ggOU
Iu34aciYOhHjI4vkWAhrUjN4khq67ldxlJxpZOTjTHtVc9PH7cq9GayP3/8mpnU3HyMLiM11jfSc
ksyOSj4xyTJbIzPMOIV/O+t2D83faDzhGAxszq/4j8VPJVarpz+2SF+d3p4aZrcBkozZADkKSklL
b9OVxEI02z92TvkvK2nxP8C+4ezspTi9JW3SZKDoJlQ7nKOqmieFwoYFaBcjlpGpBU56yJadcKBa
o7RISl4EyIZjDooixi+jw6kmghQNFwczUPDHh6eAGFA65ABtUnBEP0xwyNIIBfFOkLXQuX2Q4NtP
h5WcQW5Kiw9VbcLc1fQFNVd9+RUPyIiFbFK8J7Al3Uphk1a8ySy6YDHBOPHBfZqZcnpTHevAtjAl
XvnZ028UUWIOkXEZvwXrKr7XRdS0BX0LXKuTKmhgpSDKn8orCbZN57v+H36FN8PXaMu/1BOqRxvo
Dhjnkx8OLVWPe1HzcgtxJ6FKxea3nlkGRHTL+U3/E/wieKaH3HoTewZmbGoSmLCnSYSsPEPlCcsm
HbjAClLOTB9M5gkZ3WvkfyGoiVRstClmLlvwmEV+QiuqHI/9IgxN823tHgrUOcB2GINZJwFz4pSJ
rw9py4WkAayesxPQuKWm8N2xdDHKeajHBccyqzM2zw1uvSByoYCAdJpWWv9/kilMnsxkt2HyU9rA
ihhbL+hE9Laya/IDoplcL+rqJYHEo0onLyYS8K/Wp4/i07KGEvkQY3h+igu3THnTHAjGh66MvaPo
v4wmZmIWIdPrPbfcYj39yuSnHzn+J7mJo+PHjTs4JB3GZS2nNd9x+SyM16wun2Z8S0QIdIkJ4tSh
E+Pr3/6wLrWaGs2VGY3ps8H9v2N3c1aHoL5cEe02IfIzX147kT87NvxDIQV2ZOPf5wb2znbyoiWW
NeLW4GQiXpiBkw+pFeRzRT3gaHmb12H5rxUpcXM2NsWP17bQL5Q3MMOMARKGw1jw31mZo1Uq2J95
zP/K2qpdZh/Yhhd1Ldok5V60Ew7IN9OYspFYX7nnrqYuknxeAk057Yv51zkuGuJdx0GCwEaJu0NU
13DYSwLpOs4BmDHgjkHcmvdAL2Ap9BFu0YvgntavNySgR6sVj4lCNtGPJF4kBWKz3IF/RSG8xsyz
Ux8kE7fFqfI2uwiG9AB7+a5KnH7f9AtU28UoIwBcCDPoldjfCDn+kLYvdirbpm38alQQb6p9Phr/
qosFz56IPuAQ7BI+NsGBi1KVVTWBoxLwTarNX8GBQ69LRbQwnO2vdyLVtK1iBFzeZjPHwt8AfEfv
iHDbDlK7cvaVFWCb7V5hAN9ePNJqbdPMVkBX9JFPS0sopw2NUqpzr1rTb+mJ4dWUJFp6P73VXlVz
94SHlCokH+Dz3x5n73mSHNzxZjSMHLlxVW5p78kzUlYQ4zQN0VvZhmJZStLXhfnsyj9kzB2oSTRU
LQQAzUdvyTCPJ5Up+IZIJM7AoW2SQKooJdSuoxdRDuL/6qvUbVQQbYQqbmgBuuommZVrKJ3IQA1a
SsXjhM0aX9yHLRXky2JGYY3zfr7nhTb1cEbx/Rs2QlL6z2w2HbORVBUESVtoQmhgJe7kogB9fKpk
fQYBclsFJlsUH716KbQcuWlEj97EMs43wvPc8VofZKsGHl0J6cxgms6/0o5+enZKvH1uSiCluIPJ
VaP7F6vH9nVA2r8uPVSwyjJo95jbaZ0+hL03e6QRzcA8bqdB3gS+vpUTOMenwgUHYR8/cQ9MU/Jf
W87SRhPUN7pPL+rXU6yvCp2qfMrZh78sNW9rhcraQL9UBmCLZp/yASaNx+gbRfodTGrpaQliEgSg
9LPFEquVA/alrOEdj2FqP5gbveRiMaTpxrwkfe9MMsro9irBJ+DcwxcLA3SwNYPFPiIarNmCBwA9
8JjOc5wQSGJ5LohAde8q3PB3lhaoYxW+rtQc3Zn1gk0Wxn2XnvxYU36iTYjV98kTFlGHTB2w5dvm
h5jkKGBNVskqi9wiYhvsrZk9tHgQaRq3cN1QnD26PzyVuLRLsmz94NraeGc+0k4WoVs3cj+dxSww
v0SedYY06+MnpA3lRr+qy+DJH3PhbymXBPPFBkILS2yOqWYS6KByYZ6asU4y3kybC1UpqxOkOPZq
oNwBTKTRrozxbGPPcdePeHiMbenJfanu0pFLVDw4c7PCdoxn/x2BVE9bjw5xz2a85UsEeKUnnBhA
CfzI0l6ZH+RORhk09vyoTS5k6T5z1TdcZcHxhW8mEu9s08hSQ++FaIClwDSRpa/R4Zch4sWn6lQr
ojCYJjs6o7xYix14jBzqBwZYqilY4IVcfbSf9D152GYn+GbUwKnTMLSx7+koC2kZbdwwVR+/Cxws
Lo4YYh/NqQwgaeyMMIDDOEx2Yqd+k/OBpLhcjx3+4IC7nOAmo7Oxodh1oVezRoMbhKG+5QtR2ZvY
8BwP1U0HvZdQugfEo2Znl2mxKKsOAUzG5SykKrMPrnPc9KLqH54xk+sp4A5ACuzTi/krdPlNCPs2
2dCp1JB4cRFZPAU3ilnFpimyWqT8YsnUkV7KvG/4Q2XHmw7A/rvaSdNNH0PknlFLxVhFYjW1hdlG
Q+61KaZywBS30ujLCN6plulQ/TIwv3VafoTVQODwKIPQd1Q0C+875rdhwQkxpa++LHwHZfB1lEDj
wR2Aq/6dPnVtIejypFOp5HHs1z6nqJX+5JUmj8KXzchE/qMUERFMIJ13mGCgfkLTFTP/vPNGi7A6
Qee8xgvA9144nUdyDMCwp+d/pd9JWyrEaKBMGrihVHDHiSWm1kkpEBRyUGmbOZ3kKaTcIbYZvwP7
MmUX9ssIO3YCSr/+qPtyTciyHts67vivcdpbFbTzCbQ7y/UjjgxUvHrVk2BpPAoEbxD4QgbSYatD
7Ww5T9yPNvTiGbEIEWnFlyNj+gSWah6g+KOv/5Be1hr8OIA418cJf8emWO0eoBeA7cv05iKxoLpo
pQPZImLlaMabxT3U5a9b2woY99rJcembc2eGLZLouOTKsMQc/7YTuh96bwQ3xYwq9vtlCmAMD4ly
AxkyzHzZNwruEpuBIpN0xGztVutsnTZPNfLJK8W36Z4wjZ51X/IucHFotj3Bzig1Ei5ruW6aovi7
71PyXSikODTckbTayxyUz5PJ5MCUTs6bDx91fQ5WhxyMaT+f7mRmm+Z2pjaUBGhUCuKQiz15L848
GxpQb6M4mieOmDTHjOycZpmqaYKtjo/QWMAu0Iu/pyYQKMt5HFnW5gjFL/u9SXtCxmwBEJSSVSxl
Sf23O0Cg345iWAG1zBouyFb4XoJ1JP1BCXmrz+vIOKx4HuHRm95ywASR9OMk7gsjcgC9BJuaiaiU
KToao1LIO6H7jlqq3NWqtBIR+YB4ttkJiJ3bVZwQxnVhmlxEy8BptBBs46u1I6lB0DVb9lphIHTl
eyFW4PUEe1YFjhmzluN72SwIMnQiZlI3i1ZEvU3zw5WhD4JifrKZiV2yRshPrMbJ1widMc50CWOq
JFzFxleZbdbv2mFoeOVJGxDLz+LEQGepzEopMvG4yIuaUrrntZ3r7VkQBi/sQnBPp+jhJZlJRCNI
JiUq/t4L5Z2mFglI17/6vDVQbTrpMzKyR8srsF4l04s4ymK3tOH2Az9VC1dKAUEGubnigFBg7fog
NeyzwyrebqlLCWRP66croMaPJ4BqiLorXp1qjC9gW8IzM7VlUnnhOfy/3IQxXYvFhh1fuXUXRipu
Erxu73/rfP8y8oaEXxCtudKE8Z47lycK2BvdqcBPI8ISRDr2INWT/5bQzyium/mSC5LROKcgcNl0
nsMBI0TKebHRAtDZ4qS48ifkvVehGzsr+g3UciK/nDLDAKmbifirzNphy7GHbfzEgTJvwDmJFrI+
suoL7vhJZ4Y2m9heeCdiJKkHhJyLjVc3e2GDTfdmYspMZnh66BDeAg0xuPRqqv20nlZqTDZdWrMC
N0TGn+knBOYkykikus0lx1WpANAVeuejQZYmYm4XzytrOnG7zlgbw5BJHWg3h3nIyNlR1YxkWXQt
KEVEZP06JauCV/GS/HxZsJb+VGNdawf7+G07bSD5/eW43/vAnzaQNhiwZRnbm0SPeqliIOULfBTR
7h8R4WeT76J7O1xX4ZC1rSNg0aKRfkVqQdGxRIp+RlD9gplAK1AozF07LaKnwG0tAhaptyx0NnNI
PvKj7GDEuj1KxlfQRcEo100RfmKXtHzney9nMifAJt06bImpLfjnor7NOaQPMjKColwA82RgeGUx
5tCBoy9cXYvq3DlM0BdBcyQO2uYfamBIHXCt/DtMY5Gc/V4hoQjq5pekauzRz/zfC942MSPNMSX5
HP8GUtXrpZM2vW5st1F/DqEFRWTYoeKYYUToBl3UJfVFLXZQCLNHwLX6otroMgdc2OkXvpq+F9De
tlsIiUrfClB3B7rIwD3DDNiDizVAXtIMxS8rKYO7ZAms/qM510lMfBTeXaBl3UI1fRfFWqK4T93D
WWLJt5IrxvB+GKs7YAkObrocoxQ+QlgqUlpMszeKax7RCzHVjFknqpPQ/axyW06A9oU3YwLFrVXj
APpf6jrM7C39GyXZUUnkriDQs1ZgFFzYp9hzauCjYT4Ge25Tja2nhslOXBHBrJADvXzsnbzpVy4j
BNMnc6qxMup5XWO9Z1sPlryqCJ45t7vtJzfDsUsMSoFeruydctZ4mTqzPsXvIvpQk3bdD4GbLbdg
OLPEA9XVkB1Z9DfA2hlopdH8aJeRYOTIUwqC+nBlnBDGfE717L6/vda1FUd4+t5tbw4kALvg2dNn
xJaMb2lrac9nTiBGAbyvFRNz69kHpBk7bVRZQSVNoEq/3UyYs8SxHf30STbsfO2KfOCmnSrYDLyg
/zwXlpVdYBbkg7ZIJit1EmlUsieG1nCg94eEAGhekTHvj5iIJuUJZxu+PFfrov7xtIBDWzdmooKJ
+6Rivi4kFNbB/efzb+G3I+242KQeNpmu7hojhunCB3yV5KvZfyz2zXTSWQgWWqGO9Kp85ICJPo2B
G7X0V54NIMUccWVcXoxAAf6EM6RjNSKiT+VA58GPNz2jl3MlLS9Tg7k8cKpcXrffvysfqwVG0My3
OE/bn2mq4Yk/UwaDe2oDwCxglhOlC3L02wHc95Zkn4dFQlO1ETzjLcXgK5xAsqgLY600dwQ27h4I
tqPupjpM09tvdkkA9FBDqFu7q5h2ZOAgKrQsnPxX822Aa9Z0dDYVHMVdOhkltGl/93MzkGU7YbYN
PfzrydWOLGk03F0ORscxB41ufJe9pO7+nF89E4F4/GzUQ9XefvP2E1sFNdfBzJ++USEwTUVwK80w
vrt76/Ul0TCszTPVQy5gilCxT3Fgh6Z5SR8j7lB2ZqZOGGILuYLEGAVb8QkHpGxQUvh8OFOmSK3I
phix0gwPqPbBhd2B+lWdPSto9eRI8OI8xlqJMr3tNEyVFZSUxacGKRPy/NnhY4HY9IEDMJ+1xrfH
/JTaqDFP1v1hPHrvyZnS3l03gNh16jmMcXRp3brH47wndpwKkyjWrDxX0UAxA7u6JtvBk5N7FN5I
VYnG40u7rTVO0+dlBwSEhvDXMIjmVHJAUElZfpuRYxhqlI3iX+K95mLY5yE8cDUbjNc1wJfbeT3v
JMVbCbDv05mOZYc0y5Gv8m+b0sUCdTOB6c0IidwKxrZMOdzGIkuXH9y0pOZpk01pfvwIhUh2zdnr
qYI/tqFitahgc7rSA2io/Yp6Oes6YlXOVgkU5ON0Xdpo70W8Yy8vmHQe3HYif/CS7WuJEws9Vj+g
DKiZiVHzYC3wZ6uPVihVAH/VIKVznDOQoAQHj2UksAp5j7LgvQCmBTYXsfH1sVBzMBOnG4qdp5H3
q+uq9/RoFsPDf+ywRs6ykfJ9foBZKSwhNRTQjqdNPdvtcI4EBXr5v0XhMz0Ld/mA9zUKMROy1i1w
sly5z0d0X7FrDQX2K/6GNcAQBtUJgydA7Dk/XmUOdt9gDZwLZ+9bkss8RV1GbftpyBF1zENpans8
wbDvLJpzc0m8prCKds69jR+AtyJRhr1eHoZrtRKPVtfItRRmRByu4WadpAYNoGVYqNp1/vz1wV7h
Ml3PCEUC0D5d6egD0HrOLYYl+iV/RbrV/p8DOIJ8iSHiJZITwXmYW2h/O+NhwXMPLpoHnczvusoL
hpamg705ibpw4ypfliZnG3o7ZEtzJqipFtfEcfXZS56e69d/aOHOgOWuRYbxJls+Um4BoQeP8OIG
E7+6VC4xqa8k/b0yjJOyz7qrijnAKSHkFnel3kvxegFD6oFJn9plrEj8APnaGJ8NiCH5hvFtf8p7
IyDDQBgiVAoHw6d+7xF16UC/vStdJq1jGPIEAHVT5CjQomooN7dglIoIUeZ7gZlCAIeAFU7CwK93
oDcLbue4GouVwEbDVQE6hT3y+8Mw6gdfF8yEEBNyA5lKZ6h6nGd8sXCN1LWe2LDrMbdyvnZnue8a
2IRSUPcWgmCO9NJ92ryL9F4r7TXlQWGerbtg80wCas82jjYhWTA99XqbibSIbDBd8fKeWl87lNMn
d4h/rvPan4AgSd3mTv7NoZ3wjBpFDo9sbXPgo6Ju5kxY040PyFU5XP5l44W8w/gttNlegKbkTY0R
vTcGn7dueGldcadmN4di78+/LtNxdjd8PgLTkRn8yhZe2cV8EmypS2VCpQ9MjPL7sWDEL/Ys+0H3
VFtemkbqtZMZRb3X3jMFfcfFPAUaUtHwk+hIulgSOIJz9ODZXH7ov+PNCJqaTdKCaiS0E1SG7HFi
3VnybI29Yy8lR5veP1gEBm3K4d9dR4ATu2N8uCLQqNZDdb08/NsjOoN+XAqAjix10m15NW2YfeTQ
1Sv+eR0Bw3t+ZaIxnofqMF/sJRjRrfUyXSLUYEzFny5pTQYcPi4ZsvFke/aIbtkoOdpK5yZv6app
sIB+KN72ROvDJl7zETKDB5dBJKjBbLorFLbcgsn4sr2ppHKzUiYG9ZYMZg8wZvwIls0afhdk5Eel
+OOBRTMcLYHmLQu1cd3ufOSZnWIYKL8tUOAD5jhv2urFlaDziXRyInsTIG5LFCiIHAyBJn0314Q/
jM/eUMu/967TfzuxCEeA8zZk1AXIFiYnuQ872W9HORTa/6nBGzM8xQ/6X4LoKptBIvN5G0awWrll
N8yalrpz4x8DwrkSL46n20YxJQVgOY7UVLdF+OHbdEhdRv8dej5m/d2jdq6B0ILa3tLfAWKlRYH5
DaFxUbXhpDWE5q7FdZzeEceKVzoLUx9mEziuEZZP2pGUBhPT3TkSjtx8Uk3H1f2+C6c+2GaJW7R5
B8bek0S771OBSoxzHgyOUSiJEiNWslLHK92Ua5FuHd6e6yRN7i1d4b21dTHh/FIiCWzCArD3DYC7
fkU6Cr2ThDfYvwBEKvSoaG0l/cS5J9k7cprz0b3ixuVUe5UpfhEIbNBKLrzymKyiIpCj3myE28Kp
r2WhDh6MrZMGCP8eiR1NhGRMVz8vNstwAmQCLkOTInZAe01ez+NbTgffFjlaE8/6mvrjUEgrbq6u
29wT1mpAMOyhDudJjlkhQ9PKAX8dsnjwfJAQTErdgZ8WL5yKRAcPNTIEo0dT3LSoszh++RWuf5ow
L4kUZv+EKaZSoHFsCPpv+cDAMg4shpWqIHJq7HqTdz0hYawF7EDewiBZLhimEix+Wq54FVnsyKOf
jSTGaAPSeSjWzTFmJFOX/rCDmIXNBQcPwIHQLaUHl0at5b87IEAAOBitj9urz0+Aq6/YyO6JJDEp
u67SPSZ0lhB+Yb9D9MeQsl4WYh7tGG1fhRutIr50fW+S+xxtDcFjNLaiLXXRZycJva+bACI7MCLK
YvGnypMpIDl32RvyAR3S66JpjSeRkNp3revB5Qjoqzv4KJ7dGrBXLFgvIQ2PsIuFagk36m9qsXhM
jEbMAbH5HArjfeDQmp3rD6uF2p8Gak6aWRInKdfyp3Q94U07opmMCwS2cIGr3N+3C8vX8mOeuEj7
88H7Dezuh/WZIFJPfTNDJAE/7BLnd5utv0HJCEPm5wE+TAIAmLf+H+XxDhwq8VRvPXZruMEfhLxG
SClyqETeippCVBHGyT0S6J6I9opHXF0o7CL5ADxxUaBVTS+Kt2Hq203sea13KTwEhsTi0X65hRCw
kf+Q1f5HcLpsqVnEZicmzmZrIdB+wRbFmPnLAj/Bl0DGhjzUCSl7jmSLGyuQn6aVvBrIrefZwDge
k0hExKh6RJ3xUTfWJSXAeYn+vpfddnJVqo4NHDbgSEog+szQxZ08Y4FJ5jsEdaf4+GfP/7/rE7NK
qzLLNSDMBigziie54SGVR4aaWEwoMLAeucIf1dRhnfyM+tmnf9YLP9esDpQRPtfe265B+GAgqOvb
SIuFPtGfz3sd75fN04E1IWofd23iA4Ilc2E3gwZsZwZFsOnGgS7qqctS8qJYXf5fqSVPsD4xvEcY
kzuj+ectMZsdYH14xcCWLW/mIEql1mO/7tnB7ZUpu3pnl34isdK8oPVHrputxy6rKy4kXcgohkoV
pqbCVeZvSeaNhkfSw+M5EfEUFSTuNTtJEp1OticeRSnF0Q3a6kld9a2EIjZtvwjr1XSvcZmcIpNS
djdjOfUXPuM4GN7y9aHdrIwDhHkeVADa8nhy7XN8MIMVqp/d0liKvVo9wdbZ9WEIdsVzHpyVqV2I
b9nnABLcwr4vAdMvfUqefuNXXvT2xRG8j5UshLf1BvhPhx0a+PVno9BDIKuO9ZM8qd8ueJGR559x
n+GaUGNCwfUD+kZq1YTqo0YnUywwfy1nenqfpTUTIWgzFqi6Ssdl/fupfHNwoV2vOL1dzqNPd+2h
531MNjUYyfUNwIUspryOItkLuzNflEStUc1vsOYJmBOeRASa5c0O3q2OOn+URJxusu431CQhAyax
1YZ3dnZJK8SguCDCI6j6vGZijqk4AmmWEegcDfj8vnVH6s467mddjRrjYdPpMfueMhVZwm4Jqk6k
GS4/n3ZatfPiuzVh8DVVmm2Ok8dwYisaOqTn46esMuffwcmsVGbDIfUKzsOd/n4lm70pLCqbEQoo
cZDxT7Kf1Z9Y3BLsDPMwK0Kxz6tKeQfxSi/job/m/iOvOQW7DS03z1vz7vPZXhSNld80valknJG+
W6ED0RwvmvdVqPcSUIhepoOUcwrH5zNMRyVbIU5gM8JTgl1T8yL0CsSXaXdj5KwakFF19603wZA3
s8rcZ4cJeauhK2VodYWOVMdzNlw4GZtq1fm5yQk8E0KIYcV0OjseS290imX692qa8uWAr3yGUrX9
0ZpmI07Be2EkbyzipoOeL0Ci2wY28bXsaHDemguG9DQEzz6eLXSaQMCrqyDrHgYFXLCSt2a6qlxe
mvhHn6kCcc5mIe7gkwwev0XH0oy6x/kwlTFM6qo5eqRX3uJK75ERPGRIrbVpAyObYE9mF8wATE9C
tAPvBPPdlXxBOY9dEZ1ric8n/YFTzo1DsH28b5atccqh0l0wnczruq3bZRRxO6DYH80Z1QbBYdzc
MrQDwH+9UQ7ZpHAP17QyZZrKI2YPS6w4s8cgVaCgF/42O4IP4HJV5vr6B/ly+haoy9BXyFKcwKzT
c5AdCNcC5KstS9S2mCvv+5hyBDIDxaao6l4RZ39aB4D2TT8w4/AwREbyIf3Ge1C5BlCx/nlhKaYC
6VMUuyLgEXtZxA1i7nUzDj2YJMU7J+xsosfcP+AWc2mIQGZd98jc8wyoOS48f4YhCndfgBO6m+tJ
vrS2VsNtG9NPavwgX93DCDHg/yjT0nyhI2Hz1fTvyoM3L1/SjQKsq14usuETTAFDlgTAQ8bjsW/A
mqAg6a4yAShDNwnhSqcRT3L5WAG+QdCyf6jGs7NWf3nov/KHg3DEXsZK5quGpiiCHG7bYEwj6D5M
/J/xgLxDrQ1fDIwngptVnT2UtGxy+lIAf0ltJapeTTdmsGxryqT7T0JuD1/6uNjRj513D+i+9Rx0
0V6QHGH/ATX58nR8vHFNbcT2qKcWVaMAF1apgJgr7LvacM8ML6Sm7+pTqE7DON9h9M27uBWH6qgx
3MJvd9UoxCOjxDAdod5PSeKUcyQ6yPyPp7MchHLmdHz/ZxDvGWbk/ujFqq6MncXejhNlk9tEQlMT
5TUi52lmPrdbDUdahSxuODsax6Ya2a6mryipz/RatGGqO+U8RO8/wAbQCUjQUdl9q/PaHzWp/V//
H+2fcManA1uZQMA/SEAb69aCk4r/ItZztb0AXwtRgjawgpQDutfptFIdjUpyI3RpACKcgIR+22L5
kmhNHJ8XiWNdNdQ2W6sC71leZmdftdDnGzn31yM19J+J/e7yJQyJtG1OjGT7Wfrn9OsbPAeAKNWw
PQTtw7NneHNn/8vBMMuj0Ju+v5RRkM1/0cgwhJs2AmFTLEGKpJ2ThsEakDPN9xLLofGf1AdzLUI2
Fk5WKHfNJXoXZePRqGAHAGV0UXlH6Zcz6JBIFigSOsVv/xmoh5br0nenoWMl5SDflOqb+4i7zjcD
vlR+0jaaktFaImc2+VIcd9+oZfE6uY/L36FIs5BYrJ0sqtknJ6aAsZqgjDnx1xw1uceIYZJYansY
2q3xldwQoLXZOsF4zVUKZ4GMqV0ADSisMa4sgu8jZYoevstaOHwXpidWBLHtKulE0X7bJhO9fI+5
RN7HndrK/Quivjy8Yk38RrxNaQWc1uy4fhyYrXvx2DLrV8eLXLmSjc1PWP37AixTV3bWFEwJOxl0
j8Jtz3Eka8NN/H4WBkxIyNzBjBEKQDfB6zL0dy7GcozII0fPevIN3t25GJtTWTGDsAdKGHrySIB6
rsYgN2F5qMPzC56vrEiDh0YcxTzXE3lu973L/MYnDic8HHW7My3mD5Jp/Pi2zoj+22wkgraQIz5u
RKy1Ocq/GCmg3OC6jlAN5370CmR6+06woB/NMhQumGSEbCE9xdQ9BJJvtBzqGTj+tHrnEpoYqKiA
t0Ud3ILzxbzu5n4kyTzn2zKGhd5FXAAX9YZ8mBtYogToL78KQDposm2X9xuzFSSzbL3Rz+eMXr7x
N2y7nP3PsypUASpeL+xnbQ1ErnYrVX+/GM2xHt3x8sGUOacWmF2QQQX8V3e7ThTL+uefCteK/B7y
rHHCzTcu84IQv9MIwTKuW3Tdg0S82NOB3zIeHF2b6U6+ndU8BX3r0cC4mCrfEAQ5MH3LI9fLxpy2
q+aEOvjEebGrEv1+k3IgcNdd+XFAyRMzoqK+ERvc7qhseGKXo6YKjaPTy8EqKgAB5yXresjzGscS
HWVCLP8uunUP/R8Wxe1l+tOsWT9G5g81ehgLD/aBwBY9NY15e1+s+/mm3LLhkh3xXOp0BHA/MuFD
oWZf4V1aqXrUqDRZ9jLCbrydy2DCg/TnLWM5siM2wcbgxeBYnTaM6lC/t3w4r4lZBWHD5blfnJGf
JlkeTm/FVOfdnu3+kNeYnKRaSI73goZdJh0ezSz7YU1JZN3wEEQfCnfH7aANOoA08b4eJH9+JCqO
rD6wv8bvkuxRY0iPBmlSfoYmC/ACWnTSt0sLem/3JkJE+7mKDttc8yue0QcoSHYVPcWR5CZsm8w0
hdkyzXcv1EsiW+g4kwsjGKNzmq2M0GiqQOQBd/4VtOGYz4xOiRF2hh08jg6BCFDZ8u0qRt+1hSnW
Ahv0cOYC92ZR/RXdIzK5eP1iP8HVcuZN9Inn8NhDgbsSPFxXIiC8AkoEEnGTxvgVFK0d3V0sjgcO
NS/ZFS2esew+od6E3DDyorFq3t54e615f5HP8uRABrLnsUgbsKM8I2cZTKG+L0fOIdxpaxDTW8Dv
GHWp6a+OwW1ZBoIkLpRQ8nAZOyVT0Y6roGxsyPXxY7nmxT1PAL1y54UPHjFnvPw3DSGyJl6w0wZG
ayctCzXYVb+L3+U3WmL/Qxf7/ezs0Wd2DVVIclJ1Y3nFt4PZ5w6dIMlKzv1jwTGfHZmwzoq/UzXs
1DIRa0sX1JYDO8UHFzvXnl+j0+12uZoyxr+gJPJquilmbDToZZrqShTLRaUUJWl5xhWnVNRN+XO1
969d78P6V/JzlWBTqZxmbHM0m+cxmIe/zn336UToeic1AuCxIAMSYuNVbjD8MEdM5DJLcx9VZTbu
gzzjfCzoujnRmfDrkEuYE07FyaWfTqCX7VOuzs3xhFjg2HXVJkhhugZdmibD1mnLIf2+HAdET/6O
zlaubUv2Efx0vvTqs/14FFJFYsn/pKUI/b0GO7clMA45w8CDj6J+DiEFQSdFcGCNeuDWctTSXhR7
aXPi6ta2z8X3mm9DRnC90x00AvI9ASMNex8RE1EVjvMEEhtgVJ2p1uugsi5zBbOCnzAET1MkNFZ5
NcSN0y25w2OxuQSYC2cCg5Dj5/BcjIfAgmeybhM/Te4+il2/b6tUGLIZQ61CkNKuvT8XRyO93O+g
/cLsp4qm7f7UIwGho9J+x5rBlpqbfiDpZFSZhh/fuwk5+aefPiiJtq3c/obydCdhPD3t94FYR8YI
lIvG+XuP/SqljxnIASpYWtVJhAcKc/WBtABrNnFx+m3ncwcsZq7Z55i6gBfekbWtxZJqwKjEs7IQ
8Ugh11VIGubhYdbngu5HV/Y2uy+yyGCE+VpD+y1Mb5gB6mkkihWGugziaVC48N5Bb8Y2KXsl5mSD
gmWZ6pb0T7KoM2WT7qlxnTjEJzpVzwWA+8CbQS5+on6lseONdccQuUL+9ZvKs3mv6tWRElc+S61l
3juKWqqUPuNGSF3ijP3wzgE8lT8y8jTeq6DtsxFIaRhQV4VPlYcUhTsS3iu9IgiOVHdf/NRMeeNC
jmx/Br4ipJLvb0SRT/JVrP50asu8QEbRt+uAyCtnHGY2k4TqBn3GW+qla2bu0rVzZOJ5+Vg5ktuh
xoaGZVkYPfRH65VbU8tUcDJweoNo2t36lYe3153F53Tue27VeNlnOPz4SVsjSiqyXYRXMHIarqM7
hccZoJHeMmrdBH9K5Ztcx0L8IrW5Ly6vfjhDXRswTgUGHXrKy2z0zopUJl7W/AX8HpiY5UtC9uvg
CjfJgNzvEs+xDQ6+YGik05kWlW3UkpYFf9teU3Jp9xwX+CPk1ctaQ5gOy5KZpZy3mmneiwx803Q8
NfXfL+UFXP5ptNZWqxwa7ViqNMAl8Fin85fmhb/Zh3msGaQJylSnydRDc//DNeax6aLMYayc/lKE
HfyhDVsIKi0lpg99xqLpodkJHqsZU3ThvhgQO5iA1LkEi0IpTvRkXtI/OkGPv8x3TFVXcixTyrQ4
TPiirzi2BZ5zVxvNpNGCOzhhxD0ZIPLe7hyyhejk7WbMv98ZQJbxmNFtKtNHZpRVY8Yz/U+ZSd+1
/TAHA/lpFJ1ij3C8kVaIr+69BcUGOg1VrUe8IpSN4iSe/1985Y5niGOsnSzNfwkkSEfncidteLOu
C083IOHsNIWqcXx2jl5TxNuUTt6q07cXqgPbDZSX+uQwliRuLNcAz0sp3AKU/k0Larr8Aug0kdwk
VT4FTo+Ewe0S9BBWUAqL7ycyeazJAhA4yvuV2T/B59g8VvLsFtVVve/OoCv1FsYa2gHbaVVPwx25
jovtdJTTK9qysunVFdhb/bmbnTE6180YXIQjaApmRpsOnbpC7tyl9/K5pwRWsLD61DbWgYhOWaRi
gwQaX01p54ehIxsmoPct29G1ueZZc28yQaWGFN6UzkHHga4GCGU6WX0lbxBhIZ94UBorGbxNxr4n
ZwwYC1d5OGmhJDL1gEfiZadJtotBWUfLJtewNJ+QWiJJKGkKfKT3OtLcCq1vMKgmb/HJ1XKq9oRy
ANUn6mZYdRal6YU3pyU94X7G8Qgor4Xeg+QMAuXEt3bZkxEKg3ewBJAwiMnZrOUdQAh0m7ss3GT8
ZDyh81jWC0TIAJDpUp2kPiFlpVF52DS4FzJs/fMSMqizfsHEaaxVcIsNXepV2ENSPW99YCDNU3rN
0g7J/h/vLmwZ93y5Tx18vzbrwkNH6qkAcFv1R/7Yn3P6MhmqS6xzVzSV4PnrgzJ+p6CVJfG4qPET
ePOcLu2RqhimWbvCdqmSNFmXT7G7PKG3bPJbJdVI/iJobrzSP2ZPNxaUeZne5dJYvbpHS8qfEysU
DXVCEHlK2/unJNaRXrbZLenvJoUixZ3ZMuWb7/OUfDDh5GKZo1F+8aGHie4LJBMtF57cxv9m0uuY
X6nD9QbiBs8VUMmQH674n9lmp4mR66M02pPKwytW2ryH/aQrK8tYBCwxyFsUWCaLAM2FxSBgDeF7
/kSemrp98YO1gs70WKfIREh1XgOYR4WgI8wProUWDdBM6R9+GesICXEJUv2Pd8gRIHiyCcjIIat9
w49u4RfP0FZRPdeD05YB/zI6voveSHgTXAWVR4KmgZLVtCZjrlotp4Px4RrGVPu6a+/zLNwKQni3
4/Oa4VCaqbJOaa18zXqTajh7AijQfYLnxBqxghGEEzilHYRF580sbOPqKfrJTMTzM22G8Vn1l79X
uqifOKmQvvvf8jNiiNEyhBsScu4dHs5sDPmvrA4CY7naPyy74I3+eCewG9mJ1FWCExg2fvHJohjl
bujUUe5Fh/KyaNS4G7wLmvYj9a4MOwy371ZRW3XliBiUtHO3ozRPA6m5I42+v1fxMZZqvU/1dw1g
uJmoJsQb6CmYcPB3q6Tsf27jGcCQav/XFXiOHzlZ/AfvcsCHd51ngO8byqMhj6vYvp975e2LMD/K
DYUYMqWNRgb4ta4yF8wZRSp1HZBNMabDkiRFW5C4rllvryD7PyH92YmwVK+9xuo88/C8izSoUsRA
I8pQFn9ybWWbs19fcBu07zk3AIXyUaPwh460QsKycuwvOjOhHbpwDkWoPPcE226efNTXo5bSb/MH
gdHpQ/BMxOQI9OrhsLmtp3p53GMqOAKFKO1ghGGjSwWfQiGET6WasgxkcZtArzgeFgG66BE32/LZ
1g9O8gLgXbwNF9k9RbZ91rDsPcFqvg7HoElGBeU9qFyzn5h+Z7hJTs0iJElP64t/oZOTgoodl1SE
YT8EX9+0XlqYylFzkVy7oQLRaR2D8TTyoDrXRqygM37suVwiRaRI2mTJkCzwDaaO5gCwR3M3bW7M
C3QVHyslpeAlA2SCJJ53aN8C9vapjHc321ZuCYTrkuasxAn7/hta+swcCi4rz1ClyjCNC9LTH+pZ
20Htbaxy07q9ad/S+YHbrw1UuDDizQfmwlBIr97vXm/TbXF8vFP4x5evdtjI9mwC5oIolh95BqoD
LDq9gAZzjArSRYVEHOJvj5pAILqJGO0IeYRc9YVjqS1yrost1/F/5hZIC95ENvG53rk+7zcRIy6F
CGoScgQ946IHToDDsPdtQ+7Ipjx0syjUvo0jwnw42U7AilqQh3bKL+BEJ7kA0ivHpAbOYVqOaM2S
63LPZrfGoiu6e4SDDc7BmCDxsJftwLxRIgWeH7zyzxF5Zqe06gwarXebyeTTtUzV1RgiHEmJiW5Z
QmcNuWqcJQ7bzMvJnYXzDmc3Diu/BtaT8yl9bdu59H5e5h8hlBXThXhctSV9eoMms5uDAauz4Ore
bYJ2xlAQOgugiO+3JyQ8RkCQKfNXILtvATuG8NmGioJWvfMvQDQG6c+pnqOX9zKT+StEkQACyUcE
fPBlFy4Bjxg+510XJlSvkAxCCFsHqdcWpxj/eqKlzggG0njPOtbwS5NVE+QNuZZ0fSkU1lffGk9Q
L4nM4soEjHiQ5qfox7w/mtwe6TfXEwVxclD0dXxA5m/kvBk3jWIl3XJVS7OhyssrEeZNeLoLIUEn
d37yLkNeSaWrvlTIChGd2pygc6uu5l+Kml3K8ArvNhdw4VmrRDuV+/A/IxHTKcFcCVrYR3EqBHfd
ZcWo0kk3wxCJTZS0S7MmaGDrfMog2q1S8hpvaHRiwiGacqXcLP+sgkOVoBfvu7N6zLyIE815Rk6b
cOc31CzUt7Bc45Q9+5wRS/aAruRVu8psuWXXZGe2rkGpUZGo7ydNNYTdeCWC/ZGIT+vdAOyjSih8
6U754Uhsm6BRiWnCinBe+6QHbK9HEFJ+AJK3zcaUGviTyZUs+qe5/X4TXBrapNd9Ci/reuvT9kcs
xlnNYf2FiOD3MX/933USrJ5LLMyx/3QXIn3eEff+5DerUuxV3fn6l+1EGQ6CJnzCGXJx/0UuN9Of
SfSdG3+pPo8JrxhH3HPtZbqBZwTpXTXAWrJ3P6YJUuRZVgIjxz8Wqo6U4q+cAz54gqf3kkfXV+Y3
hJJSI06xv8KfBEgvFt3KAktEGj9zEd4PQeOLJ30zZejqLXX2RkljxDd1PAjdov6XXLOu/TWmxHBM
ONkjtXd7Q9euMIbDd+aVAwUTewOXFcaeFIe1wOnO3b/k7wbk9DtvGINDMXlk4ErfBySk5zkj9Vcl
9JDOBa/T62N2gKbrZHnx+ImJIOkGhtWFZhiqsYsVcfJwDdM0MVJ1P70BNTWpcYyi2oRF9H1hweQu
vZ19H+TI0BDhq6kMz1R7C6SbPHmsau/VGrpr1AviM/XcX6gevHKisRMNQ+45hIHyZ0sNK+IHNc3n
xceh+FsnJD0WB8+mX/Gd2x5OPedyRK/yIfX++UX9XfB03nWsXTAFD7DY1iAYgdaFrAEJ+t3IVBbD
v2J+PWYs09YOAAHVL1y/1GJ3nYdR0yQ0ixx0qDl27t4Y8y1qVyhyIJWnzwL99CUjVVlgb7KgXVSK
1nr5oemEB23T8NQwE/31I/2CSajT6/mRBQQz1qQP8x7miI/AZF2Qt2B+BWs+NyVuzDh8lzcEVb+V
+tpzcx9m91u3D54PzuQRijibwcR0vnqfJyPlImZEFsmxMz9+Jju7K7oZH+X1U5liOrohgiyxeWzD
VnCgEQ1parXr2O356nyxj4v/QbkDWMJ4DsX+VKuVZN5MI0CwrEHkvXZ9kyRQsgHi5eziN2EcHnYL
5YWYboixRaVGbRTmlNZsUurJ1xnMtJYzpldtyx08YETtwKf/2VV3zyXm/bUSreb0sNdC3wgieQ69
QCQV/KAz3NGkkbfPTesGm1wkcN/CQZL/BX7D7O+j/Sgf2b6rN/u4/u9B+5AQNv7yCM+P645qf08H
h/xbzwsuVcxaAInY72hxTE9/YdTFa5MSnNQ2OBQmAQUsix2hltRLN82AjuBdHStozLaMIxfPqbaK
WJbkABi4tH5RC/HldB0z146PQq73kpVOTcbNBvThyBqRyuS2eMTEPoJRbdN8IvYxy8ULvRfNAH5G
FkeYlog1fg2jnEk1NU7Uuv1qzbhvF0uTCkX5THu4AEkB/zwhDOOmVlgLiafWw4q/ip04OF0iPGnI
zDXkBkh1WO2PnH96nO76Sh+B+1x92Rhs+FtumoRypvo+2rlJub9a3G4kCqe0kCC53pcAwzIDcr1F
yXqduC0bhAIakBitJvdBbEH7DWajs9tZfd2yydmgaUHtQ5pXk6BrACjlGmSfyZ3TCJzK+kzuM8J9
E5t4UWTioJ0fOIsuE404GtrZhEY9hPG/UVXKyEZrYxvQDyxyl+p6vMVq8w5CzHp/d+KOGMxKnXRJ
KXcPZ+gynij/ge/tJUIFYMOrn7aP5r82i9S8kO//9dfMHHhMYpPhql9DjbLlOH3YuV1LqNAHuch5
mJShK3rmC0bTMaHPWpzduS+V3syxtcZmyLGnMfvntUKkKQRxPMY1iDh5uV2DNHKYhtqi+CQfhZeQ
Vl26Ty0J1OM4oW7GDcxcXaF/7lJ7a9Sr1ObmErx9ZdTR3JSuL6B4Qc+4NgQGVNH7EMmKRbR9YDx7
YqvFFFvBRn/gPhM59HBAHdRQ6Py+Q0HqGVin0pBTsds0R7+xS+YYqd56rG/BXS83YONhSFAwkYGq
Su1RLIoYTDEAHPhQiSkbds7WIsalMIjCi3Jt3Z+In+aLSihUxAoPcGxw26jYSZIlO/u+tg4X4SKp
dZQYt5n/m4Kc0CN/tCNSlBBx0dj1603Tu96/zwpbDcliuXZH+tVGMXY5Z/prLVGPMrBZcovWP+IB
uayG6DQL+9/RLY58u4YUXTvSNhvH/nYlE/Uw8tFyZh0WUToAsqJy9tYtFOJmQfTIFN5zNpBjL8UJ
3LcgKk08kQy3mVMFFoNXYIEsBrHkYhVzYIEUupRKH7UQII2rGCWwN+MVYChW89b2y2gBAdLzm2nc
AAJKGUWHnhvj2hNd8WnajwaZlNGVzFqt8gpoImT2heZ8tsTXLMZDYBYcQzQnXILAkf48SPZZV77K
sjX9BQOhxyHbHiHx6iT4boAxP40p7x9jhO6cZMwrVoyodawosaxNcEvACG71kSdCE+kCqGNc1Gqs
FssTsPwDdlQTF9nPq6UQTmU3Ph2zE6VuxwciiV3Lz3XQP3mxIEzkvws0Sf3dDkDKFClxiub/f3XM
OUILrXtZcYc9RmEzJnqKx+9BcL697hzWMw1Kjr7JZM6UOekthdVCbjtKuLmCGaThu/g2a5l4V1fp
XmDZ/XcfJz2S5Fcv6CGA+GNKS18hHyzFK3xmNFQpfuylH2M+qiumVwQKIr/DpRFQ/yGdm36A5PtU
n6YX5p0PlqlI2VnouP5Gg0cZBqxOXXbaRNsuG0PE5/DQuKL6/Xw6QejqtTydkgo1preS23Y8l+yD
RgcVL2iRGJK6N1ksbeATtujtD+7E9m0JXP0uTkSlFncqW2hSkEctBWdJLfyC9GelU99rdaDlcOzP
/OZfOzOyDeXnoZUVS2Ta4ExGLcigN/XNeEBoeKDtNObgIpoPSCwKdaR3nW/hkNNLktl1OyK7DF4p
2/uvdm+UFMqhcHd5KLQW1xAQH4kyQnKHqzJM/2VBiJXdf6xYWhqHdlChd0nKBDuWtwBeuUd3k9Wq
lf32xbxIZTV9EuEpqn7tyY5IyDDkjcY2jIZPRQKX0Z1SGentAfyRe22CROumEF0lDJ/71l7Fv1Kt
2bzs2fqXABoWoFhQVDLVVp1K4ZBGYMY7MbNH8LhnGvroiW+GXESS0GVjQjTlAjb3VweKNfI78TvS
EbwnLhRUhX/y8/uNNO4C2loTqw3iCbETjEMwIfE2kS//t6Kc+TZBxENDcPeJHIvCCW5qtoq5aRFN
afcRvc1NA037JUqHvsdT5N76mFOPltmtaUqXubniVMEGvCT3aHW4w1xN6lTs6DUeRtQJdTkqaVdc
zYfGuPd40tlYxpuDTPApfW0fw/zV3I2zsbkpO+3zrcmNVCjyl1UxzEhfZW4ApPfv+qlOXDntQaJU
nAmpAGJzQt2pMg3kMwZx32RQkX6w3giaJpMJwtNvCzPlbQtF9N6aMfTEgefXXqxTSBQGmg3bdxR2
4xKPrxaryk0PJY11tPAu2go7wYWVAiMz6i7Sruo/bEfK9YeJK42p2/6+GTapGoomKsu6i7DR/DTm
RrsRWU+Gyi+9yGCbqOuPF29EMcmae6LqeDs+lGRCuqJ6SmY2tc659+FfYFASXJHyWRLLYVHdUnKV
Oqfg+myHIC2wUFxROKWpmIIuLolLhnClYL4MhjsSAYT+u9HhV4Qe6B4TXosj4qkYdv3VBrcS8iFg
ELqyMrlw3tJdhId1r11w2g6gwTNBJSz5bfHDUs1awiLO1Ze4WqKetWYg7lYSqWLlzCRKVQFTWLZg
D8MrkY7zA7uCKcDjU7uJ9p9xGA5TF7vvoQ/sQjcx+ZmZTObi2xq5XtuqjFzlVMl1YaUdc46yxzH6
wzu/n/rGpty20UKcrZ7xj6mzBXPocfraGsveRecd/fnF/bmIL3t0SGJO/O/yaoL98vJp0ro3CL6/
QW4peJNjv8NWKwCC8zzlIxu+H/UOVG80a3ihHuaG/lj8XHRe3mTi1vDJ4kYyRpPLbLu6iXPNQPJM
m7vgHNK4UfLjOlf2/zWBA+sCHXyilsxb3fXOfI8aOnTjczFXfXuITcojk0gMiTFYWK6Os5g6Arzd
65ob0YgO702WsRPxQH91iRvi8xb2loRoEYqK4X6mZPQHypCG4xJIsR0kQ7/K5iID20YF5tO430GO
ntCeYU9+BjYmBbV/q/l8uRPifatNVIWfl4PAu+/pu3EUTcKcAyluHF/sZtWk6FPi0hZQELauBisp
O0KvFjVrd36iZN5v+nxizkXUNN8onwKr6+t0untD3Uu3wFCY0AK26ngsuXq1iw3wrgAv5klPGNPW
+lDKJSBTc1vfyhVy1fTFYJ9U+15iPneAVGd+TqVxcMcxlu6tnRUPuVW3bSB7zPNHxjJDGD0m0Y10
IIEPqgV/W+Xfj6iZrGMkyR+JGKG27QfXDDtMfbWQ9RJ+2wCAo0eYQ7I5uRVni+FjgXwRXk0LMcb3
jcpAIjJwqj8npZykhpL6ncXY8RGxMBa9YyZLz4TV1Kd/6e6SkoSLmkHvHzfnR1gs3rU/DlbyJ1VM
ErvFkSTMwqOuXhHCPptGRA1ZhNnEf8KyQ+Wv+rMOtDU0HVnooDAIgs7Vgcx2zOd6aOcO+lAKwFx4
Qw/cMYQlYgwVbliofs/r11rqEatJk+oj6AmrMIRmWWPPTFNbPU42r9ZZJDFAwXEZZ445rAdzfW9P
u2qBQ2ukpq4BHCU+ymxR7/iFmc/6gBFUrJQQHLdkSUZ3wS5tm3uuR1bOGfJ4S3+cBUlnoD64P1Bf
Nisk+CTdovTSJ/eB899a8/ORpCJIh9pjt1MtyS2RWh3MrbolAnB6/+nqvRaettxAqYNTMMFeFRdf
KN3B3eZtnWZMjNqKt8W1n5dDmpynMat2XtLHy0JlxOX1Es+8CaQ6czq3jtFBttkCBKLjBFX/UxSR
DTsWv2HU6Lak7BeN8C0eQznVpMybxjVQ+xf/rAHBquaReLOfb0JDaXkG9DzU5biGdclhtll1Xms4
KZfBUEoLpYM/6Pf+Gx9NFRp6QGT5anOmExcvj6xlL9NThbV4CBjBbqD+AcDl37k5RfC2eC2v4Y0p
kdgl4Q1XEQW6kkK3ZICRMhNbQYETdKvW3EwFIGVa842ctlLw20Js1m6069YWqWEfG5NxQqByVH5i
R/7EaaSzxBLiibDd63b6W2et0uHuTK1WQFxdhD1Jcy2JRWYlom06Ke668fYM2DIrMOChDf+hhtd9
iMhPgNdEd3I5ThJhZAb2Wp/2Z+dMborLlrH29iSJVLy9rAv9CHuN6t/jitTR1u8zWaDPqf82KeIF
xWdi02tF3shToONBHeq+RMfoaLm0aThAOrP/NW6BLRL/X/Tf9qCx3b/KjkzmDSRkO0uXyD/J2g2l
XrZ838RBQb2BAZiCB500XzxtEQVFfmH3oJ/1tUW1N4cNoBWjW0udTk58JUHiiWujR/df6F72ILER
OzUH60mPWZ5+lSGdC5eaZsKIDF+67UBVSeBWIaUWUojzdqADfrZKO0++GT+NePuSKIMMWgK2rPeS
7nhIXTznzX/3IMnUunfeBMK3tAKzJlgIR2dLAb9uvnucDXds9BHB799Z/C8yLzLnPlwerjqDH1Uk
UcG5L1ss5Dmk96OtHp/WWKmHYURPkhGAmtsJPb8BZhB/bOXZ4so1I2QWn75IswzhHYNrkSpbvxa4
K8gI6jpPggXmaoV2O7I27TM5WGM8DZjLd/hJoAl27oK1UzUWYQDMUwmnTNy+WX0hJzLHbKmz27fq
ZVmICzsMfkn+5kBC0VNFLwPLy2Eekp746PyNFj5h+4kFjPnwtrSHphsV23rsfj902+kqlQRXnTiL
Z/BWNR6OYW4NMagJs5kLgaD2jb1OEb/tnKDq06FB3E8yRAtllqI2QllrpbHWTZz4U97u7QVsPj2Q
I7Qem9YD0CTMOyHpK9u+oCbU8M3z1lLfRf/q2ACa693IN1T5Pz0Gfjlq/XWKEbyA4+YwSHrotpQR
xw0LcjJPYD8R2naPXE9gobYryHpWUeR6HW8AQf3HBTCIO1+EXWGjN/99/3l+ebvD3ur6EgbFIIYg
vrQj2PD8Lka/BtTadHrcA+psf+KUcInZ05P/VPZmzp/CzR0ghjBVT/8/DdPwR08IELjdCYRDm5I9
F5VI3cCFuPqqXsRHlcLdG6b7If5gQFe+ljdoMZfvcqBdhGQv4t9MNDXvrDpjZMk8s0GcCjktljbL
DiFCXABGPM14bDU47GPS2g15X4jg3JqMe5lTR/iByW+1o/Jydnb10YLSQsLZ3w9OM+uCMjnTduNX
Y6jgOWM3qFImzQ/oWjJ6jtubYTo7yQ+mNSSlfdqV452kib8TwDxLTyP55duVxl+naWu5ROFPYu20
LMHFkzilpR8WTZt0KHDUlYHCd4W+scXK2/0hscVaIdQ6fiIRiEkj9K4P897S2ToZlsx7UQ3KMoBE
8j0/Mc8qSGH7hA8moMtMak5xr8W5dEEUUEQ5V0LU6M5AQ1z6H25N2CF1LbpchKHobA1xxo4nDIDQ
DoBQH3voSRnGxDlhQ5rD4kqnlKYqp1VGi7s0khRMpPcmJ7uvvOwOzoO1mX+kXb/iFUDsL6ygDtUh
Rn0bpC649X3VywnAvpv67BhlVr9+JEdvWsLc7lnO7kLm3+pb0q2XrPxgdDk5C2YnYT5dFqVZ7hnN
Zn5TSzW6BpzkmfNHwBYcuj4LDPZkywHIyoFDQB9YVGbvVSTLuJF54vzQ6DcGaiTyFqVlAH85VaNL
Y+NB27Bq2Dvq3neV0fgoIbP82WYVhUaOz2fzG0jp9cGd2JMLGl4rcPu1lES9tt1GZqZMdhZvwKgo
pucq+ajUOy6VQSqIhTPn3NRwWbSTMrXif/l4pArdtYegC8vq8ozvbOZUSebvnqHoeT2GU1O0rEC3
zuNPg0L+4d9OqYoh3UQcOU0lUB8/Q0s5VHY32iq5Bxbz2mJD0TLu8K/gtYod3HoNIaevmaKu82UM
H6QzOl8E926MhkYZJRLbMIwdhxfOr8/NINCIFv84hA3PB2kg1h2WGUoEB1iT/7OUoNfVfTggk+CZ
OS0Zr3t55/6s//lYb3WcsIiQ8kLLnEIGQq6Kba/CIXbLWhAj3Uz3BScV+dLdfPgsEwJXwuRFTsO6
4fndWjUgxz20mR48qjkBq06f/J1z5emR01Y50pmV8s/BRig7GWul187mtoev5ZZZf7OPI1bSJG3C
TLF4j/E/0W0wgEPYFu0fBMnCkSBv5Dp4lvFJAzyQVOYsgN/03J6EBJU+T0zg8O6FPclynEdmO6m5
+bVvH6ZqV4HOAa1f8ItM4okXNs23l7ko72hqEk2joP1Yas09YzES2Wjngbs9lENdMnZXZrmkEX54
B2hjgBG0kgpVh7MceKf7zx1RyE3qfrOtiyenDmAc5Zi9N/4lrzRm5w6V4iVKiXhlkNpfV/cNlC+d
TqENNOGCwLwmAdm1O6ZOZYM/0HWju2zGQYbD59k8ELZBCGfTlltN+T94KQRUJZPFg8RvBRHfgB16
Xln+QfF+LJonDd5KDt6swYgGRXJ6fJGRml301gZC4Se4isSvhFcxi0F5UoDvz79kKdWrEh7nYBVG
a5adBN7v8EdesQNG6POp29PyhnKXdxsz7dBgXWybApAepqrL6wc2GDQU7aPVM+tjHIWfekuD4MOo
Kx1Dx0O6z7Gu10MxtjB5sqcNwk3xN4yevLYUSurq9SjaJiQSeeISZndRmMjv/vs1gmfUrungGSzK
4+ghXmCmGAhNoOaug5F8Cb0U16aIB7q9CUPR7CKMbiGxtv4jE2ScBKXOmRAjdjJCVIWInz3ex5n6
ViaBrj1TMENn26bJDVX9eCDIjX+JEpMFOmcQi2mRpf1SebsNd/d0/PoHL05pM/RldPw00e6V1mFx
g6bHqsuQeSbUUAzxAAXUyEwRnt8xmJzbecFJ1sFKJNHE10UXOr3chkLx29yqTedcBCM+qPUDPO6H
HfkLjjeT/kfuEL2L2XUoXOM6qmaIHCKOhm0Us4r9kMsone5SkhvJ8HTGUmC/qlKcMN04pP7rxoIk
i/gtlPHs7XxiLGmogEptRfyYOiUHDCJhncZ1rQxbXAU0HrtUJrg8umrjAjy/wDP0lBwGkuSwN6XL
nucklxBBEx5WJco9iU4zT0rpPqsXW26AMku2YzB79XpBGkfJlNgT4wnyyTrg0M3VXsuy0xWb3vtt
yzqOMnbfHkFBXVYNWLMZ1VITnGiHKzxat6cbWbLNXfctJRXKWR3+MLciksP1Fb5NOyP82xQ6G87W
ZkXCJT9KMe7subcy7nzHKXiGfVcBwd3wOv1zrNejY3ShhSp0O045Z4Mc1yB6AAX7huWQ28m0rLAk
MxIoJPPcdBvYWePOHIYInWKAcStvjHMpMJ1PbQt0wfg1Yph3qJ7nof4DUaVwVQ7TBCq4tV2Tcblv
ZvOwTtnJGb/ut7/cTjnbSBalSus3oed8iN6QWwP/7rhCQlDS44y7QbntsrbvNjXDNcpLEO0zeB1G
ml7hoiPD7I7FBCVIeQzB70W/aMlTrWz9lRJTMIwXGmVjbWdzqbj9lMOg3CNpQeW2k1PG6RU2Lm6o
7ZFxaLooqtg6r2LVetmNYanGt0CjRvL6h3g/fju80Vn5tztkfomlZEr4nv3hGp5/FOPG8v4HnQv3
AJRBbXvbfNEOli+n0uMisHkdxqohrZNqXeZTWdCFJ3YGfwxRfv9tKznIC7eqwYJU/UZ5vhm7xish
w60d02rvE0dUkhXp/AEELRKW+FUSwEoTO6FUl609L6YLhk64dXOsvRE5tN9NzF45ELPbjZTL73/W
FokaEbfU9oeoELAEH3VH7NkVVafbbML1WBgSj+314n7hA3y/Zs+Hm4UOGymtwq7U5xexLHrlP0Xq
dO+y95mmWMtSNKPvhhFkbhKM0o9wLswVtW+zUgcbiPo2tlx1XxiHR5jZzpgwGsIBInODlTyjG6wx
RpFvSARS4+P8BBs5RRR4xjZaBRQBcaJbaNp8NudBYTYDTO57s/VUjuOvOVye9EU5QlLKPeNnASbz
2Tq/oyy2sLzHecU9Cfz9eWW1Lxsgsx78vG/lree02Jw2YBXP5+ADBMYhE/0jluzX1m42Dzhg1HBh
w14NhJmOhnuArVjwRlGLIiRXdRDgWIaSlVVaXjM5LsAgaE4Efh+4UzkhfD+Q3e7tZCSbegBQ7eNX
8CldQg7SJ80gsglo+a42l0Ov0pzTdUjtEHNCbXqCouyFp/P/2P4n4kxrR3cdFCwTTAdknZ/7q7t8
sAJpfvVxqumwU/iBsS+SkQ3Fq4ScUJbhnCCXGO6DxKPAJFcjdN6WwJzpGJdQNCt9O87hXTE5uuoT
EXdbytDqLjLkMheOaeq2A9pCW566+9DidW4Ij04IOnQqH6AuOpAP/EYQOeobPF+QV5qYlDedrIJU
08/NPmBb/NdM1XFmaVh7vC7oNfKR/SXhDJnpG/jSkCOQyrRt6iW4QNbU628vcqyndLTk+LqjUNwm
9IbgQE1HC6MMQXECxsoW8Bzw2zuo+/3oXryKhx0THoQxPVT6EpA6Z5C0xngZOEU0AqSRXdWqhxXt
NSXDbH94zgdCcisgwn+EQYBGJY8ClhzWDPJsdhIUauWMYSNJZFkfJE6GBzFybnpv31SllNLPC+Rs
/SXh2/yLH1enCVwd40Zl/mgIblMDO5tEgjWp1zdewAmgYUt9W2oLs2KXd4e0LZRQNb2Dm5O2U9To
llmNEbbfdLZhYcLZvkReRd5YSbDmyrZHACQRrb8meuZjjva7hT6P4CM9ldtQD3eGkV1WIroU+fid
FyNzB0Yl92/PTXpSIGqobc/YRZqf+YSLI+oe8eVtPpVndur0uTCzsAhQlli3LgxHBv47Xf/uFt4u
OMsUgu+xdFL9N0t4ZaxUB3YlLUGKGQrYtBUJXXZBaUmd2kL8GnRZJ2aiYgbU/U9Dc34mrd2ZVPfe
Fr+1WKZ/WTVNNxMeoygqs6I05idk/WzX1CPU+oD05Pp7mxU9sKyGuvs5y/4sG90ewJFtUr2hp8UT
gkA8TmpLciOUEK7DhuFRXB/B3bkuv6ffPhtcyj54wWpw09c6kr7GCc2sr1GA6hulBy58SIwn8Ymw
mObjsfsKCkBMf2wJmIV2Awafvq1Y7lV2z4yUgeW4kel2vuB42Nr/lNXMRn55Ap55v0TBF9paJOuA
+dlBQ7t6M9xvPmTf1tFNagsQod4ZQSxrBUuTsbh5qXZTNd5/bdeMkc1QpRn0/DouKR5YBWc6fp4r
13JnCXnt2P2hq324dTdcI+nRpgW/NJEjvmGeEpuPojYHwvJOlUwVi8L2cbmutp0ttl+HlpmO5K2g
LV3Q/Z+YvFqvDT8taXtI/QpfPugeOtK4noP5leKK9knNae1ZzjvM4jKPf2ufpZZ1ARXGYQvQh8NP
sgG5uv4aekffM742bopISYeL4V5oj8vJAk7F8Dq4ZpoUDiHMYm2qnI6/M1Fwb4nnbwkpK2brBD50
R3uKhPwTxJdE8I4vCUvNex7NiFiZaEYYfqDnn3BO21jWvMbTcm4MJqWi8RdenTJlHqIigt4Caw/7
F7tNbW70e6kzH6GFkesB8DXc94jQ20oNgS15UOLuoNrRIJ5t6aiEzcucoX1ALFgBGsTf3M2erJA+
sb3URg0X+sjzgPZnjST4zLuyMLj9+V5/eQFA8ZiLgHYx4HlmF3Gk3X11ht3vhWrectvV61mSsM3w
6xeS+QR5mOYMnS5kIGJZoi6GCoPQ7nEYPy1XvekD+b5fbBjafOAj4ikcKwXriPTV7Y86YnLKqbCB
ejULbT1pmJNjnHI+6dFvHjSKX1p7YayBFrTFsvE3JerFEgvFXr0wtIPcEUC1JmVt0IeWSTQrr/6E
guhvnmSH0A5diO6NG59GUmH0fbPtrM+oHZ5zWjnHYykdyIk+v33dbmbnJg1w+gGb82+JcDTtdlZt
/kL5SgsBYuBE7c7Nm6Lv98qZyxTRz+TZ/p4Culbi623jLYUZSa5qAyRZ+igtJIODSNzkeZE9rYwY
Yvtthn/3pvM8Yb7BNBhmpKeqmmPCgK5cqBGXmYR+AZC1jZLxBADCoTJuzunCm0XI0c4TxQO8LTm6
zXgWagb2Pz5GJ/ibPU2CF1yC2EynqBW8k66OsELq6THT3kLMjcE9kaDMjUYbVaIgRiUqUaStwWrK
guTAJK5Mb5vHVuJ8hOlDiIsV8jrl060VQh0lLLB5WBRU02ll6KiW68g3riVDe/eVcMbaba6KLOzz
znu+7Rz7Y9qi9JLy7GiY17S/wESVIPueydBGl6qr++7WY1zFuzHIF7zVLjLzSDmLbSx/B6kRkpXm
3rpQvFmvMk+wZzk5RgAk/TguuQNDGB034HJjUFKrn/50euC3y5Tiw0Mpj9w96DjJ19srqDeDz373
hlT1XaWbSQA8lj6ezPidAMkR33qaLebFj8Pw3TUH0CN7jRJHGC1jmpDdGhKr+mAARPsuK6gHopn5
ljxGm8X7kKMbpHKjPy/GLwtRidAkcjV1oOD3hb+AF6MQhzOTc8sjq4S6Fjx7GHJqGMuPVlX8LZhc
kVGe140N7Ej/Mfu3VWcKONavMR5ExFi7VEawGyW2Gzroi/TqI4zUwzDoc/caZpiHKDNRJpWJpwFy
yI6V1r8I0RYfGOL81NF0Gq2SUhXdVZgeRsYnaYgm8PS2gQer1K0TrCMxHiNckuaDUf7ySL0bKc7l
zsMCRMvFzn5Vb/NZVfRR4fCO2qDQtRQkg/PV73QbRjUvzfmSP1svI6b7WVTB+2cUaGec9dTNhD17
8LCnyrOpxytW/ZMRrKabNvmk6n7xQV5ylcgmVLmB65RUk/vDm2yGLVFCAFOYlcANzjZv9TaZIjOu
aRveP9x6LjlQGm7Yuncq2E17od2LPhNsVPL6oxRbOUkTpCHQEdvYiRasT71EOD0Bos0ydzZmIeji
OH0/06Zn1YmaVTHTKCRKgb0+DLGDuDEW2MQaevGKNzOFQU7Vj4a7A82qGGLeCRUxCnf/o7fuhIF/
xuImYwcCaRSbbhqz3cLcGeY8PvlRv4t+/9bpjSx5RfF+JfYt4eAMzHh72VIUlR1wFTLlI/cL++Rp
pMjm7bkyfPtzMZvZyWYldOyXHz/Z7UndkCzPbebrB1TWB/NHQUz9wSZSmdjGd6xdddQKFbNtY47G
yD/L+wt5KIu9RKmnKtQFMRlS44Q0zlCNNXZuYXUk1g5DrWILnGSMtCocMIvFKyTrwYIMbjUJU1OB
sGvoK4qQY7E3CWEtHU6WfeDSWwFq1EQ7Y6/rhQ54e3KdulTiJXsyafm2FhYc3BUK4QC/cQ7Q6yl3
1nocEq9kkRFNiPTGoDc5hIX0vmLbNKLzb7HLONCpSFwQp574qm2QO7TnYM1FKlcDeOwYjWQmVIw/
oK8SmurwGmmlRkWmOg4kNust+LnC1umaJbSDB54aawGcPjaDl4dGOflQd7VJERtWIii7sv93R+k9
hRqqLY1iEOY5xQOUsw9KAnazCC3NB/V1HJZvV3eVOuCzIJ9isKRTJ0vR22qhYB8zWeGYsi+OAgCL
rfb53gubJnG7Xi6COMjtwN9csir9BmwsWNViIw1PKVBdy0z94dwdizHJzBlhYa06wopUBeCd8vzs
+WRxDXdYJD8C/9pPd1CgdIf8iXCC286KDResBbqdSJRYgL4itZHI1ZdRkB1mTtiMFR0Pqiyp/TS3
O+qf45DcR/mt/uZkTd/FKkiLMrfrdKmA2Zl4By6QfUiChINWBkTcxNWNYk2xaBjON4qe08SceDLi
bTaEcjcpZ3ddYTVmuADVogMOQx8RwRmkzOaVnvK6ja6RREjVpQuep59qrxuF0mldnX0lms4lXE3N
aPbcdz+6PqCC/vU05snzosxQjCGevnldh1GcYZCr/EpRplX9zPnBMdY6kRhXFXAl93VphGhrp7Os
xsZFZF85GndU8+fuVhs3UOldq13bXGl9+Yqra3siUlhDkOhTk+0r648g+Ul4xRpOvzqD20RR8QIX
8Yw9uLpM2oF6ySo5TfevupIhUSf1UiCupZJrdEGzNFXm8YImrjgMeUbB9oMc/hcWo8ZNNmP1uBUO
ve+i6OWbbEFT5DpuSQDaSnOxXoMtsL5/KGtgZGvvyES0Zfn9u3K353/KMyZaPY04OQzf6WEaBqZl
F25P9HTltB4/AiQj+/RYWlC0c4xKN4Lgq0o+PDY3ip8h/6JEWI1JzMlziFqs3tmylGNdWiGa/UvM
StroRuTyY9BCE611OQIWwBx0cQKMaHiFSL1Oi23XiZBPKqv16Uxvo8PzHZO+clnq3My+mLzRWBt2
EASdbZK4xqb/PGuj7dB2tXrUiH7NoD2Mw3FS1rUo4SDGngmgU2iDQok0SPViDn88UTWDLkxlJvXJ
e1E+6dvl3E3X5gpwahlBg2tPU9FXZZ7kW8SL4wHfkbZ5M/0r/aFV/Iyvu6c2e1Px531gvKVNRe6b
n05rsLSbz7ku8+P0o2/vzLf82YkuBJs+86kseiWj9fTeEBYqmFS8+xHeguwta6bsKDNiJbquv0we
3jpw5w6lE9TGF1Xj56L5B+x0mp4s1783O4iq2A8l10W20aOdWzwdTZs6aPAQKEdxcLTdlNQaUhe4
ywMZNz7i/a3wfpBlINIDP+fl6uQw60+lWMmCqK1fYuWuSaSQNxYJ/v2FdPWx8o2waaI/4ZUih059
dRVkq31vHK/QaRhq3v//InGIbHSB0N4GiJ/fXL8Ti1F0nCKqeVoMQYYtadYdMITjKZTFtgynGHJr
zsfFkYfB/ExiHsHAaa5W8R3PgRSX9FvC2WrpuDZRMmw2eYF7pPLd8VGwwbX9UdADRMXdfb4sEQc5
CGlju9A+VQOu1kosX3ItUBxWenlRTXVzP3HAxq6Pri06W7uMb8o08lDh0ZaxrVu0Gk5Ey2UmIWu7
drInr3dYG+kGj2nTPW0IIql2MO8cxyQLtFDKUUwSmNZv22Iab91z/21DkG2qBcDEnZAI8NhxVK3I
qSJupSH+yxhW6goomF6+TBleqBppN/kXWwwzRMDc1g+U6XtZ0KYYv9Zv17PilK76ZZDpTGpyH5lQ
P+EvcfbkBFC5x+dMLwvL+u1Tcmv7cM3MC7Qi8VpMzQ3IuPMKY+JZh/8i81RcafTO0g8ZPYA1KEd4
fQNuWMU7I+R7nZoVqos/njCGfNoShNVE4cbcYY2X0xqAIxgwjJZZ+YHvRrSmggkpb3H1FSArDR4j
CVACIbIqeDlJDI4UHy4YF0NPWq7k20K6exNUg6w8UxZz925nn5F8Rj4QCeLHlKDObYIDl6Q8GyDe
0O08fO3gJLw8vr+nopUBut5TFL0GoJey2Z7NpLv286KUK8BtDuB1Rbd1UFnC7+nXaw/2pDaCWbC1
Rl7obQf5FfPUaJ0ixcmyGFwRLxnd3sS106OCQHDBf6pyZQewXdBCHLb3tlP/JCmmDk41kGf6qbp+
Ud7iKxFUYgTG0pwZ+fDg5sH5WkCczntkiseir9923rX0M21amgpnL+sA50Kq33zfkor8Bc/gHFtD
22yFJYUnkF7LTW+aqvLXv/knavXRyC7bSlH1pdEQfiJw2+k1QJOmNumkPEE4yJufsjGwI9gr9lhI
LrnbFf5wwT5uCtR0OWl61EZnQ4/jbhzQTBFV8nRuWCfuZ2tARQJcX4ZFTap4HGM34rOngLACoXMz
FaghcH0pm3A5oe+aOlqupG/PYW/L7UJz7rc2qlM2+S005cgG9CbKXTZTCCoPImuoA4vXEqcBh/in
sV3ETF28Bpv0R5MJl7PzF7Cjq2q+bHGv0mYwAaT+hhDOkMVI/zcwTe/NWiIwnbf8BKxYHezCrvEj
G1K2/9AI+OojXtzKGMS5hUqPIm+P0984Fp5jqnZMDEuHI8Pgb9GnLPQjwh2AJyFmyN6/Bd8UpRfO
FBTHPrSO7ja4ACU6Hj22cT1DnRzt9cYLx6QqYI4Jnspjzmzf3FKt7rR0++Bc9yUIerwgI9MsUJlP
8haUrRJaBck5pL2ylv4h7eP/Hq8loNyt69ZSZCw/KAhyPkz1Yck7sCPDineoDFn/dILeq4AUwhzA
KjO0yx3IHae/KpVD8GFXcghrWolALFI8ASelE/SdnBkxBUjEIALHv7QSD+6FsAdlr0tlNBVWqRAZ
4EPU/PFGkNhKJS6ImcRTWi3uXpK7e2m1jEWKhvP8GIBusbRdEG0eDAlyGM2KgjmjFhOlCmPPfmZV
N67bwRblJEv8yHZBtdlJxmUHwyQ5EPwo+TJbI6R9IMuTMTuZt7GkG1TX6LQxwDj1U+gi2V1G3MxX
YKZzzPQzCiOpaoOfCMh33fvEAW3VI9H6/iPFtbPbhyTntGKtspbSZk3UFi8hq/8/THmNz1AC/1i3
V+SZtIyMCoCvtotbNCbXc7B9h1HJEHcvBgk+HcL7mNxzmRaV+B5K5OWI8OFnUcyonwRbxcLURCar
o2GDrVU+Zo59KfDMXfbi6LExO0P5qsE8y55Rv2N0fCLUlOJi6iBHgkwGUp8tqyDWj2iaJ8M0g86S
hm2xYbnGdSndnDiKSKKQA5/iH4+kYFo194g2sODHy1wUMNsFNKrg4txU8SFhhGeYstv1mDsHGpIb
YM7AalQR1vmoQNAH0lU1CR3OOCVBtYahlwS/1CkH+TTKHqtnT7bTxP1E6DsUa8Xz86B/JhV1sXEq
mHdL7UW8iWrPT5WbPwAQKv7gieg3JY+aOSqGQWkLQdH8SwaV1Z54AOM9NA/vZCuoCgEVExq4F/vY
HVgRdfNS2pOYXz6TekrdOTCcpHlKIFO0c2nwmxYDk1T1xT1MZqTd97HK8cqagoZ/FnBW3JW27HM9
cfZVT8OrQ4GXURqAjA6Waf08VhYzOBE1zFpOhE3Oytz02nx9qunQkutVuQ5wf+tCGR78gvWV+ITn
+Ou5NN9/9wnNEon3TWo6i5u1qHnuJbBC+7vuq5+KzsM/+CgnEHeTpy5KeXISRDbxDAK4T6XliDUf
T+MeHSfHSczZvSOhglD3Cw+fQ+cKjn2jCwsieyZRobzcWeVDNlykTrcCcu+6xn5KPb2abeE/VH53
1VWR/OWbSvkSmG2S7LaZLfrpv6qwSzdCPJGbg2e0FIOv9iURlANGKINy8NPbOsHEOkk4bNZa+m6B
z1unVCu20Ig6EP1lH7mOGrZCaIzm8YWupAHwCOiwuqqEIgWiwNJ/LxCY4mCkySn0mitKT+V/CvG3
RCzXWz/Cyc7dyTje2Yrgsz16sq7eFuSqV8cqMMyZESdaVxGKwLac4Xk/fxRGwWXpWZZfd6tYNAQC
6kTuznhF33ZmHg0qhVqOgl97Gvpt8VGG33J4CPST4pUUbp69iEPBSso4jMpPnT5YciaJTEflX5eR
V9UCpc5ZR99AMseJkmgAorhRPCeHSaMygAW7yY7SnagsxaTeZzeuWIKiPdrZa7/DYyHLXlcatkE0
VFdSK1M0BzCZRXyb1RpSwa7hnKpKaa9jNpsghaMzJJD8EX1y7gVEXYn2+ki/eOG3NiNL5Mns27hn
2dC9hcmoTp8egJH3na/06jx6G/ntF1uwFUvKrOTIp1oLLfCBn58g7RAQsi2XoOQL5zHDMay8i9t8
W5r+TvFfUYlC3z8DhrBTmDlJlC0QAEr8OhbXqqwhjbyiWDEjRfXjGzyPfM660VM0hWYSEua5VG18
D/gDRtb0ptvmFZw9wl8Ab/pm3PQJ2nIdrTVmHt2H8oj3ji5qCeOmAqdmLlIhPhLQm/5gW+lz7a46
rSh0rhfQZ/cEGqFe58P03IRfWcSRO+aBrgR2x95OgfGsgjuFayU5axcfbcBvhmc8Kh01buMzFONb
tAiz47D+sMHRweuGHvmBzF75rhCBDjU2NRMFm+8cvV+ic4GvxNyiRT2r5A1excXRjKRjrZtU/N0Z
aRhFUrl006AO8HY7WuTf/xvx76GeBZpjpScdH+g+HMLPrS/R9JaPSZuM3pUNMg25a/aUYKVIL60E
W4gIvDsfArdl+XhE0IS2O7cQPqL4KNBcgHU0yKcoZaH1CWPmQji8NaDtf99ebg64bTBpyAeOZYu/
k0v1NErXDfzeLPCSWS1RSOymRAMwvjiWNtsx2+HoZ34FZoIFw7TC+Ym3STzlx8Mc/yNCS4D4RjlU
84+t8cKrQqUlOWBK/FAEZAY6048KhIDUcjb7+jTfW5HtpXNrR+R0QhlurVWKayN7JmT6KmGwE+zC
YX+MxBAjvLUZdlKzw+RqUuGrHXDbLURRgpbejct8IV62Wgp/6UKi7zv3NRLousgsdaZeOf8Zxw4M
FXWb33wwpl9nAiVrf0Eq9bvQPnbp6XmKqNPfXGdAPJfnuEeKIvdiEPh5TZlgORap98JXJVI7a9NU
5jT1ULufSJyyfCndEmUD6YZVKCEIAVuzUnynvV32L2LpedfB/mJ/lH1IVHlYQ38yhwa0KAH6DE3B
/Flv9LQ4s5odv/Wx+2jkERfziS8C2OVP9aPOYF+3DXjLCupOex61N6qpm6wiam+LFQLzOTVAnRg3
0O7Ph8ma42UkZDKIZU7QIYtBl1qznCRUtbCatpVr6/H+E9qFwcQRkK/zzrRxXzm1Z4rS/IXJgFEi
MTBdrYY7+ih+6UN9KSLEvZLedz7Jr/G6iO605mlXcevTNatRGVQaPPrah+YydEC13kScWNSeGFck
TZuziNAX0LcA8kQbU2PDfSoFBd4kZvXRsDjP0eUVFy5Mju/2GKmntWRbBNJ2DE/Z0RNNAbYU7DHS
4HktQHntU38VLjzHIU6USxUhX+vatteXSJ58l4/vWSMQsGQU0ekzub1Mmr+JIBPmEDXrW2Pr5cRu
mEQ+r/Ka1J9PsVNFvd9SVJCgd1xQK7rCh34hSfxFHd0vV0UmtlYPo78+n8vUEj37vq0dfO51wWLz
xY5t2KmtS/oeLYTHkZJBkbTpIzZe7UUxBDjPkBdNsDVppl5BMoIAUeN6kQmyKz4sXJ/Fgc3QIi2m
Nie75tPAsb7GlR7sznWKxc1Uia7o+d9ghrs+AU+15EaumhxnAOLCv3Kes/pXsu2ozOGT4J+AUo9/
nirQYLmCnMNH8Lrs8XYqxD+VOeYg5IDXpLwCALR1jdlgxJ2q4InrlToSZWzfsU9i+JuNz/UWf9oe
4sbZp9NkOTrc6tq2B/9XNyHqgZmeQGdgZ7FFnyElX9oLsm+cFNZ3r2jmRB14QwcuYnNJhhdiJKnQ
xTv1t4eOk8y5X0jZR485nj8fC72Bp2FP+xaM3e03/WayElAgXsBAOqNsIuyEtX7wC43Iqhv41ARb
7FMHul+e9rgupFEj36Y8awgiRED/nbedjbjX9xkFVNTK79in35LSJV6GWLsCi/VV0iPzr0y6CRHw
QNbZC1oTxU7ifDLSMgr0JzFb/RbNOrRC/Hbq/o3PNCq+29rXTQSKhEMHxpn+yO+1Xs2iby423NAQ
6Twtq+0XOPnOifwzD51af+rjqsb6c0E8Tg2mgvrBu8UCZeJoDakIjjUgjrz4DWv4HXfmctFsoM8h
/Ij/15o+6eba5UwIAjqI6fR7AF/HU8/re0C3ESzttJ8JAhPvudBHqtKLNV9Uhrsx1OwLF70aP4fX
dt/uo9rflL3A2f+rayDkTSNetdcJwUTkZkzzyDBFPUydDDFhnxNmJQO7Sqnj+Pdw6tp+ypzvgck3
52P7NtpEommdWFN4lMZ/UMrktXasSx5QaQ5SNbdfaGDqQ1gNTyAKd8Rg/qyIIWD/d6xRRL6M132b
PjeV0y8EDtrLf8kwITP+SclQHkjMb9zzJE+wBCFav73G2wEUyXhRpSEvl3GO78pQX1pnWgvUXFMc
kgntb1n4nwVv5LDtsAvMy/eRq7ILeb+rFxy6P+iJPWBEcs+VyiCb3ju41b/1Kdq93pxyciFrbtBF
Sd9fVoD6tnYdwkbfEGUlNczTGFI4f1sLaouM5cDu7EhqXijwztrwIXhiymJiA+lPLJ47To23FSpM
l5TWTaYMDrO61oppO328Ln/WNeRP+mJpEBJuaqzrxIyWdszWPQp48yd8V3jNJrjGsui0m8Vv0QsA
ObMKjQeEmUB2kdEQhE0tbGyubWaqKacSUwfWlFyvlFT7zD5S0WNbXl9VRzYPo6kC8dRrXtRBrbVc
wiyoQEQcneTQF4JS0JYlSube5wo23cHg7LcipFs2tHUl/T90W1FlT0MKFri8HQNYTuB9jeItbpU0
K/7T+Dw0k+fzWl9YoNDFsTGP+P63wJC/en8hnY2nXBy1195x7Ze3jacyI0PhOCIww/mtM2fSSLjS
puRvc+jRAVbg4oY8XQr8+rBxyKhjenh+TN9DEMCqVHkQdfvpIrnz6Id+dnMKJQ0vl/pVJ3UEYqyw
1kiCpOnwj9dK0lOv8aSoGn5hRH5D1cWh4Ajoy7oZHfJMmziKNXCPKAO428XpMb8aKjqObtpWPDof
/bmxLcGc73ootjiyRAoCBV8TAUN6zlKmfrDQdB+l6UoF16DELxJlYNmKR9q768FUIybXg2kQ9y00
cnwJ/XTzaVlmTHTIIgcawSncQ9dVOZnPf0CZcl3B4vxkNL9rr9HlKm51p7IPLUkY64Z2iwZHlKx0
/4hs+RjT5MRBgREW5BwTKupumsEhlwqZJ7StIM8+2q1uWrXZaYlMBIGSu5ptu3REk3ifqjO5kW6v
w9JAEd4tymC6qNrIC5GEkHIve5LQGo2FWoaLjZs/KDPtzeQdyGDMPzuEGfzCgjQ2Am/pcS8fz4zG
134Xi3NiKqvRkEXndZkPH1O97WqC0iTpSszyi8gIED7YaQVBef9i3ksl9rQXAj0LqPUsH/vBSOj+
Qw48gLRC208u9fCTgkXbamzu45kPdKI5TaMQPmRb6iIYF9TzrDudIGjNvgRp5ycj9Jd6tdveKCVi
1SLVctmTWkt5Lv5bD8mNXYO90rR6/Ld+/6wl3y2pTPoTmFLpYiRA0H93Ustr8eD7R1HX7uUWl1is
GedoTh8LygUFz6o/Av/cSV6pqayRNFK47zW2tzIWQtA6wfaRsgJkjEVgY19kwZ31IkH9kiMQVFzA
ZBWN+i8RaxAGa3hYqhHnGj9MB7lHKOrT8BpcI7kvVyN7T+npAqVu7a9L+wjkPvgcbukgVHAXdzx2
enTjfLULWgTsBEHLlno9/7QbSVHmvL55TZ8W5jbaSIDYwlAExu2RyyUusOGslrbXt38CL/bCw9Q3
L57p3uoZjNlVmeNtHqFMNPT3yVgBr8TNihNSEO8oBKGy0PQPrHPhHvlPq4Y+6Q+Sbw/77FDikq/l
zx12W4FquakppDgn+xDaESXaB32Q2tVkiKVSY+Yo56P+OvV6pY4oPAUZWJ7Ydjc/v79kVB0h8xew
uaS9ENpJVttPmz7TxnzPP+pZBemtJQGXRbkd0Hb5CUlfz2/dgQCTfM6vRaqMUbwdphqmAiZw499G
WgzVh2+SrB+lhEzYn7sYaJLDdFuUp0MKfmO/kLVEhTqgJGDH5/Dk2esk0WipePXgcW/+JAh+v5oo
jCUdnIqvFbXpgna3vTkVhG50aVeN2H+ShhojLxhOX8ZlHBYjAmh2h/wVigtqWkrm7+/xIWH+MajX
+23o2Kqe+f2bUlAsuT5/IZiVIaAc4wBhBlQLEcqh3l8HI75Bt7+bRJ1kY002JAc/DAlNfnYKxk5V
BNyc7MxEAhEqk+EAJx7mvqYhHCsZowgzx9KHxcWndaqs5+JhhtG6pgMZfDQYbhCqMvxag4dzM/nd
x3h030JTRJp+7FgRy/qNMxGgdRQUZv5jSzSf6PF4G67T6rbXSznzplAnYntA5lfUkWRnf/hQhiNM
n46Fv6qq52SYLwEfMgsgMbcIHXRGY6nAteSUz6t4z/+kj2jCwfmNYTiHh85lcXDt4BS0lvxHfXI8
ENWYSXNruXi5MBatccksjHcxQqAoCgEFR08TVawWLNesS/eer6pSKTEuXN4LQsGJnKPf5WvvKA6O
5DhdCH/n09MNdwix7jM/cLYRDdyf1Zb3y419T0JdXewkcnOOPdlDR9QSqDYOiyKTyx2XY0zHCVws
YbUyN03pcyyNS9Mwoverqv+6npdyP8HuuwvLY+Go3qhq4DMXxlLEOH6WwUec9eyTpUreJN4C5QBR
7QLvRfPfQLWE48WK496hQjMGjjSgcOS2pu9rSpSvDl+shQC+AUCiFHAIPUaWp2KCZno9Le/cdYtR
qmJymZvSuD5xxNE7x3L31ubP/Frr9hlJFazRPhU3wxU1zYV3JKWa46t9mgHb402vi55CL8cpN9OE
vhbTrF5NCULknPE9RCSF+7yuCK9jZ4W3ODfPWRRlI4cSCJ+c7xmWfKbzAKiOMuYM5Gpean59H4/S
96nUE369+4+lqb8gSmcEcsGGktyEAcDpTn/pEKS6y+a6I+1e+JiQw+MS7JzM8a7TX7ajkraFJ764
qUVnmvnsGcfMwyqg11VjtlRqYyo0gSzTiPNIJrm6jmqLD1RIBn1N+bG1kxosbh5f9R/aZPZA2oTf
vt7cEpKmcF9gvdMPpZasHa5CwnUZdccC2xa9e9qQTj/FGk1IDu8+k/jR6kHPilWe2qJ2Ou31uV24
/GOw/wKEcqMOoYSojgKcYiIhpOoZtRTFn1a22JlTS+JfMQfkqtJQFQTIAHDjul83Jk5l55hddF8N
CWv2J70iirLB22LpDDeSy8upHwf97jbKocl6wsvS/B3GVUQP/+1LoPTdIq5BnWSrgUoUJkByb+nI
LVAFMtvF7MOLPHUZpm4c5OYEVpVZDi9gMQGpuJJS0haK7e20HUe/375t46D+ZtyQxkCm8+n0fp9A
udxgxYkpvzgeVUIvxQBY/2XvZ9pM9tvSePZM1uOZhYaNJjaalSMM9bWdwG/aPQ67v+T3vss4CN57
spxvgrQgcbyeZ7KTne+IKVdkN72TLRnZngXoCB+4ZAWy0xFQrWb5GCUxyG/dXGUeOiz8lQzQlWXP
QqsALGpaYQrOlQ2laMuQ+3b7eUijVHB4Re0d7Ux9WtBKoG3nRcuoprgV6nSYWtppQJKeubWVszwu
r4CYUM/CIXZB7fgxBlxu/nJYyg+LCOOlIn5X3CXCu7iz+KUup0bJ5z8qMscjwDdPe5hgQQU72gjM
7k6vPyBSzC6vm2NtqGJy+INqFdvkNOHAs0DvehshjkXtwMdlmiB66+A5ssuKEANab7PtYddZ1UPA
C1WpDHsCe3EWtrcK4+daRpvJ0IFzjDVusAtaicjIqsB4TXijv8TdvgKrJ145+wTzwHbBDcYEZFgl
kl80obYQEOoWAe/KlosqQWriRwewD1ABSIXCeXd5DmIWrOQ8+Hs2AhNRI/8zMm68qMQ+UzYAlb/b
2qb3Mi1to30bbTWfKI+hgLanf/Jhc6E8U5VqXqZs6sDY7ISmXIHyeTC8GFTq5m8htgy0VFvhrnKd
dadhrQZJ29+hlXKJIihCJU4RRKyUcPPKmkCj+WNOndw/Y5xM8Czcs7H3yvwzQC+n33FoHg7Yjp3Z
2PQ4ytK4CwM7Wem0bdOiM/eafFuMItAPj83ZpgHZCY/SqNhB16MvlQ7xSXAvHnQ3i6abzdZpAJRI
c4oLSYK0ACyX1H7P6Bcq8bcZTYF4TZZADe7D9BhyEwfF8QpK1/MB+PFMYsVOoX4v76SYQvi+Esho
QvocBNe3TPL+H/oORMLxtsGlzXslH0o0CF3brv4hPHGL42ceYCC8Znarf1PggmWL8HpWmtiKsC/F
msgJ4tmpR3VGKuIXUkwbX88OF286uYjJoMjh+SfMa8l0VLjJXQts7JlGUxvK07UvN8R5pxHlDwAK
RMRdjiA+C6YDUM1/OTafDconye3XfTGt2+dkqdl1bTrhzk/SUsutM4HUBq7o3O5kuTIBI8CCLkeh
/vOxrpHbao/lt8kPV+YoizyZgRFewK9/Fek2UE2tAAk2W8He/o7ONrjT36/PVl+kKtlhhZxdWySR
7kSmTwuQnnDA9I9uHays8coKENniFACxzk8bU/6LjRPB1/0xl/nnngOzqGefs4B6+aJp7iOP19Ax
bDDYlElP6hKGHhygAxwdBi8nliGw55lsTo65qCpkO6X7Ziup63wHvZz68JhFLynHevM8h34krLOt
Uzp2UOxaJduXJCfK99ZPMn0FEyulYsUJytn5VH9bd/WhfnkC6lCXTQZm7mGrv6ksmPz2xVBnCd0z
gT41oZxK7t1mf1hpZ7oiZQxM9Hl27CEk+3b8sUGPX9UE8r1VBzJOKa7S6mU9sXG7nzT/IyGDn1IV
8XBqoF9Sw9KZtg2EWh2UEryeqUqb3d7jlywEm6qmAuD553aJI6uZoB3QQdq0Mi7TDA27zLFWAayj
3+1kgYz8pY5zr4phPJ3RofP8sCQc8PheDUQUQzSka5nQCf/dJ/aEfY7Jik15/tMCUNL1Gt5gSYff
HyGqllW8fQSdLRQZWqbPy2yHnnT0tzfatu06v0R1FAc03M0LfO5zbikJHyOx1fvPMsAknYYnC7KP
OYJ+xo2WJoytDz/l0zxWT/QpxVsvSLi3EhusJ1Tkw6aKsca+Y1MeJ308HppYaK/ILW67aawfgAGL
ybaam48K5DnnqYd1WMRI60mj8HxRXAyI45iqE2KjQCjDa9pcklLEPsv5bCBGnM/HPSKFWbx6spkr
M06Pe5ElLiOhgLSR+ljY36vfixcLnj1JYpgXZQoIgT886USMgJEq5Y3F9Hk8P7B2f3yoPN663ZDk
glNF9K/kcKZexxAm+BBZBgL4UXowZZZ4hkIv36Of5RnRbA7mbJ+qja0TFGIFXVrmQH3qBODISBti
har6TUAdk+0yq1Vy4Q03hq9JqgktJ4MVRUpJd0OcO3wMEinU/mjDXPdytxmBvhWmgeDB5k8p2/R+
8Qr/G/3JOMo6jcHwhKrZnuhsq+cc/5FOL3hkeQ2CvaHBEwdWFu6Jq5D3RyUs7D0IzUQST6XR6P0x
kFkyvT24sksXiWN9O4r/g43SVMAQ/J4KR0w155IqfbjGCWmMTqekPc+3xChEEzlkmgM/FKF9Q+Hw
8WcEXdqFifOuXYJhv1b0DdzDrjeoDkPJheq6uZiIN7vvnpRdZ/ho5wtLbqmnw3h8ytNo9+EXCQbl
VUu6q4Kxemw2SkrICPncDnxOBPkUooeCCeKyU2nea7OMtqQ5+FoOPs7Hh3a88DNtDNeBdvUwRngq
y2aLIFxV5tsFlKYNvLq94vWHtCIpMn2atWTMm1Q4eezcXRxe3NFdcYNxf5U/n1QOkKT7jTEXD+sX
jx/KKEb5xap19/J+6TMjGiazfDq53DjR2Fb4LBlzZFRpqDWooK3n4VDR3yhTGOrQxdkFtKWwN8mA
7oid5enBIkR3MKyC57tAfcf79JR5rnJD+QtgBkjBdgu3Oe5WUyPgbF5FuQz8a2ZHwdqQhpQeqhVt
e/tZu/LplmeG9Me+AVOWDKwl0EI0y7OloZraUYoeTYyFYGNJfU5dYb9PH/Db5eumkau2BvPOVQn/
nnzUWGW8ZgvL5q1J6OsYvy5i82z7gshaYzz+XdM/MqzjemPFAIMC/vbc5g7JThgPeArQPVsL7art
UzThqQBEQKkIG4ff/9+WwIIim47ts2u4qjFQpSWEnGQ1Yf86Us9Pe4HSDjnrjmumVgwPdA0r2UGM
PxLxEAIIzmmjDNIzzXsHL+J/KRDf1dMVbvk+bPp55YIdBHDTDGDT5+nRDzzzhq4yHgSoPFjGy3jg
Luxm3vnqoIouorZczfjvTF1fzh6frYP9+Cszavx1Yll41sgFTZTVHm6vQ1gLev34DnA2AQ3I1YIM
8kChP7JYhB6yp5zwjJKhWNP7NixORn/uCkFqcpvxFu58rCFmwpKZ39khn75IXsFNq0g+7K1B6p0s
YDt1yAWQPoywwVPi0YuecFCABfqrAvkDFHa4pEGqpcKmZeZFPTqrEHg3GHYyMZAqzi87O6OGY5RE
QFsu/Og/N8sSvAUaIuVZDRkYU7hAqj5h6X8877QXO6Ct8x34jS+q5xrjh2/ESy9jHLnQK5KXcSVr
5clQ3dZsW1z/cSQZBAcTpPriBt1+GkUBZEfo/lCO7rLqXonImPJDe5nZT60GpzJmNUFZv95/v/9K
H8kBgVrBhVz+SS5DIi4FyXK/M0MuKZHs6jZWFo54egTfm177XFXJkQmlxrJCJJN9PqBALNbttv4N
CGo1xMFpPXIJ6Kdcbtvrl/yJZl9sNxCNqSSlK+S//Q9EGrFM1krIELzlcFNl012sk32sJ4mFgxSV
sjG9CWobGe6O+REyBP/nP4hFrbk6v7eqglo1JervYWRfKEbWJ0FQla+tDLNpl3udD0ZUaXs8Q5aD
KDaZrr+8rRfhtq6xLIb7UeVP2WCANV8/VGMVhNy0oUaY5PCCeQnF5oawFTMJ7DGF8OSQuoBdYyIn
jP+gJf+admtCQoO899GO4Cg9oSyEqXCeyi3GF1mrk8BI3of1GwJyY5HLcX6VAdrWzdAlYcerC426
lKVFR/g9MC6kUZQhRLqc3aEgh43LY9lAFZFWqqffjArkS1lfcHtPLC5A0gi1fkWCOV9Asyitdrrv
XtsC/HS14bCdpJunGxMTlIxkBK1n87zzoMup0F+ZZHCQlaLaYiEHlGboD3rABcij4IpmRgj2xKI5
uS3Sxf6Pn9U5K59wokSSu5wPc3FmiMUzvaBDYEgd1i+USzGBv16PDoUZYDfVrNWbD0M1trPEhwUg
muYpguY9fLhyPwOyUWp9G/iNsepV85hKo8ygjt/yXTo/LNrSTlpgTrCbzPtQHjDMvqg+15wgdIZE
QKZK7ntwak4CUSZ3iOREUuKjoIq18/YAQsVMt6LedSX0V4927r+hdC9NWj12xU+sakjnZ6cueG4N
MWIR8y4ksfmgntybc8hK4Ie2SPAXrtu4EKMrC974aXBGowqKQi7WKBQzNWiSmAstN22+SLA7xB46
svtK4C1D6rozxuh8AZErZPIYTadf+L1VSD9rwrToBVyXN7XNLqAgiHpbJOijm/qzyMNi8y91/W80
mllqNnmjBO7N3o2jodrGOOAR8qJlLDRd6JuFjQwkqFBSR+OMRbslcfKjttcmdFpY2PND8g5QGt+M
dfdPOLT9PXz46vxVKJVPRYFVOdflBLSPQ2oOtDZf7W3d9l+LDllocYrcz7lszcZEuUHGiWGt9XFx
xfLwaoIIfM/tB2xfpe4EKB6KiNg/ccs8KgkdcblPncLskEw05aWo9DngbaRT2sq5+c1xaPfAcRQ/
o577UCQX0s/2NGJ0M8x4U7dShfOzXFIRcvzs3WuOlpQGkqyrF04+NP2Q3lXXvDvzVY3rWNJ6CSgE
MmuwVlpFzgsnAtg4gfqbYXS0UdtQGmDFWFJnx9AQ3ED5587ZVD7M2jBTNdwniYjMog7sLke2eoyU
GsmxR4cKhjpG/pjr9MHODAT52OtfJtC/yqqelirgGMx5V9EHLg4lw1w2BrquMcfBqCVUUkk47o3d
m2P/h2SOpd9m0W3PtCTAz9MD8IQWIoK4y/VKXo5rjxxOO6t7fxg+GHLykawH3P1tYHR2TWvpp+O/
HfRy5nH1Pg5zWkAqrFWvs0/RDGzgB+mmU1FK1LpOAoQyaObSHKTxNixhlIsBqmIG5xRKcJAhVpqK
dGBcoCcIJDlXHYH3d8tdEkU7f9CdKod69MxiX1duwZ1fXQf6uI6PM2f9JTzRWosKMJJoS+AxTrke
ZP6/dFXMo0YAhNBnTvEjcxjkxM+UVpvdXR18pwJRZUbzJXUdgS03jxDCs8kmrzRgX+AWkbFrO9pk
BrgmM+9A/KXkVbPXWH54vSKAChKZvPufxmZC8zovG5RGMlmIBWMhl88ggtJ16f9RmxCH74etzJZ4
XaLaZx99gz4TXbGqqVcCY3raviAbRxDCHkTh6D+ehRII3cb8y/M75ZH7cXcxDdJ6WZrtwaxh/mHU
Pw8ZG3UysplMC1/zyBZvexVdHIMfbm0EAfTX66aTUoYspmHZbs0d9Mc3GlX8Zn1iV6gcPnCjr6a7
CRv7PH+guUZD7VlgxnUpmybx/BOnQBhctxLZ93QOWxY4j8UxI85AGYNMzzXXMzdi2FSfLaGNZNcM
xNFXY6mUCAMwLJvXFvCmqcmVYkRotTcBdjQxycjv+BkTcukHSCY4W+OCpM1BFMnHxBF4LNnsW3g5
eVbM3wqM1I0WWj3F//KhV58laCtJPgE2yzDHqplvqpYkL9ay73gykgnR+H/FYDJiOwiKUQ6WQbNy
lwOFsmIxJE8a3487q8mFOPzMD2AXBbyBofpD9F8mZbMxR7LL0wdzQewN6+TQzPd67FH844MwiMuA
3qngksVgqva0ANDzIKHw7t0ea9kzlIGelOXCCDgUfZfTrhYAIhwouBHks/2Xp4u6cPK1qFF7jFZL
mKio0GOqPtJJg/FMaPz16JDRUAQupwGryD3Qicm05ECHjiwZk8bBAQ+Ywd7K9b9j8wg2ug9ysCie
XLsM2RT4DGv+ixzH1WVAQqy/1PqCsD4dIl77EWC8xUVxWP2eDpAlsJVE9k7WQL1yYhH8pMqWteVp
/g5HSwG6O9wH3WE0GE2aQK2+WD+h674/+3bjiXi0DpaNt7PNkb7GyCb9NsmbRSLQ6uZyrrEoQKyP
BlJ0PhwcifnQUmCZ3AHePYyoC198mgwrrEEGwg2Y4ZCt6oClew+PnIPkCcrZx2kPBLEy2Yesuz3m
EREg5/Odez0HVrrA9wob6feJ0uxvK3UZqsVZd/7yaoQzxBEqjYHfa0XO7OM/fvki1SN8W6xk1YG9
C9Z4FNaxz/AmRGXc8SnHT58bQ3vzsw8slk6krsWzCJezPn79H7YlJnbSvcbZgwH2WYKHhb4CCxkH
9In6OZ3Rr98ltAvZmS2+VeleZGNP0AQ2QD3mEhUsN9bO5yjp5+1pNS7rqhQeIh4eRk9H+9JV0soC
AKwHe4tcL2+3I5LTIbdxiFCa/h2NdBGyjdlYrtjZ4QjTz2iqW5pW0g0i2bgb8vJIw2zVRBKM/aGM
oFgOLYR2BNS4d3TZJgTQzpKaJ4MryDjJ5MMXuki5qO5cwwH1xfOyS3swljAx70DP9m9Vj/usJo4P
FBKY502iULHNKd3i+C6S3CHKCkbkfISJh9Rb3UML7sJ1/7w7UzhhKPb2RgIezCpY66tsSXqWIxTT
rpAHtM3pCU+huRVDB0X29pft7r4tmVxjYcw6JYBYU6bk2rg/iUzR/lU0izM5bGJ/dtdoILYqF3WR
pkXYGM62nzUGdNLuFN3Fa3RJZYBKimjfirIMkLMcf1HxAAOlbZwbCfbJxJfG6Ceij1HSHaTYoo6k
MEybt+JJ4G95MbL9sXX/pdt6CsrLYQMLdnWYZ3rVG/Hdx2VqPKJ3RfZPOtlz5w6PT+prcmgF03g3
8WJ4y/4p5X9OUS0GxOaoFR2yx5LE9dDHGwR+HjFrS7KYkXSmzvDvzrxYtUDSvjvXDCiQmw/Qw4ix
3WYrLFJtp11g7VT3CDQCzFpsJU8teT/Q/+bWRg3n1YseAU6AGWGQHffzwFbZflHq/rArBCz7OGpI
lkkHozFmGMFNvmbMawWxDV9W1PrIr7yXKjbjbrtu4GNXQJo1Mj328HZTxbllGLOpnOUtr5NyzSQ5
EeONRzh67U21JcZO6h80ZFNb7JhqV/CMi35UGoLEe7fNjdyJw6LhXrzQSKFQL+8UXeSZydtWhOT6
Hudt64cFr+nMF2qzhxJ+3bx4v97eJibc2aXrt36lvEmPCq9wtFAowq/Y4KYmQUb6FCvCfzpGLkdG
/d/yur0XKlTw/AC0LVjOA+r6RohigphVee9bRuseIAvQh7f582qSIzYa7ZJzuHIizoUd2Kth91xj
3MPZ3HTAqNqIIikwxrSbLQJXnoXzLBXX9gcZMrhiW+YNIKc32N0Xf4k/os2O/mRWy91gVHpeXCpF
V6voSi8uUojaq6kn0seefVa7WCfPB54LpiwcstvV0u8oLaGq3iC082B/YzgGRYDsyu/2yoj8aIO/
9AY1sU4MK4zAKTlWvdZMnEh4Vn8ddN4I9S3aFfp3y0nci5D/ULLJhB+LMIOtMm9ZPzXUt94V82ls
OrI1/aZuxOKLpGwwmjw7YBg0AS9UUK4hRC2VOhN1BGP2fIfMrhMcmDXVNiJOv96fN2q4gVUqH0/U
d7SJqIt/UsaxKA8F/QEf8HlJVK6zQySAwrjBMgaVswgkjRkNlOUuxH2si3hTPuOyTXf28HGNjyFS
9FkCiXohhCF/m1RgYYv8zbDr4J9eK0DA618Xsxa8nVQ9cSSsfREVezkTXljkuSe8PORHXxnHX69l
XvLePRMA8KRR/QMbYqe8Rw5ccnGUoLLi6hcBy8Us7bYORHVjlRNQ8+mNd88omVIag03EOgwB+ptT
eJ6Cq5HMAmbEjRLBTz/ryEy9F/HI4FZNIzTfDiqfMALQKRkQUkNR0iO+Ir/WR/tFEb/xfe2EQ1P+
dirslf65Y+76nIMRS98aV7Ueew6VGVCXuOf5zyG7aL4Cb374GkhFoJYUruwHTaPqoqZXRRZcL+z9
c41XmQzuAZBx2iA1xh6MU8R43pjcmaJKiWUojzbgZBTGpoXcib1wH4ZD180KhyUgVLtjqxjt7HLV
9MOHy+qrK+h/D5ZMe+qvF+zAqIJm80uqdA3tJasYtqqur8IlEEgJ04y6kgkqDGoSQjRljWbiHUlx
sWr9TnJ2Kuk6B4XB1oeJFimgPNQ3njDuA6HIirKlZmlRfhUWCC8UTkvFGztyYWHlRSdf6/1Eh2oE
/LzRYSCTReBJYV2AzfgiHwI9iEtl3PGWRa7NTlS35SxHE8GQI0zOmL48KOWUrsOTNBT08W9Ahynq
6dBnA7xeD99ho+UrhO25YEmgrj2zo4VStLBWo+w9lEdDHNh/bxFXf+I32TSyWLoBOfZ5JWmYEJ+8
c/RfxMW+STb4MC8Ej5OKUV805VtYvFykog2y72uE9fBvQOyUXJby+ayvX290rhJuVKkT0F76pov6
BDtHEyp14au6LJvB5C9+S70KIhE243jm8PUeepgGfiRP2wblixSdXRecex4md0nthL05SZMkDwYr
7IwSkNStQ8glMA0NimmvKJB2iIjrpMHUXxBUxV1qoSrhizPo/8S18o4BzBAdTSI/AxkMTbOPupXJ
dLgfJFbQfh+1Are2Xcoz730b1uqEc6cPm5h5UQvc1SoeS6cL4dHozqhITxZiPCVDR87nkIwmq7ec
PqDekrrDoKYH81JAU/LlfYYubP+Q6jE8h3SllkoLrLm4a3XAfN/UaTEUYdfoum0K7Iu4HL7YVMPE
8/owkorVfSFqLNk+Y3Xn1zDs0x5fDHfYSEE/7/6sSx8S1p+HZJIOiiM37fqUPh2Hbs0/sKRtwZgR
UFWdwWPkA/dPlgSu5ElByPKpn3PFCV454FjbCDw+ftqkvEL0mUjM7hnXPR5yfdoiL1sBJbl7res4
C0tm0XRg8mKAMEE0NxKFEjU8rQi3uL+qvrZsbDbAgPCFQyaOWoyGFdG5ArS/eYFjsgV6sd+RvZTu
vGwEz7NPXLNjtVTQZXXPK8GvtmN6l222qiu9p+Liyn5YeoMCmOjgbN+0iIEn/rkTzkYVN5m0Vlfd
xLay1xuIdKJgPwkawdFn/d3FTDTNEE3KuLSEgPQD657UpVD0ZwX4oAY3kUL4WBLjVm3SOk+/pV5r
DfsaJAV83BdkLTyvKH3ILy2a8T6DL4z1sIOKZ0JXhb2cs1dBAtyRpon0JVGlyM9i8zpRlnbcA5fc
j2AKYQIz5CRfvHqGKZKWKgwR7rkN28jDUN8Anr1ez2/Q6JvkkAtUcFnK2ZydukP5Dz2MBdCYbq2K
Q23rLRcOLFHnaLZM3sLNHzsqFrvrEjbF4gtX31YpWfGJaki0v1nRoIqhmqr75hLtUL0TGyUpuGzf
qASknIE2+o5eX0ueLdnWvIcoTOTa1SHWnT/lz3o4c0JRgv4tmxEfCHbmLI4AxoiUKC6++9waB4Ws
WevVAKONSURETSR9IvtuV37h2cmQ/njD2rQQSAOiWqIBo8YKW2FhG2AshdXiYqdH0SSAhGvf3QX8
lN4f4z7gL2qO7DorU+M3UDC05I8NwxpsJQlJUgvFFGZlA/kUxn+YTO835a2G+Jn8uLAurGSj59dE
/IJoyOLtT9zZcHbtnH5SfdgcYk0VXXpBn4cKl3mdZULzaTegLsU8gK/FmYQBV8+HL3DlvHksC3Fj
APA0Hvu4RjSfksoOsVhXBAKKx5qEYHXDmi+y4en9o1c8/62xF//ZuHAH+dqfZc/4nxjrhpAPReIV
XDCMdcFWKuO09wKrHXbrjx5xXhrXpcAAin3+CezLaAuIablJhVz+cag+gKH1wlUkYmckUJ2ZzIvU
zP93zpBKsERaC4OdNtC9q0EjSj4Foam2hI0UdtanJtu4QQYuIaogxsw49RbInLqYtdPy9016rEPY
viWjn8daEN7f3eathgaJVZnplyl23dW+vAX6h3o0x8qAy8/0oh3cZ1ICFF54IyVWyXpw2HsMboIf
tCxM/M6J4OlvkzLBlm7zpsH7r7vpanWNyLmeEBMr2KK/i3RSij7/O8sbx2/zK0dV01bJa3nswCD0
SPr4gnA8RqngyFWkDbtyNpcOTj7rixaJHjMyt6hoSC2b+B0fuMdyBUFjlD3DT7AvspRAU6LMQIhD
6gvw4rk8vebDz2nQdRSND0km2l1bqNenWA/u+JidF31W7ipI5F2KUT1Cvmi06i59b4WtK0wMTe3U
yasoOuJu0XloaUHKmYDilCviDuHN50PQCkqP2uUaxzO4ArKubP8uEZV1DlL1k1yK7RABJV1t+co5
sRUigNGMzntIY4/k7tV082bxLEnT1Gol6XKTmqqUrC3rKg8ZyTHv/z1YB5R6IMwnJffV8e1hByhZ
XI1Re2GroOYInjzxUlaQsEnR6HyoUWed+nPtnOGs4WAmPRQ6nSXhQ8+uqb0UauQta7V76+0Xfj36
CN160/y3JyEwCiMsAhfcZxfwCoGW5weipN/hwx9vCgOsoSwuf+w/IKP9jR+MnaoMu5APmPnKlZ3a
5LaSl1lMxNGdEwCev9Kkg9MYx/dukDSWakdFKCQDuKjqeTtoEcJlRWYRr/Y7RdRiDePw6sMnpLRN
2AzFacQw15Om8I/Tw4fu7NI8ZmPlrGmiYWmm03ofoI2QsGCNVVSSfvUpiZ0EbME1zGlSLITv+6J/
jFevatE9leEqsmlHIsgELlrOqMMnp1uUU37eZoNZFldNUIXjzZQGWaWPAyq1tkMZ+0lpHgSEc3nk
dgWmFix2gIcE1mbFOiMJ5jxyavlIjsw5Edu93Bg855NTiVngxGD16h78zJXVhsNwwigXw6gKE3Go
2wrz0/v6nCALfJMxA3zaokukfWj9IR1SCSsPWvUQ8oUXlIHIdZvI/8w5LikrsZNXHPK4ZRuK4LQK
HbxWzUcs7yrWD72cOlNaf6kOecqByWbBtPOW6WAR6crHb7nLsl0CmAhszZu8wi6FZpeZglc+aq9c
3uPGkCJgu0x4bkKm1ScU3k3mxdMYVWk45WKMVIyJAk4r9B78ypeACTm+hL2+OgEarupx1o0G3nyD
RclNrfRJB4QhyCw7bP0U5//NHI3WUyVtN8/nPc5KuYbFjDyuqId+lz20m0TtPI9r1fTwVcNxIe5Q
swmrnjfSaJz5Zxj29qX5VZL+AOPOMay/FFAY3jQi3LF4OBtK9wMJO9RQjc59b99okhTeQAmc9XSC
ySYnc6Cs6tFCZf6zFOevQIhNY1nl3nNMNVJcFyGC6RiPomIS7ulyfaQvj3IvLvSumB065ndJ44mA
vRiQZ97fcnz2QSWKcH73rpw/54rxpIdYZoRISWcCR7L/x5iCwAF+2edt38Z6WVqO7TqQNB7AD7LX
fEibi+WHBN+zBGF9Uh6DmKjNTxVltMY4ImMQ7NwaO75AOAA94WgwR3POl9bgMcAm/NpEH26051GO
Bm3/CiU0R4cqVnOsQQ0oNqr2vjA2uSm29gOAj8D9/L7KzkzB7YZiJS4EFpE2K5XHEouvw175OkWv
eMRGf+l9iNSwnusH5UOOw6kWatr/airTahLe+YnAYWLFyXp657L0xDg7RyqCa54Y9kwkS2bn+c1T
3IvvJZrRdzyU1XuJV5KuF4v+X9g30coq/zxcDKAD0vTvTn9+KDO34JFuLUN4JiMGLN8fOTJs0ihg
Ml1p1ESwkhs0pTg+b/HIJrazxYMoD8bJgz2mecsIErHjDBLBAHoXUR3mGAhZdtEfjLgHKyZ1uoj+
wSJs9CWUUEYpdNlkeOJ9faPsjw6cUo8MoEJnKZXE97tnHob1L+Gf8pIaR2Tx4ErtM3KhITbDloNt
G++ixNEWjtkKwOukJCBrVFaO60k/CzKtBibyh0aepWH7JlRybOrU6idTJFgzRYbOmecsUIvXPJOI
gQDJK6SfYxdb8U7UIhLnWlgDwo39DycJVGYTB6tl0wwe9+agXId1fhL35ngb1f4MVs/87OeJKniL
ePbH4+Rny2Dgsq0lza8jj3+FSgIUpkDqi3Zblqmu1em9wcJuKkdDlE+Nm1Q4KATpFbg/fqupaaiO
PEClLnDt4Pc2c2M8VWBM1EtG8KTMyhw9kBqOi1r1rojaG128reN7m6MmPOxgW+iYw7mbiI8ApDP0
hGo9qoswFZVxbDq9xejLspQMihUICmTqCY5La+pDKtxT+mi2/CLI+Ou8IHD3zZ/FsxFpSNxFidlO
wdE1CYXjptqrtpeECy4uuCpwPFhrB+rSeLBdhWvjM21YW/7vFZizW+v/ev2QFU4tBuZVrm5ZrEZk
yFw258O3Elk+C2Ub7M4+0WdLC2LJBVa+oWgGS7Ee+JuLtx8Fm4gK21VhwoYYe7RJ4ZyzZRtEhAZ+
xJxKUMCgyN1/KPt98l9/DTfsEp8W90x4KrZ9vRT+G2pQi1lgjeRZFnC2kyq7kHFsbgqj4e2erzNn
Drmze/6lyzbyf0kuBVA0+FoYS6X6R2+yNY8bnPDhv7mptz3ie3R+CseexJGxQEOpNuiC3S2u1NBa
4r5CcWQq8hSxkOkPqT/DOkyitrtYS+1Os+byatuFunYvle10U8LKrER364vmaol+PUlI/GOzKoMg
CLBuYtb4+7WCXLElcHxuWHzDeLtQVOcdZ47GbbJqiHyicf61hukKey0ORmX/qqozR+ixmJ6CNvae
5HtVuB0NXzG0JiJsWwyDbl2G8mTkIrKG2F+WS5OsV8cwPSLgLbwfdocAECthgMGsFFjO2R5B3i2t
YCrVSHYajsLohRjyIGuU4Wivm48ruIKEuYPy/uB1LYGrMpMmzsWGXErP5KPQ4cHYiFZAol49zP/n
lAyH+e4soNgt4W4TCqFeSm9Hlaq2L/oTMa/LDoAAC9czFS0GiQA6wBaClsw7rdzVEAOo/OBr1ovd
GwfZJOp4JehVXFwkEK18rJzFqdTaApujqmjNyc1P90n/eh3t7m/kM49QFBq/wH+DmMh4UVNeOsC6
jQZu7LRb8UtfxUxX3XanppSGqXYNLUS+vZ1S0hsyCKuk/6UB2Xs9IcKetHxDic63eqL6ahgBooZv
OF6oP5pcLNn8C6pEEde+K7Xqkpgc329PnVmYWwUCgZc7BXHmSci+lLd3uS2YjEVmXImzadmAQKQN
gKfgShi2sD3uFrh5dMU67w9ZRPDlGQEpGHSJKQSXqDowLEqpt2ZaYl1Quhpn0aIX1ZuRt09Dvj9M
NsvqxveUdZSH85wHNwBohtyChqtK+13ICAYMikLQygMXmgCRaU2uMNdOqBDRvzwBmaBTWWdJAV1z
i/HorT3OqEkRwyooS01GtlZGuZwNQc7kkB6pNqJ45G4oOwCU+61yNaXUGEX/2ej4B0xbo54o0RgB
s7zMiMysUlT7FOMjZqS1rdqlJ0mfVHcia21fNBZ7jXoJorl07gLs53fPWjP9SKqKMAk3QvHP6pd7
2JHBAnv0VOWrUxoPLp77SZJOQd4dT7BYuDwKs3DwkTuuvh3MEH1okw7f/dr2y8S69tYWlCeCew1a
5DDXnUTJtZmh1n8CbpeF++OCnJXQmX61EeldsWDE5j555qAKrbhS/5P/JwZXT/mddW35xGf8ZcWu
KPrFEjkDA6iaBEHKlUb68f+U9TFxEIUwZTIMw8oZL5S/2Vcwe7eV0EL/I1M5tXmeTJpV3DaC+4xE
/1QJYAPgW+Nrz6zaB6mg9rFaoq2LoVxXMJFahCDKl8QT1RyGj4DA9yg25z15Ux7V3bH39MuliMe9
UiwBRGtQKZMTD8LbaOAG1I8qdvETPRKYpyF9NNO35lHMl5GG5zEzJwfs1goAsOmPUY6GdrQHsGKY
+d3SdsxBZIPmLhxlRBf1n6uJSF4KkGkuY+f544g7fmJsr8MWBSt1cpV42D+7v9mwm9I3OuVahHPi
lOlWX5NihQYxysTbqMoqni5vwb1zrx3kpA0URzRFecyu4Qp/677YL2gQwwGzEAItQEH/w+wUP+9+
ZSMAhzt4Bu/MnA/7Vu+WaZEKEsfjCfgoM9M/RXBXYQsvVwN6unfHp+Svwn6bCoIf9UoFXXC89Zjm
JVXxfxsD3lxJlBXlBgrbzo35AwjEE7+ONBv4uTNvfLySw7ONmFWbDYy3tXflXfZj9/akLShiiCE4
Irj9voeHPjsOmFaOmqW9l7DL2Et0vMilkXWc+VYmYqUTQZpKGN0MyNt1EUG2ECKWWa2zTSQGPVf7
U4oW4c5PaVj9GgVWhHniCeIADGspmIz18RBE22EhbH5N0p6COIVw0FP8vUDq6zNv/SdDY/5dpm4J
kr0us107ePT4dM3r2jRlIQEWjZAF2qOrcoNhoEHl7C4RBbYDuMiFw7ZFhOESRi57Aj95gLy7MXtC
FTsrDsx2TrLJFqLguU39v1jvfHckaO444fvfrhiRDy9O5zqy9TYtJaH+KhYZUkvFwuolFI/3un21
cLP6ax7kslRwMeK6ckH/wOffPM1go6aD6fPS3Go7Pp13bjx2TbYLgCzgYYpGMNuPr6PmGMCS3xjq
D6Ajja+Lp+Vl32Gg1CeKCYavk4oAxtpO5Cwmo7oQBTp5SaFgyvGNvW82a8E3nWfd5J6uTJOKUGaw
P6b7RX0TR0I6FzXbkwnGG2zEexEEHV2Mxm0Y+LJ/6y3i+B+peOpdSHRaZe84uXMgY8RQ6QfSV5BB
vC4SQDV+xaRxUkYKjX7eez0fXs3zgPSJjhBpJOotzYUIcX/6QanrM2Kq0o/4nUxsxIbXdX0Y7ZSk
mNN1Tohk62QXX80+Bc5/rAZQWv002lS0D7wb+RWWVPe42oAKCB4YAHfR3vdJ3NglOxPv1fcw8utZ
udhp5oC+Dtk6ToOagFtAqOdWGwy2pmKXKm0XwdeidGlRLG3CI+f9J1ge0oGTyRWJDdGIPI8zueeq
CfuVT/oTfYENYhsUTUzDGgIPb5Vi4n7Fu5odesgv6tBIHGEwG76XKNJK5RAVugYUGxw13iRmoxaM
T+Ptx1jEHj4Nwd0MkTJ9xdDM69O32COhziLeXY84K+NmY2/XUYsbgyKDd9iaiaEgPuM3fAyJzgM1
A8aU5VGu5NB2DhazkfwTf/lWfOf1MfI1vuT8DPj4TYKDqrB5/HF50b/2Xdy9kvi3dclScOxflsaq
1fHqeXQ7pK/LhFepXcAQMEdfhhn6hUzevKusEv9AhP5ZX/KcwqM479SaluZzNSUVURmS973OgOxO
/hZZZGzbKCMwxXe7ZtiSJFK3iOzDkhmXxJQTiScEn5GdAVyfZGW90Ib12lopIf17VzXYjH5Lod7o
L9T0z+Ubc05cYh98Y4maoy/hd0LETrPhH5+jR2Fwk0iuNUVOPNogdy6ZsS/e4BOblwssOB7VnwAP
LLOvnns02LXEdnbvOseLioCgMVxp/ka4WaebCPCgYNXff6JYS8FOFqKGWJnQiLVbVcKl57HsiVCX
jHUbq5r4q6fm8Ofo0JTt8LScHLnFF2wrlbi4UeHkQ9rU7UfxGB3oeVMDM09kjauz53gp0kDcJANs
KBUMAoQ7um2EnZmeENTnRnkaD8Uk2tsYUjGWmFj2e2bkao3N5/yjWXpv4MStWuXU0B+5ZEv20YX3
2sPg5E3RrEuOwYEdYGl+qySnp9Lj8VV2wUQeABb995UhA1GzgvxMPtoQEanEYpSEzj0zpy1VDEBM
l00lKkCFQR/CTxoSwUchKHps87AJWGUxXzvV09T7X4i26nqHE01DWGQlKwW51BTYSVls2hE3kx30
sSUjSg7b87uq66ZTCsxxVpZt38Z0/1zX1HA2FaCzG6mU/djcz1LTozhaWMJIMbBwDiguxbyB60j6
EfZnhg9lLZNPg/4wbHyj8kWpKmMcBi/Ti/FCZDimUQ0FdvtEv/3K9YVONo/uqEGk4kh5m3mVEboy
ED9T2Vcp2sNqoeKwaXatpFFuZ3VwzC6u/KB1fMKteAvWGbjCw1nRzbHlodGV3eyxzmhSrmE0XbEZ
nMcWXb0FyNvr9UV2/qABGowaHOyW1Yoy3DaRy2kxa4QTNMO1U/JnjPKea8YXCqneXgUp2d/6QndS
fSH5ZYMcxwK6+91cB1CYWvBM3J1PYSa8BUn+xbCaNWT5DVpwS4HCNkc+A6XUDWDGcOh+pZb0VNsT
D9GPKUoKY6ziKCk/+DJ+VSSh93SZqIGDn3hCkLdslG7yTr1tVs510aEeLoED7jOPhHlJkKKoNGwE
go1y8Nx/Yt0q0w7tL0/3EZaxQFyGxsp/ZSue0+IwlN8cUYXIzCkO2QAlUlKOZwrD8+pzwk4WMEZO
zaNBox/RNM5fttX2pCI3KD0Ia9oPv//+jdB/Re3PNgSAUCUiHGdhTuaQp+rF4o6flguFG9C50X05
dFbvP+FGk4nI38JIJiOPcYdJ3vDKorCaViwhtfuZdxXe/TIbayWYlYMf/y1033UldEiK1i3nTJyA
lUEkmOeX+yVX6Ptd3YSTxsQfjFhF7ZiSv5tdZmsPc8ylFfBwDpC+cBqOs7+xppL+ShGWJ3V9lz7B
/KKMRvJLtATQ+sxU24KTaQCp2N0Bt6bULMmAS9McJQ1qLUxUjJyvz9wht47m2X+Wvt9pdr4n02XE
EtSG5KOFvIXhzAxqpF2FwF9yyLqSKzUKyrUtBQkDYfyLTWa+Nc3H3hpjh4QJdd+86LB5zSR1Kb/j
NyCFsEJKqgJRSmigVRVCYd2rE2asw1d7W4p/q5xrGCATDEua1kqEE47n+MnAT4XMTATRbGOtsxus
GK41hA1sdjB5jUf/t8nlf0OqP83XpB4vo48BZuGjZXJpZhs9VOwUploK98YUA3ukvJIALdU/qtnU
gclJKZWmWebR+VyWnMl4uwmPzpDI1hDF/PLB2aSE6tVCYsTV72VAeM7HjPOSr1nMMCC3kf4lclD0
Jv3AcbxFTybpCRcW7j6TjewGKPC4Fjf8REwkRCrYE9dYX8Qrko/gaG8Y2uyeZ/fI4UUezd2/nnvf
qfp0gLnrE+3/V/MKRC7uOzvFhtKH4omBubUO1JZGQYw4WHSsool+STbrcPpJiOHCzYhOIkEKkrOc
UC+ZKXpdCY+wNRwQXTfASLodq5q8XfpvrHUqvTWx9MJBgs30XpJxvQv/SPkyoE7dBj2YYudxL2uL
0HrfVOPxhmFJUFyhfSoHw3SdQ/CQEGeINhlX9x+CWNn67iCArNcLOdxJKQZIYjI1rOBw8xhCOIVv
UnSOun8Oa83O2WSr79wg89Kv4WUlhM1Ox1jfzAvEzxqjLvfwEH1nWxI0ry23avGrQM1B7y/hd71i
0weV6sRiVjDOVIwSZJ7G6qe6jBVt3lwjtYl+RMFG6NyHQCzlWJxhf9rSbf1Ll199OoQtvHInbL0Q
ijOMHmP92biSrn2Lv1P73mOpQkelUruYhlwyWgvOGKYSPrvEV4pzszpeHKF5MLVQ/XzlWY96Dbeo
jqeOrVSzD1oVLksGhOHCYYA9Afdb274LbnhaveVDwLH4hNt2zONbiIwOr4bah4uTp/C8jUYhYv2W
98bW4rGEfYppDCkHgkmph5TXFJrwUEaVaKeL2G2c4hFR0POLuWbaLYgiJzXY8qRDYrraYiGA+0pa
2lRSpGC/LamYR+feHsD8YPVxJl7JwZjz4bKAP3B/ttLeX2jzn9frLmOXcPUMbiNhubCGvruqvw2o
ZstdNj9JH4JJmjIehJAKP+VFM8Rb9QIyoF5NR3tn8L5dfcD0Qq0rpeLN2Tn1mZWdqlRYjMi3W265
iVt9YZi5X4UscZciZ25nePw/ZOjkz+8THtl+bV18obNv16Udoh26RAStTDMiZnPcQTZQeddkGQjQ
7H4dO/Z/G0bVc++pRO9no2bPdntr6JMcywInxAW4nwUijzRX/5alGrq0YKmr3y6evZ+tWLpK130I
/w4kqoehN2BPtLyn/7AfnL9c42wCnv+y7iGJ9nmKB+84rwes5CWMfVGgQ3zZ3tPiZGsWLlJhy4pw
n9WGDmqnwWZ9d31YAoNiO3LLFAcqCufsJiycWYn4346U3VxGWshNv1dPROQFU04jwym1ciHWTLCG
xmMNmZhQpadnLkjlniPFJtRMjLuyrgOpIWBrz//1YBKSDXuzaXMjxkLwFDEsZsPj0Y8FloG/iIzs
cSOP4QwXzOFDa0IVsGVv6QGPcqPaQyH5Qk9YEre09cAEzZGErqktCJMVnQodtRpv+sHJjAHGY/3r
2IGZy9uEHhS7x7rmCi+/YItaHRcbTyQdyz3JdJ7CklmB2BpDTd5fF7xlzSszX/FoKcykoN6VRNJC
n86TL/XiLHNpnUfkFYcjPBbex3VYnaa39H8m2ury5+N8URaxIXpCL48YRtc1w5/gOdk3pjYmZdzj
2TwG9R9RzmL7dgaYe7jjEtUxtQUuZUWhi161yYrogjLO4MzCZMyuyVxW+naQfzQ1HyNuXlv5zyem
eJ/jpO+hOUsPq3yQroPaTLSsK3vxmYPFOV+wf+iq+vo+VHqSHuXtq9bQsdOWw4WVue7t8ljo2Bxk
nWLUeU5X5039Mj8JxtHh8iRL6LPtEuO0G5+wrh1Qp2NBXBeIZfFVZIPy0glTLEcjshUgem0cLMsQ
1Y0Vf/ApNfmV7KW+vwC647SO3iHtl2BEW8WggcTkV2tq4GQ8+SiD3OC6HgCj3NKqeJczmOulaReh
TTI4oxotm+YsB6SpiJquviE5xLx2FLsftlOk625YnkisBdG+EvjY4yTiibahSoO2WRsSPh8yLdUM
OGFrfWZWzIOUHgwE8h+mNptj70635Teb6+zB5CMZ5ovxntp2e8VZntVt5MAp1WBryrKG1kMxDuHq
+L8+swqm20N4wD3OI93Gvxg5OsfY3daalLFey/2++Nvofy7KTAgCYl0AYWnmUQKzOJY5qhjfcc4X
F68f1KiWD2y+ZLDln0/V2cjo/fc4lZvKj5IM2brFeuXk4uRojCZnqMSrDIqdXpNi82mfcepBbjvZ
2vOe/p8AyWtGTttQBj7NcaORPSH+T0opINJgjn1Dj18fzREPp1ab+yc02eTKmsf5LU4lcjUhYWJt
3D5LGZIcWCxCvkvu4p5nwumVqyudf6RowNeLT0Y1GQ93pQ3BbsZKctkTBsErFfDv1SEGSg/j930T
uw5jUo9R8UKc5mOUm6mS+EtmOKZUHrdR6/tt/v79eH3bpqEPh9S32NeOhEC76J55tJv8DZrTi2EO
5golPJuLIzZ+AbPyUbZt7Q1lvD6WSQdkTkeWlZyYtnTHorv7PxdmULdxpVIDcNUaj2aq5xKrorjJ
ygGP2s6/iODKVH+mL4brbWTaRYrXXwyE8e4zQi7AF90t00/goWzF80Gglx6nA3JlTYeYbJWpYGGw
Vv7skSHUW2MZ1gsxELpW2axDL43Mnsx3Kf99obkWG/uFJkQsm6rj137TQjQym/ljqnXOQ0+osxY0
PeKdqrgEZsYy6euc0Chk5m9K2j7xi7HhsAgHYzmVVR1XGL3Ykl8Xq9SvVF7ZWOJtmGJ9EpHClJfx
h0DFForXkgMy/fGcfoBt60R8xeKWdMmdUseZ652Tz/q2Lv7UOCMw0ELbITumFoLdzZ+UjSQ1u9sv
fJ7xrTuN8b+ntZiX87av+ay26ykliLJD7W7wxE7UlYbbdFqHOUJit0z5iPDCGeW4psvWwdt//4Rp
PnGIaFQJMyMz8Rj7thBTTryrC4bIoS0vvp7cTF5DBUZ8CcSi/K8QISONZ47uMYDjXQ6ZB83BzQCO
gyepO3arcgZYVYHIJB0yM3Sjz8lnuqT3m4E17QTavP4+ZGbYi5PjLkQbmAYwQOo8vGEkCnOhbGsM
AXdFtw5XmqWbZzR1dxRrI3yzIGsSpxxWpAzLjZyO9W0SnB+w1Ott8StVvE4dhtbQNuT0dX5ptyBE
1UzRxGx8YsxbLuMDK0C/iO2KRvnNTeL9vvx9ElauF9qbpOdpPik8xcAAwzN5hro4ScibsDLIEIFz
mMfMWX5L8As9dwVIMMWjMDiWdMuxqzSzd0UeV8BZpZ8qB2m+Pq7xhXD7myM2MmU/bh4CAPkRW/xN
CKZ9Bct7jsApD7pTszlvSHEZ56WXo/FBVbHRgH9bR7apF67CO95McLEEhfrbEGc94b2X59vXf8LF
IF4Af5qc8T7Y+wwdHnRr1ydEsDFKKSKnNoXwtQf4wSiWxHH0iTzsMiHeeMagJv9OMjFNZANAuLW0
BTnryg511Yj+Tx+ymdVSqq7H2jl2iGFLPqE5In9F+yoK1MwUiW+ffLq6U0itsEuoiXlz8PqBOREF
831x6ZA3kgwIG1C/y6wj3mkACcCOuaXQ+glTUII6947/3C5Roq+yxXLeMzh+eRcLfrAXr+ULElWI
NImUAn5BeAkv4FdVUtxwFmrXubUHKsyKfqdtW9DuaXlY58NReFPDIjbRVZGARIXsilcAlbJUyNYx
swOXJKEcj+zkMqI5IKdVA/YLLKNJuSwhjGqOHLkBOrbWoY0j2khuY7yygXtKYeMRPB2JaQ3OrqMx
0nXWZ67bqDG1b9IaJk1pQ/CwUuaXhcG0so4au1awXTP9T/JwRd4N3k14RPPUZgQME/gjX5g1Vau+
gw69198g2jlcd9JHIMEhK75rUPOG/AF9uTXy9U8VuPu9MRwJdQAmfSZPUMZvSoWz1wsTiNR7J0OK
MsIExfIC/ETzIcsUBiEEtHaooyFypArjKG+258cAi5nlAb/h6BVrtNsOOaoNNUKnTRdPUAZiHu3l
AV2qEY9gog8y9Lwi5PYTHTNAUfkK44cLZvuZLm4VvfXXHAeDgAP6jHTD0Hp2bgp5xG3Lvabozl+Y
CNkwosjBn6xq9CfHT3f41TxLdhQwOpn+tfJtH16yHJdifjOaR5+KLbuNyo3kqzdEj2/9tm+eEPgU
UttiZg0nSmm8FkDZ0CZsYvz6zhCmvmOoR9IWIhLm0J38NbV6UBCC8pbszulqiTz1EdZFchg5uJVq
ARxXf9CmiOnYBarSShdYI7Pc0qrzZqHls+zhHpbfCnwEJlsUg3dCe0T74bpJEFCLl0pDnI/FF3PS
oTOsGzQyOTzBwM9xHO40zWkHUwWJSLF1Qa6kA0qHKtp7wPwV8Xc0iF5lq0hmeeTEyJlO7VCZLa4/
osOk73PTVZjBJXVWNsgju18cnGW5uYm5woifgViE1GqLZpVZwAoKxyWHg1FsoFAPEf41xLf2MfAn
l0j6oooItg72XJyVuAIEEM7PC8THfFmlt+BBfWOioEuCxQoy3gsqY27z2E0abhewmYW8CB6a4HGx
JOfNvvPgT8KkumsZtjPG/FuS3YSLDJKgWdQYrliu3V7fI19cH8yJavE6SIiclqd+PsffK6JYPPTL
7JEQbwf3yu2cr4y5oKQ1CMu1rfjWNt0lYqTPZR5yjvxO0NTR8OtVLXWV9k87gZRy0UQT4JdPUadC
CBTM/gw/OE7U+eTVJu4cRjBrJ5nSranWo/Ovl9y2F7nNDz2AiPLz4aTrbO2Tsf84GCAFfiYyoTzg
Omi8Pe8EC6n4coFC3wAW645o1fYNAj/8Gk0XrRWuuUUBIljbJeOxY418itXZB0Hl1XTQbgDn22c0
XIKLx62iXx1a1yM9Ab6ZB+bhe2zpwjxGRVbr0wMGInplFGiJHuSurRwSs77zYjJCx4fJrPBAMG2X
eMksy+1TigoWyQKZWbX3a5Fcu89cmZdyIhOVi8D49UuIvH0WdP1vNyZgUrEtnk+p7iSZVF+sWac5
5/NDZQg9hKg/oVGtZ6oiL/ah6afz9/KSAnXbzNXcjyKQL5vBdPy3Kz3bgK1cqAykjExztWffvCyF
0bCwjpbN3IS+cMVQg7r3hpJ3RniIgA4DSfxfvGjsWA7xL0iPGVZDNdI5sSwL/HBJKS24RAO5MJ/h
9b6I2z8pwT4X/iHFuAgh8NnNIVK7ZvlhArCHVsb5T8+VQQt8ZmGFO9EeHZ3cEMWpAi9yo4/mncP/
e+kPYe9iRO7+PDd2Pwc5pJnzNyhxLtlXHbdccjKoJHFp9wAw/DsKOLQwxpWdVTOc9S/WTfA8xpOz
KQ2QLsr93mYBgjfQ7TdgI4+Mbe/1nWAb6qiDMAkTcyREGsCi5tLApXYd7oD7kZ3LYmh5jigQQXx3
SEUxNa037K51UdtOpqHNmlPc4fzo913aPDwn+LekoLJJtCPO37zTmbeXz56W7Hy+uOQxc0CBOoOa
T2ksmfmUFqc/aLgzLLbIU1vjMi+m3f72y8hFah4t/PJZOOX7lnNgnq7nRwu3cpI3nzj8/9YXKO4X
5DoVbe+78EbuzQ2biyUjQv1TBFv7JsOH/KDyqrnUcoZzxt7j4nqlfjW3kYmzemy5NOAxEKeKTwBl
/4DU1gpKrBmW4+mVME++K3r5b0lpMRXS84ttrZHn/zZjmHTzOJ1OagC4kKOWpoC9u85RV/7f2Dv7
8LOK4LiAqYzdaOFlqJsvt9AHbttmCU8YS4VnLKfRYsnODdnFETo353LIhzxY48OYPnos1/w5h/t0
0lHIdBKxL2NFwQRSZGeFQRAjcZizAeF5dv1DjMJ7waL0Cyp+aDIQ2SdjvPYHT2k01xBKK0R5PLCM
cXXOrUUHuskel25eOyJovfuj8GqR3tA/6XnIxkp59s0MJxTXvPLB8dF5zzGuazi11M/cOyGycoys
mWGby8E66R9LVQAdI+kYdCahoj28JhuHZTzzmPjq+TCa59WWk11FnAxIDtzg/Arox6JSoxY1OJq0
r16ufUN2+UCjyQp4JyB6FliOon5aLnUnX4AmJ8ZEjyb9ve0vfPgak/qzuB4Co1iZI+gzguz1WUiH
5QXD152BSnnK2IKp2Izzp7fzftb/64mdhO0jnnzuyFMJ1sXOCloU+e3SwzdT/lHrdCSwPUy4QHIh
Gf+0cR3cRXefphmHypyY1XpuRy8PQOgN8KbDEFHnndmJSg+Wkf4ew4ryvbBDjkvA/TQomkQwtDqx
RfnP/tjtWjef1KxuyhZYdByduNFmcu9lBKF6d5Y+vJIsxsNxIrbcy0XgFItyz8VbMZ3/mOIlSgW9
d/FFjWzSpNxhhzJbJANLzE6oshNbQY4extEtAH6aCn1Y1uXX29CUpuf6LHB1DRhLKGLhKobzzQUf
fgAiq5NBpP1ho3cKeXmJ6YxnETfR2vkMCoJda6bgWXIuUZyMxm5lthhH2ADGyGRQV0/fhg4lb85G
VkHHTT6QnOmiEY5uaZ36n10FcrR9KRZMiipsxpp06rY/Zx9MQ9cL3TkEF5O8DPHjvQKd7cB4Qi0z
pLSz7PW83/WAlxfa7OajTcTL3jJwdDW/DgsJKDf81w2/i5u8CSdqOyij+E1jEE2q+XKuf1ugke//
QMrUcC3Rl7vynR018G8eueXJRyqwmlASoqIUWw+b3CMI7889syQlcAI7t8si0a7ufv5Rf7UlnRR8
0cIuU8ixLPaXI1xQ3T85d6R0zB6NQ4tvp/mVk9GopCT7EL4kJ4iKkAWGv/kSEH4UlY+PMm7j+jjy
x2YktaYyGF7582p08JqTacQXL/877sZukJKrPabCPeOT7R5njT208t0Fz9Z2nXBxT5unZ39ytgIJ
GdrMBrMiAHEvoEnaVHVK1V+xfuGseFsycMdCJ9B+wxOPx2yQA1XXtPxfdeWRh68X9gtppfhOxCLt
AYbuONqjOqkydo72g62UNHryd2Po9JZ5pUtm9M0LIc/RjaFiHL//FvtA5Aaa5V8ROT844tby8bGj
Fz6/CrBG86OmeXWrtqBn42IvyPRXayCFKSWp7CMGpahHn9kOf2GeKCM3sab8ZhiWrzwZdj0BCLQ4
mE0wbdOnfi4qqZNLYqwEAeKE99CAfnCN830Ptx13igrwzvWLm70yz1F7HixGcSgko9d5AsGMmn/d
FrwlGa/tOAPmEwIRTOpt5gshe+G4ZHbARt6pIETkUsJMgI30o2vxzeRZ9zpsnSpkJttDDg49OqDj
AjRMcgltl4mCHnv5CYdgXk5RK9vTVNAEwWHOrFqk56GNDneR1P5CYtUbDl5x35rDKOmSIMPjgC8o
XqMI1rjUDosoq5J//bTqIznVshpQN+AMZOe+Gg9HJfdtWl3BrglzS5BJca4m59iTk2NsAU8wu70x
B7uelOxSOAVRetelIZ21tuhtNbQO4P0uelqdglo7M0jKoTcOROQEYybTsGApCXhK/glFrzz9EkkA
/PTEr9pSixn1Z/HY39hm1FOasGea+TVp3AwP1PEW0o+IjJesF7X3z2/ZnFF9UElJb4yHhWDVIw0J
vD39KUR5kWEIRkGhgOLbtq+558FGLiYzE2nv13x7p8FXT7DbxLre47sA5uQBTfHbUlXtuaGpPO+O
DbQ0c5R6977b9TDJN9japPuyvNBjdM8Agz6cN/RQmRszapr+0kpCvxOhIp5HwrWXtjxzMpSYH0Mq
UJkOxgwA5mgYliIOT5NhnjDa2UXlm9XopDYcXv+dO4OjMNQPNgUzqPzhh86PD91DANjBw2cPSlUy
TMBa2yBlS3Mi4/iyu3A2hH4VaKc3niuoXTut6jrzZ1KMl4D5YzdUbVKRlGM9563zzKpSuWmaHjGf
OIWIACJ1JDlyUKKu48juWPke0OdKscj8KcO5skSgkZxef5rUsbf7zv1WCvS4cRD7uW6sACENRW57
0P6ntkTgUaZgpai79cUQItcmtuMVsZIZFX/vDjf7dQ7iIyEKZStS6ch/0WakOXScGHL18QsSkHFp
PwpYQrhk4ENFqrQtCqKBCmuFxTWlVpeF4x5oXzgVkhnRnRxSPa12smSMYwZFEcWY8vzMTPbuqHL4
ACusKZsUnY6dqNvgSwDVSa9sdD0XIZzDSwR8Ij6+JO9F02ZHx7Xe9M4KxSnXC9JlwtiE9zynxl9C
DfcVcK2duXE5v+7mTHnJS9F4sHBoN2B4sJxOo3q+BFnJ9qvFI9LCjhr/NWDk7bzhubgYUs3XCwYx
+PqC4WJ86cyF9+YZvwO6YlKEmJYgN7K3OtWVdPC9iEXMyxGJnFzuoATYC9Ill8Mu2jFTqL0gmPyk
OhGq/gTXouJ4c4Wi3qWdzzAKm+tkbm1ZTno6mHffvcS6+K80AowFHEpljFZ6BTisoYNpK1SteVeh
wofTrP7yhaTSGZvIVR6B96faSdro/TD3c/sagZ7/c+X6I/T4GYlaK889p/BrYqOIstMHVmWEHnna
7cvnXNa64kceJZajo2FvnMmpyt4d9NON2wZ9SrzqJ4ZRu4eltOEiH8d6M52nmWWT6fXwuidnZ3uk
sTZUfVXLMx69amlSX8e3fmDHMIQ/3x4Dhsi9POhkBT5djkMuVl5o44A2u7W3QkcO5ZMYwqY3eVhJ
5u1hCzUWFey5LT+MzYyo/KcYhNMjiMv1iRE7oVWPJpOZ1f/ZskaCaZPP425tG2w1WCIotS5tpRNq
XbKy5pY4njaDs6z/8b7PnVKC9/iCLwtLrNb4t/Cp52+q51oQl2jQ0Qdpgqf//bx2wH82LTSkeuy4
Fy/OR/Ad+3kTdbS/RbjuX012ebwZZhzerP6ZalmA9RrfY2f3K5Y6MUXjUk8Bw/u79VXOUSWHi925
L7Pkg3/NlLO1cKQ8+nCaq7FZ/898hXA36QHGbGi90xFrGW20cM6j+8qWwWyZ5T6YnzNyHflr6luW
GwmpCRwmjMxljhw9NsSADaTe8443RyrAnetcUulcu5Pd9pjI1giveoet/SU7djKUavIX/Oe24dUU
aQSDQgLiRSIr8UfGhcAynwH1tsDLTKDbf/qLA7hhCmfZxeN/kxdiQrKx8QWSwEjPtVOppVK02s7Q
Hw7cIhoVDPyYcRv2wBRIfVgkuCReNvIcoXabggXmEgu7yu6jMK9aAqZ2OHlQufvqwvlGNEoIj6Ql
TucoLk1tqHo+DdQgEMVE+IcDZ7ghBJpg0gSJp2RUjEh2BYBHh4O2aboDy/r9Wi6C9hKc5KHx6/pq
Azeeih+2kCc5zFvl4NmSBWvpDYAYZPYex+b8xxuFZNXP6YVnA9QhFcIn5jyNM5imsnQWmMNbp44K
G5aDsYcI3jxEOjyLnCKbupY4j/aVPNqp/VOWF4SxU0zZ5KJ7AgLHRjzIPHdyIy/RGWTH3c0H8twr
nEAoSTr4xUg5khWIkL1QTap9eZtG7UWheGGzklyH5Ttxx/tX3hsb7R/ySYw2op8vlCVcXmtqnOBm
YOmLeb4Scss++3CqUV+aZzh/QnMo2IuEhfQXp+dT8vgQO/2S0dz3ikkmgcarl7WIHiDD3fGH7T/Q
X/VJmqe9t7H8RfLJP9hqmGX76EPiv2zrNfm+uX6eXg/ezMHUQaeRbQSqRSB+Z6u/vVNNCUK6GRjL
61QybJ//8Ac92U0cBgYWN9tBvN0IDWLFFhi0omJN3oC1cc/Dmztvtkq9HOoOz87t30Fvg11nk9WI
ajMkI3R/IAxyB7LWEbj0upK+SBL2ireETJ85n82WoE2rxhmlTLgiaRhSHdNv8z2NJxg22fB30IgE
HnvLstnZYGL1ZM2F6hKPbsxiAFGntedBxwKBrDdQHt0qXHSyEpry9L+nrGnM2zdbxB1izcWMWd7s
OFknwIIDNtT4EDbw/K0NieNVF9bzJfrslHtMQt+LqTKyp6oQoAzF+UYjhEi7HkbcJMeK/6tkU29A
jmBltN4JzB6mO2y8I8fw1tye9osTmdCDVeBa2bild9TPfE0Zxc61fSomyV7AqmW3s04nzy0lyEJh
J5h2PZNCHw+EwLS3vqrUxdxkNLrw7IqLquTFId48kZMiFxEzkF8T4D5IkUVpthohi/IOm0Bxq4tI
iAZRtdbsWo6YdW44kgzKV7hV6YPENChzmCzc7TRlRdQ6KDIaRiGkEug6xrnsseFXd7DuOn9OWOnl
cM5JSE+Wzbbgq8l9ve/DeeyctsWW4VUiFK8pcqpKeNVkTculF+8bavkpymwSN+oFOCykknN4CEw6
fNuiO0hnWQ1jvUfnRbfBz+e6/MczWRPd7CrCHheUwCtYH14szIBtjhGerhN6oECyu/3Xb7no6E9G
KlWgdf+mZyi682Qr7VzjynkgTKnM1NGlYbZGdcc43BAUh7CsZO4QYdZZougo2T/8wykQh/SmDR28
gmetet7cdMN5EIbwoA2raBFz5NzJX/ic5yzsV01ai6Xdbcy9jyXHuYboV1EyWYlv8Hzh/RX/OLyo
cPtfT23K/+G/d96zB9L921eAolrcw7c/QkFYmMN206tgkw3D1qt+tRUeiacvyouklbT5HgB/fpZF
MX2HUEPM4HbwCEB6qDtVGujl0QXqsvuG1y1NXfPMJ09bQj0XclC5lXD4iYFPUMMnjEqexAY4yPYo
wzCJnNEeGuNY04UFlOUDNedbcqVSkEz5A2hEwEfufXtyDLAuROqTHh90gnk4xB+yj6pBEksRhyfL
qWcHyacCuyfdOILDs0uGPBHohpua/8GxtLaYR9aah2yoqLPQGxqWhYz+73CeeeF/3mtEmlRaKtYu
Sweqb5W+pg3lyVvmF/E2htaz/Pw85I6I9pbg2lnELFj2X+TrZkDaP4K4UAUNV4oamFTw8KhkR/Tz
eczObitghqQwx0KOMgu/EX/mmcUp5xSpuNaQnhmA6by0G/3cIvu9Mm5HR5UZqhWEcM1gSHID7eTr
Wvh8frlk+/WHxJNErxt7t2h4qemien+MHli+TYG6j6AKqY4YgjLjLzJxbAHbzZ1ZDcAED3u+7p4e
86lERi+1OIOoSQmO5GAQZtqSIpVBo3VeoquN2abagafk4Glg5gYdymTOI30+hx/ts+VXKuw2SbJs
wSV/Put+63xXew4RQKKrxuvW8qYvze6Xg/UV2bpqtQ/hNuV9y3HV9coDaAgHHW5qI7I0+JrrMmId
NmgJhjxnhVscq+greNVjT1RzwYb9uqnbiM2W2ytfWXmN8NZoRTA30ldaG8QHmkgoD9140ttQvJZ4
+sPz/cgJZv9Hw5U4VIfKrE2cVfbZBXCHMyYf6W5uH5+1pLNPXJlAGBfJXIhX/jlmfeHEpYAoLHhP
zsV9z6LaDV4hVJu9wKxivavOfrJn8qIRYlx55LPdcswVrFxnOALXpBoEk0ZC4EDDEyiaRHSuqrWC
5mqtyEz++Z7gCuGciCjTemvOTSeh7EkY2H77XULP1GmBQg1ZI/HxukJgkoAu/PDDc2xnEesEd8e8
V5fouoDM4sLBFfNOjiZBj5NYhP9SG1SmfFaY2saxlsmiSGbXWJkByLObPEPn5Ld208cRExj6AUPb
vw8tkAeTX3bf8dmvI6MD9UzS6sxdMMwxPpiVgAUNKjB43NvAGFkukImrS7NUEpXn64xgq/Mh+zWn
L9CLDhyYZG957Nf7ZmCPEBHEHdWpsK3NHPb57WEkkqARLuoz2iySoKYiQp9TGX9h1VbriOBklZ5d
lzH1g9u/dWVBTMj0Y8P8Xd4dRy4GIlFZNRwal/hTgOlx0w6A7LEbEAyIp8i9LHUGo1p7e0ae6M+P
wpRSSo+FR/EgutbGr2jQIG9pfXx4s4HFUKP0QzcPbt20o7sl/onld+YnyDb/FT6+y6Uo08eij0UJ
KStSO4ZdlsK0aRVo90+sRcAXOKkry4tc8UuXxnwRDvVnO1xFUlK9hzDbEaNIrzC8mTTTtCiW9isV
m/6A5++qRlFa35kBRlB8JlQp4133dw29rTkn6Krq8+g1ceEDSn/lic42y3jJ7W/iGtTkcifTj9BD
o2vd1M0b/0/X61v/8xVIs+gQp9RGbC/gqi1YHojODYJ4R09evCJvxQYFJA2rsGMG924qBUwTapoD
S7MTJ3Du7qXnXTDI02rRzHgicrScPdKOC4pgePSLKasBeqiixe9f8n/WLgsKDDwbh6iBcU3l6wh6
XuQbC1F/H7Qfm5GicWG5lbZCxXebrnRp3JZjkmCcqOKO83NJaFeI/zLrK5NqxlDT27E2srI8z/42
byZXwZs4T3ci9y5oRxQ3vtq/H5HF4aLf1h4KTLnDefJ0TnK3KFZPQ8qQ4HiDArnfEKVm7yR0Oc3g
Z2ayzZMBXAHiJZErtBuH/R3CxmX3jQ9JakDaMFjeKsH+Eu2vH+ge+3Eigk1s6IjQOsUgWI/C6cIT
sFDPYSXBfmWPBRHUhJJDbEyH3T+JrtMMAtTaxE+qQYk2O1nQDPnmBNifrS4cSgwGU/VR4fTubdQG
RNKppml4TaY1P5xZQmC4bX+RQ8YqbtwoiOWL/+OL3dV2+A4ANxlWLd36jxeS7y6BINrHug9xLVxn
Jxi7L6bizjtr35t4ym8ECDZgHc9HuglDS2fnDz1Idn+/3fQgOnfyYfYj9/mswGx7Uu4l0+++xIUs
ogAlA0OoRNqG0e9/50pdhuFvwL1JLsvnpMCgpYzGUq0+dScgPrTMz+vJuFcABlYgHxZD5i60/ylX
HccyVMSO00K8x60ACy3LGERp53icCtZxN1P7M09zsXpzZgdni9+cDYusijxUfe71fZraq4ONNr/N
bvkD37Yt/azcFyz6HImya8kP7RtcuKSwRKbdx0k9X0PmDpmp9ga95TSd9Id6FAjw+kMwn/n6seXQ
c6P0MJYG1M0MSYZdmvw8jkt6M6tGtCzM2xKxpuP01DtNyD8yudmqDc4/Ycx82kKM+TMMoHDMpKb3
JLd/iDac4rsXCcC30u97qD9RUAMgUZqr95LVZKNhf7kdKL7/EH/AVTkj+ABkomiFUtOwwi/IKLgd
CL4T5NIjIV0bHtne3O6bxMKJ9p+UG4hkzCNz/FbJYUjMVkPQDfuuIrM9CXXflFu8/EWy5W8dyy4w
K7y+DvIZOYcKnSpndbla880RBIMO/HFCfZJc/uJLuB2SAgpnTGR+4g5XnVBfakSvtUA4f3Y4H6Xu
ucc9ByiIvQ8Nfd3if8B8iWcRzE1lEWdccqSjG1NZFx/11ZTDmTh5AoDgzA8uXLLYT2Pb6pkrk2P5
8YwmhUB0y4X/1juO6Hnt2EM2BCfCSk0fcU8Z2PUPZ9VZUKrvtccdxa7zRXKF4QtT0lV6SEDmTb8o
CNOK4i81gnhhAWq71pIuabKzoHUVR7vJQUVvIYYtIGii3G1l/GXW1Ja1wQDWM3upGyBMBRlYMThY
KfSXjcVYd3aJysoycrtknRv0Cs2lcIdaHIbdpxuiNXqv2zOJZMuvqNnzeRIPC6fZy8eflG1LQq+N
a8vfr3nP85Hz829azmAdR2GQFX8HFD5fq7oawr3lIpTbGP1kgbo/g7wUKoVM9re1jzR0GHGYYjf6
zK7LelJUHoJxrA5N3mpxVVkSR/eqILLBM/kHBUZBAEoKzv0z7xP+13mhX77abexCC7FPyHMlwA6h
qrJLu8L7z6P3J1Z2aaKcT94CSawL1CsN5J86ZPopC0nfQxDWFfSRRyANdUsBu1mPDtJSIEudmths
Q9BlpOeSptNKPgaG5dKnY+w4RqgkcO6uCAFpVu6DnNUwcs4OXqhyIEFbfggTXi0XgHbtuJC2UUUR
Trnm3DGAGNOPdhvXm1KDTjD8nuHl6f9eJ0aijKajynmUm+cBqw/cxTxQvxV5CtnzOoGVnbxLFovq
4C19VCCh2JCr2pOMST+YTPEJ7TnOXr7QB5ibKPlJ3iBs3jq10oaRmLB909v3S6NB+pBqVljrbrn/
KgrWOMGcmHdySlwBQAoQyml2CtEsbnBGoVt/CmVYGsz5AuEQqc7vxAVk7meZrnmJvMNS5ua5G2Jo
91jyuhyUcUNiHx55ds0vsYVOwO2wG3MAzIKCMsFtlonKhFA/QPmSLUrEctgsUmKlKvglu6bNadcp
Jv2U7hIBQYZHfaLCYwMdu4XVZCHx7aDwI+q/WN3/1HjwN6zGo5AbnHkLAKKkY3BXf0IKIkdRSl2g
LUrMNS3ZC+SmkS+rUmVV81ixUAZtJNZb2oR5RhwbbMpSApL2AxYpJIj5nl2NqO/OCw/V6Ls83ICA
AvMNwqG253QrxcizlaHLduhIoT0lJB+F7LooanIyHXF//r3PMupfS6sthnZt8+tHR37Uk/scLexF
vavlGGLb1R3eL1T3gsG++v7elCzwgUQwYCMkWb884N/Ldy4ehHbp+7FXHdVIPcwcwTzzIWV97LqS
jlWZpDNMiuDXxC8Pgw+LIUlLtWKTY4968T6tf6Eul4rM1wmT1jjGWJNGrTEqHz2qxrOagL7YBLul
nRGtMgqOJkItD3nafkO1BFgGZxtKjLr08a+OhvypsBlDfsuAhCxgM0rcz/M3i6eXOS8krs/CyGH7
6VCCtiupcJ6LD47nQ7z2Yjl8WJD3zrCNJ+9cYInaQ81g7ml9dGnaNOP+1OhVO/oo2AYenC0OWBDQ
nYySKL5syPqNqGq9Ab5qxt0I3bxfXRmuxnChV6Y3SrSGXGiE5TIbgw1OoOp+blXPhCp4Lk1Idehd
iIp2M2KdYQEvVXruUOT/OwCel5UdbXjfKzD2V1HVN+WhYfo5sh7qiny2zPcSNfcgjS/Cw69x2M7c
Y93kqdJFrJdll8wKUZxlYoV8CBg7zj/zpwszYXL1br8ZL83O7AiSzKiY7ziymg0LjrFwhFCInHl+
mr39BGCWgVdKrTT0BIv3XbtTMeqV69r1ekfuIddvFIYt8awa+7q360Gkj79Vbx/1XBiwqtWgFE+0
5qDUx0Hz8lvy9XfaEDp0wjC3UTjGYAvfmqY+NPc0xczIoNvXW88XHFQtq0pzJ+MAW7FOlzqkc2oV
4lOV+/3mUlcchNO1yumKUzaEcr2NXuRTddEOKkEt6lFmgJYP2JPqkWRyngi0mwPkRUIdWtefp7ME
tT0DoaFh1zyUfgZC/bNYBirN7FKy1xmxO3SAtRt48CpLdjhcJvCodkq/pd8oZ17Ojf143eJic1v6
EpOC5HO0no7+o6bEwoaVvd2rUuwoQ+ffG3W7c1leNiPs2qICIIR4HLd2IT1OOYUgiB3HgUGqT67r
6QzwMeBTiYYgCb8DmzXpDCb91Y4je9Qp48+UByqfGfenevOg6nUiosqIE5CQT3l0GwU2I+s9n3Xu
lHaXMcfvZlGquiIYbbnoHpLYEsq3plhkfPPxxhX69QAd499Xk1Qjj9+6GhZ/4KiXJqImW2nlbW3r
NE5ZCVbizBZ9rWDHS7hBx7vr+cIS5jan+1TYdhisLPcR+1iGgHR+ikuAIHJRCWjxRvADMO7Vi76A
4rsxqrMTeZF389itBnuZjFwhGlZtAKyS8wWd8lAaZNkl6sYXU30MMs21y+ICK1vS67BYrzDgPl1m
i+UWORiAK6S6A7DH8DExlDTxpq6B+Ynqx55/fYuHGC6mvImLapF/l5RxZwbvH02ynh4If5A7VGKG
J94ikFznBOxY8xEFmK69ssQuvFZELX1PBKr5qReRKr8jV6Bgw4fbUriT0Hi8cVQiy4hIKkE/TKwq
DSnKheYrGbjF1Cvun/Q0BjMVwq+vyXDXhZe3aYpKds1mFZVSN/FQK6vaLiGtZErf0DTyfJTyUpvn
5VJoWGocfS338+xUcDLR7PgO/vXEN362w1R0k0MD8TGW+3nOrBzuNWz6XMfy0KDkfn6n6NlPGZW1
5y4VyS7E+FjAQslLToVO7hjmLrHYQlxBiFvm6CAp/WuRmOzfqWYVS7vLYhgWrvijXFr+6XfgV6VG
sdY7GQwS+/JzPKEqEu2e/ac0I/fyMJUY1tqjfQ5v8BwJWRu4hwVa2/SxyCUeDvja269kPEM5RChZ
vikBzNiV73YYAYCoDyHGSdsdkRr/qKekuWZGYcGarkcv9TIXc7QcuM0OVGCKc7C+OsTOdJ+9Qy20
WQODeQgHwvz7zyE7n/SpYg1Akx+0IhmNyfSeIS34NNvUfHPEG0+vrOUHu+G/y2aulA9GT9oQlHwI
YgUxfGJujCE4U8XJ0GpABMAxlyWRHTbNTdFAyO2DE2JBxwYELEKqvXcFIog4wRDcB/CRb5cE0gCk
dGnKstGK9c6O0vl5M8b/Y0sngiiO/28MY3rcJ3uh8Nm4BR1s5tEP8ViMG05t2qHg3ftZmpsPSUy6
vL5bMtRtctxqnIMpH1XcRZ1I0F84DEZAJkY8of+xnBwvKsPRpjjng/jxLKecm0JiXFrR/C65V6WT
dkKU8udDmCXZTPoNbWtqtYoEdwFqnFOc0iR8ZwEqdO764ObBk8lFu9/atUgXBAwH9EF3pGOQkof5
rwLnBj3zGMFcZPqHYxWuiXDc8jL7J8gy5PvBERR7Xt27WVuD26PsIrbtXjBcJXrUwaXDGOlI/LR/
yHZv256HukGLsePH/b0ULA90skXY9BRLFZ0CMznHlRMHP2n0GElTDitb/Qdc7wT25UmzeiIEfjz7
j/Xg1nJRgnAfj7Xekp9csvmKpG8P4Mirt+PS8MvB+MkJFIrqZG3xTI0hwSWADN5AEBsP5CsIXwlC
sAd/bg4XEcoeV2rmkGVneohaHgZCUJ8KtyNlD5lSyZm8TOcAgqqC1dtfcgzcqllQI8sJLRO/daSU
rABPNzOpKY6biE4uFafoC3IkGDE6n8oonw8W57b+wTcw266Y0uH+4uaPdo7UU9QrQ4lHLJoGKyjc
kz4x2pLlA8Jb5FZQvz29Mfdd2aqTiUZNKpT2J18WFSK8/cPIgD9w6Qf3vk8fgTR+wSk/FuS8HEWb
imCqmZSS5P9Q/Ht7y1piyw7sAVJWgYyOL4q2nktB/VWdlXKE+DEoSg3I3lwYPTFSktqfplOYlmI8
7YCFnh5PbVD+J0l90VgXpWEtTb6wuAtj+9OtSQfi9w8of4nQZNP1OQdOFcqx4st2QMIaFzOEwU8v
kzifs+i4e0soFx2jG8ThjSpLZgE4Q3pTPj+a89M7CR3STeTrMioVXeAFVbOfC0HaSVvJYJXznO36
LZLwFpT1BAHsYhCJJ8CXnPf97HeKa5gJnByKWoHKIYjnQGkCoX2DjaEqhBWlI3uNobTJ9G8e9ekr
zfApfqlBGUMCRnR5lPGIWlblszcQlJ39NapR22nO+cp+35QqaaWuG/N4KbLYZS/SXwrZFapzMK78
gq5sob6LvPA8U2mDQH86vzqm40QvG8FWBXc4M1ZG3Zz8G45ARtXs0AJV77Ga4LfJsbAtYbwiRack
eDsutTzc79hUB+5azGWXHxcfplcJKPaVVHkHwBzdDiHwS+yRAtmLFFuo6skm6++6riZczOUIT+xr
ayyOtt8NDFsXHtzkm/bEhGwQ6Fsi67+fbBBRpBe5HM4b9e3oloWSzJAU9n28OuDYcpzwpnAckgn2
9F7AFzMPoax2xUsSJWEOCjipEV1y+Mx4ZTjkqD+3Iu5VjtNPhUz/9/b8jyVCSgnqAL/eiULR2YFl
MslRaye4fnWGm9o8F53TPIc4j2FgwJG0xraj/GXYinjqBZUkyJRfPbv0r8qZa8IhuCReS0mycqNO
JO9boP2sGOi5BJvaIlk+In9Pv7te1I8lRVvTl1rmFp1nus3UZyU+wA2ZhalitB9raa9z23b3cO6T
loZm0Duhd5q4K1onCUmqh8zAoRwZaCSpCkLtnUMsJcqNt4ZUPcNodIUMyr3F2OqyDqtQUxayWl4/
YpzoGjBdwjA4Yo+XF8yPOmt/Kw/DQ2pmmT3TCAWsnfzK0EmWaom5jBgxwjNksk0Ocg23LoCawnbB
GfyjCdFFzL2E2nnMaRV3k9bOtJJ/g52Pi03q9f/MKEWzWvUdci59+e4eda8l7La0bh/du1m0QjV2
gcBh8sk/zsYhZpXVMCnlG7xqT2sAd3JopJmV9TBMjW8IUETSfSsGEdNJ27qdTV5si0Yass5l7EVq
x4OMP1aM+BSPTTdYqFpSnQMKvf63S1uMv3ocWfjKGdfUFeFfN9Y137/+zJ9vMVKfUBxip9Ihtxp/
MVXMzg7jXTtKELAVAenOiCj9t2TPxLhpUXZfsRYcvnVzLHOSPbgNJQYR0XHmK3jV8wgW+y6adKFE
zmgHId5kRC3e/wNbO/1/Y8tj3+RStM+kH+DyFLZkzDr7XqNDzz7SvCrqMk4itBNB1xjlH0tC57NX
6L9ZyyX8wzcI0tehEHtKRTPzEAy41YE14+FfjueL7FL0U8cQZqa8NDsOwPWh4ObLXMk08w6IKmV6
QS0jiXop7RUyaD6t9YlFKjcaOyV2Yd0zWTsF+WdTkQysanOXm7DnNlZ8cP4hYghK+rP4qwjf99rT
DIwHywWLbcMa3a/ofbK8twEIcyG9/iUJEnJoqORmEWnJ9ufVJZUB4jOV7GAg3QQmzcw/Dtslqxbs
vXdFV2+H6kCmNWSYJXfSHqYaHYGf9BXclsdOAZEu3NsoXvCUidUl3o975kBIgFo3/RmLEIRNKvI4
Vlrp8q8yV7Z/fmAGyhvtNBj81TBVL2+xLmE27if9I/j7z4xUJF4gwQCPWkFfy8QfnLXT3czCi3i3
7U7gvAF7cdh5wqeRMBGcmXMUay29HoRVPJ/oj3tKAKQ7CxMPT/BCRjw+tIdDMlVlFiLFXAsT9FLD
i2Xc+Pc5VcF+VxNYXyZIaj5KQ6aImJ7ziN5irWrYGWe4ARyImgvGXaXyqb7X61Gwzm/86HvXkp94
VK8EZn6FC6NvcB+lbDOVpcDoP5cWi6S8tHPOzlg3eO3DjhaK+E54FA6PSbNN0DWYQ8MAbduMoUz8
Jfp6EZZ+MenpgvpD+sZQ26zY/dRNLwoCwiM0pTRlSJRbzCCw8RXwZI91JZX/hdbTqxALPt8FTBtW
iyF11PYAegUycWZLIos69KcT+uhRBtUyLfNhXAZbPRzmgiKCdLfHEbpTapp2fulw514MvEIdyTfb
5aYzugpFuoNqcblKzdKMeNkmQTKy3KqdZ3PpGlcObHJNIcErejaze5T953vcC6GFrsuOJ4/g6kzs
uT6hls/NBYkLm1fUsbAosVPb057hCL6jmsX8ApGiroxs23URHVfX4cp/MyYHD5lm5dE0N4QovfTa
wvMKjGtHXYZoqGsVtfQLEHzQUdHaTB+9dFB/4kzN84h6wepSYNmFYsVdH27XrriW46U5nRm95pv4
mJu7sNk7EUK8Tewhc7EDxzUidy7qa8YB81sWoOMkU6hOxZk+eny91HanD1ndGCh34NkTHPeCdPFm
nGa9E885bB+D63C5XR8ILhkruEGrrhzUEhcazAWtm9QLGDQt7oqrc9/NWJfFkrIodMKWwjBxqoY2
sEWJEofRDNdR6X0e6u+/SEF3/Wc6u2fDeSfV8SnQtabqFLXVtVoIX8XMx4WginfDhywKMh0m7xp7
dV9DfUlwIeBkUM5rGPWLe3nS8R/ORN7JEmeJX4HRDzPJZVTJWDxIxEbMETJa3/mIDsJYR60OdfTs
/q1kg9bxzMuyZ0Oo7XUYa5WmPozRiD2fZZliXIGhrtlai4Fw69vy0FKppxlaFZrlzaf7Qq5QqbH8
jkjZTNBaC3+4znnlmCiEfwZRUNZhrRVxrQwhmhLdeI+1a+kXcU75/RK+P93ZFf6x3poYTaqaYuzs
aUQWWugZulntt/I/ytXDtgs5OD7+lrB1vITDLQp3woOwC3R98FYfPQZQBtRvNOyZ5GJ8QT08DijQ
oSIs4D6sJ3Y2EzS0lKqf4vWIp8U2qEn/KiwUQyyccPcuuJdkLXzj5G7FTxyhJMAgr6WoEbl4gm6F
AqnAP3fLNCdFZubaJzbsxGXsvQcZWaSQYzBq4zk/eOmLGzURb83KpeQqcmtNsYBVW/0V2Ycmq0SV
cneuXdrNxDxP5h4xEtmEvV7CEIQsDpYkF4inO0twVKZQK4pIxT6AruRarrEY90BVXMc7xhsYNjL6
vZw+4beyLTasg+ul23enGm5B7vp2lI8kuEsFehmPJmDIC0HzvD6q5pxOPMIfwFFEteZfq5Qn4A/c
0j+CHuKNBwDdzPMB+Aqs9Q7cpMETVRIZ97RE76ytT111aov2d/AICVfRKyps5A95+VmQZM+lzSEs
UfpHl/7lENJApT8TtQsOY6DwXUXAkDJoltdYN92mWDjtJy8V1HO8VAzKZXcykCipGeyO2Rs9xutq
wLrXQ0dymBNnb09wLJ9IV2MR5l3dU3Ij3QlaOqza4yROjs7Aqt237/i4HZTJvTjcPCCJHvEIHZhN
82Zvuhw1ISlPFgQ/MHNrRC+81uIlL2svRnpMdOm88RmRg1K3iRQlDZWgpO3fQT+oXDKgAZNqvEki
N838iR9glNy7Lwf26DjfkTb+HCzZr64M8yrxY+PWCn7f6BsWuEuug/fil/z1ZUgKJi2ca/gcteyw
y4odIZgitXmdLnDmBI4N2g6FwXtfQhSOeUiFmmQxSPpWzB17iNWZLlwoBkXnb3n639rYTSjKPdNR
g4C0iukb+yWmWSuQnAN7SFUnwkpkHr/tBiGoZfd+9f0SsVpPV8Mij3Mz2XP2VCHJ/ruB2budwbZg
A10rUR5+zxRTWrc9ttlWvw5YeTKqo0E2EMYaEt7y0+bG3ObTt8XPSqDKGgt960OwnJGiofdO+s6p
/JSC4frAtfJHttZ23gePdZDKw7LnnLzI4nygd4G6yc5IBzdP0RixPMUrNgFeLzgbafpMvXo41Zp+
Pn1Nn9pGMnB0Rs/QHkBeZkryZJIBX3zqt7QP1u+ZmqN1AcQVUy9q32fPSBgwM3ZE2yAn1EIQYRMy
U57Hy9ykQVZY9L5KxxMpT/RhHrBsEa0ifSf6OQrrBF4egDMPxfWzS6QBhrb2swVvgtOa1b/+R56X
yMLRPqfcFiLtVrRNnfTfDl0xMNbIg7i2Su7VrCYBQU0v/t/nMPjYNqliH4EbjB8IcB/JdY4nKc0H
kQAIwa7SRgdhB2JMYvPNzgoqLb5t2GDtG8g+05VLwEcWfbZcryfiYf29oYIIvDBDBycCC0ZN/YLg
+CZeLXt/266mRzNGReetcP+reSREWxTwYFCfHnkaEutx3JDIa8ZpAxMSIuE44tZSuQQabYIGiUGZ
FWpE4ZilAOiIZOyOY/aDaVfZizlt5FEkjKmHPisfxi62oYFocN1JdEbAEhYT3OYSS1X+oDXiWPOT
KkUXXOAUd6iyl0Q7fIsCUbQhMyuLU5vTPBhuUmBwHTAU7uRhPEBjTvmxAlLFsl+tFbBMQEziU0nb
3B114N6cgxhbthujYRnNknvxqUj377lArdZKTwXDT0kpat9t8nfC5DIDfXgr50kzdbYs0ApQduiY
40woP0KB7DG94/eruWKGhGrRcbH5EHFXyW4fAtNf/3jXiimUkUlGwonjTlYz4cQyu4+0RLtX+GF3
iDz4UsD918tyuR83CyXE+gIeqD8FxyIsevHaYNddlsCYFfM2HRv/LKw57/ZzyFPzblhluohHwyYt
ponDkYfTkG0T8vhIXtgEaN7TVARM9hn4aC1HPdJiPRu43CyrhyC9h0nx3uZr8OVHEYdilpwC4Pk0
S8awsq1beC8QSm7oPh5aOeXkVYGMJVvpCFvwmyzKvjcf6OED9nTu81FaK94HWx+ayOYLzqO+KtU6
kcX4/mwBjsFREeDMvcDUWHWHWk3ZKN4OhsxgiCkDso6jKNUR/BTerg4o/boIGUqVv6fJMw7mawM2
lJEhpTAZDq14nF81LTiPDV8MSernHGrzxqzAMIc5ixqVFavkLtwBfDFV0aTDGWeTx6eKAcJRKIst
fEEoBUrOPXKpRk3/MEQqlzY33lKy7/MFsWctsMfZvEicOaxP3qgTBphel56jBJ8kGw9k4FMJ04aM
xgy+yn37a0EzeK5ncdDGwlE4uDXXohXmu4iRvHs7U4xGv2d8/rQWVqQm9rx7DrpNXg9EQgDYMcAL
37H4pibXxZ4UN3cT5pxoXdKC0D7hoTPHDLkePZzp+HYoGuA6S9m/3d0qTWdNct7w80OKjPkMq4Nf
Ot+GtJbJsbWSFhnQ0WzD+exH9NbboLrZfdclAJk5+A4V6eZw5Aeq1OCO9N2HFPAQgRU7LYLJ6tFj
T4giYYNrcYVr/hWwkT7SiDFEagmGuwnadLLUdUn/3tMcHKCddxCxzWodJvcjzPiEMAHaC9dopxPN
8ciIdrXodODo6XS/CFz5LzMIPuWRCx4Ecp0fpqkO9r8X0d7/iRNZgx6Bp8dXhfIVe7wkeClaeMfu
ms0LXt0vhx7EtvBPl4qG0DbZ3KTYyQvfTspQ6ncd/GTXvaiEnxjhLpe4Xgw6LlxsBCjxuCfCPkG6
BEHX/cRpFIKzJLe3QYSs+FPKmXjpdad8xweopO5sGh/k7SuXhxqApg/4/h8P1DwOr7UDyJWOmeBH
vP4OKuaVWLdZxssiFl3L3vIk3uGRwJ/JSwJ1DzLlw+oJ99CEf8fze+c0YM42zHpBQkjwFD90Jhwm
RSWNUruYlEKySWU5zHYhOSKWZT/YUdEMY4T94vJ3EKQY7WKdEQOHJr3eHKY1Dzjqnm4qLmYnJAml
bSX5NjNyyNryXRuyDokvFdLpb08nfrgQMN+4o0XmqWsvVPuT9PZfjErOHGBeAX6a95tlvkcazG0s
Zs9tM/Hl1A8yxS9gvqFpYnsVbXE5mbLHkAy8VR8MHs1SzCPwNX9S3onSwoZSV43ys96zZbn4IBpT
5Ffin3btxgs3/cgUkMDMgDfU8/v6tE0O5ADvSk2LzLuIgnk/MtVwI7WuEtPU839/LxQa3DrgnO6g
Y2kTFs8kYz8eBttB6rOBZMXpq5uahLtITufZlCr3/OKhfWOy/yQigTIGp0PW93Xb3OI95rwt31nZ
UuiWk8jUGTGEmNAhKffmOfNeDOoJE1m08yAdSeXCZjEpkPLDBMi5aYpLoWpl+pmzBTO7n5avCwAy
yicVyJLPFrmjLCA3kQGtuUJQBJUFkIkR6lVEiHLNdtlTz8D3dCglCrCE7HYayfZSbvcu7j81eWsU
D6RPzbgGzlXs/TAsmpATRa4N1cJrD5MlxTva8HOTy1ZNT+s7WOkKOi7oWWcWiy3wlaWNIpZ1EQu7
DXrCQlAX25P4a/3AumUBVicmiEe+PBTyX762XsM2MCyS1AtPCtcaXTnd3OiM+kNsg9CC30ZVuy+A
N8SojyMTz6C/WD2hHuS5leaOVN8F/SacvRUgBOFjOgnkYxyh6/p2hEYplSU5hcs2fz7TnmbakBRJ
/cuRh/Q+aCrsEnbuek/pS0W8+zkCd9Z7fGtYoX9cV6pjFSYQargSnsnu+wxOkES0xE+wAUV0kWva
n7DG5OfkWlsRfisgQCJ2GmyA4kI807X4LOX4iWwRGo/sUuk/yVt9XOQ1XjTdaK8rAoeSohRDvFoE
ReRPxYzisK171v7wwoSrt76ZP9xzbFqLkWzOUr6H/eAMVWsXKkrl6ORnFHgMNKl0Axmc1gc76Mla
y5lnHKDkbBYYiS9TM2mpoF/hlXGmQSu3kocO3luNpjlJqH4OoPfh626GE6KU63PLsWGYQPqbmsT6
PnXI/jVHkSUnyI4qKPCZixsG1+E7/8jHoauw65l69b5oaC+kGorxvNkjf8l795i3GencYAej9LyY
8RP9gd8RfTNgB5rrSGMjgpiA2lHSsMcg8kBGs3C3qlfJWDE/OnbjZ6f0luOw5cK8PoiomkrWgH8L
i1MoTP9LSMhsBn4OV3Czc14f2JxSMh238PKSx6sZy7C6uFn3J8oneUneRUGJanF2zfS7v6mznA+v
fgMzqzSqzBA/ikPriT5qixZGRk4rOVGrkq5Xud9bmgIKOzjrsBl6B8y8KdWFmF692q9likRmbY5e
IJ0r4/RVqP1gpRlsWRy6dKSoA9/Qn7P+sd3fKQnD4xDU1jBGyB3tnGR/aAw72uR1L8xRo7DCHBVn
7F1AUZvbS4hCHjc41c08HviAoHgk0QQqrEsVAnPFXyC9HcBuwUE1VRqcbOnle3uyMg8DaA8R8mtJ
Skh3nlaJYO/LEffZEz3n7a8SMEVXp3uCXZCX94vyOAoQj0TiJNkBvweQLsjjFNTTKEYJgvLajMBj
enV09jQSQISTv76M7exqRqlQqksLfFOMxvJ19MUj+/g5dp4TkAavUxFdtU4E9S7y8E4LX6blmQch
mLOak7t1GeC1DAUeU4ya60IP3WuBoe8mKIyXFm6d6Zi9bZKmXzS6AbFk6NeHEAoFW43osRIOuY47
paYAmYMRikyspZHFrTQtlChZRcV5wzNBtt5dUeRZLhyMGDZYRT6hLktPVSjLZA00nc0wEwbg4YtY
/4mj2QDpXO+XmuvX/g6VTEioI2pj8gYubu2195oNm7elZgefjfqS7nZs2VE0so4gQ/tlOpwJtUQo
TM8/z4aIy68RBc6clegpPSTzjFnFiECJCwGEcY2kX4Rb51Src5+ZRHcXxiVyePT1Jn09Q3IAmVo7
no5+wBSvqeUk0bX8+kENe9sC7Tc3KZQkXvReW6oXqF+VuwzkcBZWPTYEajQ1V+X8W9gYPbmgxlei
BRrjpk/AeuJdynTiJOGoxUmspmCq9mjefsyKT2FDrQjLdt7LomTrHbIDWGnDtQX4RJw+1LoNUZ+d
pJmoosznQKc7jqkHrdNGrmUmN08EnnVHx+T0r2qqNE5y2DDzj8azGdu/AF7BiW3Ab3dsPy0756KQ
y+EGUS84VrHa+5nWIwn9xcKVcx25J5tZNmr6y0qv/8GS28laQ2ZGu4wiryvDr9+u1GFuVJu3agbL
/WqRQBrPdttC/O5do1TTYNYAzpbThVxQHk8+XKg3FDSChT/hXja6j379W46HqIJbM3aEN59o+2sM
TjkoNVUES61SjHL5WmUdsZezZi/vMAR8atd8/klx/uzy3sj0EIXTsT+4K6JKUAQ41bSHC/6CR3ER
gEtGNtkoqv2Ujo8e8F/ez3nGtvEZ/HTjv4cR2fEpxbLuhbq7dzl2y/OwenAeeacb+eGqzHUBfhNi
aNR5Yplc8NiXPMWdp6rjBcdFZy30z2kqmmpftjfhtFvxgxSAwRa3RmNBZjs8RETuyt6r2Ycsbv3Y
IhjM77giffwJrwm/Vt39ZiO+NkHI1jax+phxdI/0U8SVWj9dxtnFRYwl0xdnBPDfW3gfck0LI9JQ
i6fDsWIsYsJzUh6aYgmWVaZtOD+QIV+1ItspEgQxCsQuDqIAZmMe6S/TJ/GOMTZQskhWPiFfHmxJ
wtcyog0VulY4O4xPO1tdmNO0VK9Pmu7pH8GdTYu3rErs6xt5k8EY3HAAcjh7KyUEdEybj2oYtK6X
DCLKQFhCsXtQBU/t5ZzKj39uhcOydoBh3KtBh9KxiEmUHAEEmn/0SnOD+Tc97hibbN+zepSnZUUl
VuYvh2OhWtaJJBYIioJ2ijeU4Gx4pa7c8+FDIVRHbSCZUFJmB/xW4TmztjdpYV944Wd3jRHL5dCN
f6Q7+yt/PfL5HnmuFpRfNvEa5OgI3Ud9QXC8yXRoPvK6l+2ZFPKxXIA6RUD/w8GakfkxfRGcDt+Y
VVSvbqq3I5ZXPfGKcixkDlWU/nR9NOBe96LNMYRvQlJjrBf+lQGEiXp2SmwNkFMs/9jaYa7KRrmJ
V/UbYm+Met1+8/+zdvsYmCKa8/cIXiOAcfDdR0Z2ZKUgQLDJmgQnkq6thLr4mvD57d+fyh2TxW4k
Ea3S6xbatC0XYVb0T/j3/eXJ8iT1mFFSwePYGJK1zx9xt4OxmClhziCL1frQq8pO/oClaz1Bfyr/
x3IoSPbDzsNbvqd0gdcXZY+ZimfQ0Z0mItd+Rs39WTkOu176UJOCr1fo7MabPa9POq7YNTRRVwrV
3PYIY8DytF1LdRq/DNhDBR7KcaldFG1FtAfeQGLZg9VgZlWTQwP5YVhMOq1e6PnNEWS4+rRWcsHH
gwZuZ1SRDBm47f58bzP4T2OPT/9J0H17NjqoixYhEFJqOmkHtggvNLQ/TR8ZlhVlVgmTPoWZ/EMv
Cy+2mVeimRDuOzJ9k2/RP9a4WqXYMMh9HbfxEQiBV4HtKIsMtxdSdsYMSlkfyD5pRRGl0Et7k+6x
J7fH6fXLQUesn8bcQMBrH51qu9oNXbKvoxqilrUVDb4hsNhX2k1kaYVJOHJ1imDgEQUxIEdrIKzr
Lb3zVM8C3b/JOce0pn5hsVTHCJ24Nawr5m6/o8RGfMar50KXaAGL8D5fUID2T6FUMjhEqzkLrBkS
9L0hHQZeFG1Wutj4byahZ3YfWC6Ntr6vbpZHZJ+V92WcUsKzIviJOC/LiuNmuuHtcd6gauM75ykN
zAoD1LyreDJ8qi39WPXVLunLlYCUQyrG7flaBfde8pzV0S3JwziV/Q/lHeiboW/vCAe3+9bqkmvu
3TUkougN/q6V+44nuFMj2VgL866MqaI/p/93pQiLRduzRoMlXuoXcw0RiXJeh02ihp/Zt7opW2AT
50V2RtrNlaagOSrt7zgVkE1WLK0R7FfdjsVb7fgE7cHzdXWPFSOYnxpe1XAQvXjt+OZcKWiJvqKi
KeXbFH4k9wioNixouYUdLWoLV9+6ZPEpN1GN7DQ7NstG8SH0pdkYwnjm66J0C8V+YePcy0UeESy1
9weB1MQ5zQPYIic2d4AeUmS70AywaL+o/j1TAAwnBp74HsO8htscDLsXY1xyW2LtXuKpG5JL8/Zi
0RPlgJ4VrG9dlxmGUoW/YJ334VypWsShdL2atNNyLf1zlsIx9WFNmX4BHs8N7BkN3oAcpkjRQkcO
ws4RqVUVBZT5m9j7bHpd5/2PWH6EzVRYww5IPN6gIv6sLSHKOB70RLYboxRR830HvqROTkVljbFb
96JzTrIjYDGzqysmFoqTVoueiuqhG0RH6qufcZeOIM8UGib9FUrFKBtCTRKYeotZtSCRPd0S7ESa
vjcHOx5wwJQ3PO3qRL6JGbi1gZ6GLjMOev4N6td0BYTzngtlW8UScSJqTqs96qJ+apNo4GCztAJT
vB+lGH0iJJ/Wq4+guc1trE+BBuS2lWGDKpfINVLTkGtZ/8oPt9qZUBJzr8LdNREA2TsykCq+oVCl
Hoatiuu7seg4C2Llr17awSf2iIDL2nxLbPION4zs+aN9Xx9GdijI+bCoVfTdiFdXG7pK5Gk4Cc9M
vM7dVcSLUeH3cIeMwIezktnRZCuUGGw0fqQBxZ+r/yf1Ro37R+vsbowTQEWVP1RRTuPNG8Lq89cz
JLgMxcGtAxnhyCfaTx5b5w18KWPNpTuQqVgi5lfR8LnvIc6BUEY92uRYHoOnqMpxg17sLY2V4dco
g6ZwuPVOMiTBpAJJwJuQiY+M07MHbGcjrmbetjGUFI5Yg/mD3rlpZflujkQn5lJw1ODjmau0lgZM
4JH33aS62f9+h/SANdSy0HiXki6XWUqB0RTxZHn9unFKTHgF56WZFFVLlYZoYjXecl3KCmWNoacB
d+7kOa9pzBC7U2EE9jIDJu8ukwXEzr752zjT2DKgqb2Yk64qnz439IzDt4qAqtBCgJUZdwm3Ya9q
Vw/lwcyijYoppy+ph8yBE/HV7r+lbwa//7OCy7T9aUkc0cNvsY55PFw/ApVJ+mgCYiQud1cfFRJ+
ocFzc5ucvGGaNCh3J/g16ghU7sw8Y6braFyZczryy4+ZBW4BvHu5YZekNf0oK4GD+S80ghCm6yEU
tyhtKrfz/mR/wbIVRfvwZz7c9gAxh3T/8o+dF4pqYu8+jxbRkt3RFVc3DOl+LjIQK5LYK1NVOzSL
Q0Nfy6RVSbTkLA03tpDLFWB4zoHJPNmsZXsdcq0dbEY9SxTbXe04DRCTMgH8TzuxArpZ5YPTUNJW
w+XHEDWAfe2RvKkZMnt6bICG3bVK1fdLL8Aj4m/PNCSPQwG04iccqjwgbT4Dk6IwUGg0XpQZKEgy
1tH6NN1z053q1i5YDcpcW/DovP+ELCNlFtz2vjZ/dz1L154D3fAmOjv20KfITCMbH7AvA4OvYMxp
5YwHhMJd63C1seetTrp6Am8S71HrayXeqE7KHvuQGA2CyW7iUpe8t5USd6fyUoHPKcIJ6xMbngL1
syEuDcLXj1A/SAFun4kS71lwpORfFdXwOfAkbqQaWbx29seKKNjq5+jz8YP4FqxeAKXsdJVyYNOx
8fWBYFn6rT6uMHhIfbR08oKqa/SCtVHPTSHUTMxGl0dUi43vv030L9DOG+JadCvUQZBpCJ9XN+dk
fSGZpy1Z0FF7SYn3FPL1CB7+oyB6bEHCX9KGeRfUcCFCV85+8/GVd4hCRipqibbqE8Z5OeVnPxKT
TrU4CpSpisQN9W+gHedDDaJ7IE4vIeONnCQD+UnCMzeOH3nAsdbvch0JaKYEyC6RwG0lLdyzetSU
QWAlwbXxduULFhcuZWJRf/MVoUi4vPSN1Dl7HgrsVckzGaG3ZqbU87f1fhd3geG5wi2+HQMLe609
ZF5wtqb5cPduuZVVT3iFSbO+Nal9TVbpTUNq4ZgmHvCNcQnXo6EmEP5PuvnrbIL153+9qhgsXjZ7
iOp5pGJAV4PnjwVDdxb/+dMzT2scfbX8/c2kbaksRJ1kGT7spwvW6hZqdT/fcYvDt2+RRj92Snxb
LEPBfKPqJud6MLTprC+swKnzT4safG8RwuVDbSjrVkNzQ4AvEDWYNsIXQV+i2AEdAUP/dFg8YWUg
kmHc9+jR++X92I1jAhj49z04GDdqkEJ6JW3W8NV18vg+lf/+k6hB58NWLYq0Ljgi9l6WNjT40AIH
scsHoqTcEHJ2Rw75CKzOZysP0XntZn+ojqae/PmwIJaJkFVC5CltsZ6Jo+Ri6Ynqn8KWzyIWcXTk
dIAoVDiHMARMf5QUu+mmqNjBs5BT1mNa+3BQm+4QXtwbZtF8FPh4IZp92sRWVf0NBzCj2ncLG+MB
dmdKzSO0aYT7j1S6iYGUZ8xtu2w1oc+WeASdXKXdm2sBq1a+icFRA03Ik0/bsFbyXVPGuZqHixza
aQSC/hfz47HAsgVqyPdud+9oueQ/NtqTaWoGVAtfBIL/CR7PY8zMgKsvb4SmTRuDi6jVDAXYSr/J
MU4WtILlYLnmiIRLOTgQnCbSdqud/kqVFQNe1mauhMMkyG2aSqJDAtApJbYBSRrnuyAWYf3wrH5S
YcLbwG2i8R4ZdMFGr4zjwnWb87RyspKwM5DGJSebAww2VQg85MobNMo6OJyxGlIey84Ep990pz0e
WWJBEVlwTFgpGKbyi60Bv2KTKRk7PUo8VGQZXSmjMHE+IUa1QMYCDdJOO3ucOhQyV7Hfeg5lJoh3
TdE7YLlfW6BxpDDYpxBEGSaccWGFdBeSVQgaPZWCu/JJaldD6zz6IeTohH5YPss9dNm9SKVCHp1S
iNDaTGrzdf4a5rFrGoG2eVu/hnXxj+XqsJeWd80K0WYgrxT3ZfX2OlbyAIhJsnnlCmaTBeyJKkxz
9Lj9N05fzXj0Q2osXqCcGYwLbuar8+4wOWXqHD+rvYbny5NZ+ZaDJeSkS/EfCXxzd7TNDGZAx4nq
sFeSZ3JMvQSb1qQfb6JxRn92KoRe1pe4/fZpnSXiFpx31QEDZUhYSdxSsHeY1Rw0J5O8qoU/NFCD
3hoQ9U1JmWimrFai0kUb02JLQOScL9zIPDKypvOim126IOE0EFryv06qkNcGODjsMB3DrviA8idr
3Omdx1vUJKE7SEc7EGvumWRAfs0HPXUQktXFHen40RyfbESqGWtAlveZAns/tFlTmJv5qRHsukMK
CUdn6DSFqDEzX8fuENeu6a1ov1WqtkS2rlGEV4zuYJPeS+Z4BRLtcodv/RTAFhAMMM9avIlE2tE5
iP5bx6oCKYyI/AoMKVgtrq2n1aDMbUraVWyIzOoM8va3UHswBsOae9RpSd13akanHjpAlWTAADuH
ZsAavFXodDr7I+n1rgnj0O0Hzxw8ApolseoxJcms1jhADUOGw2Isrw2XSewzSGzB/XfrL/GNK1Xr
ktdx1XGh22DPEQ9e3WfHicbC/AUJfREQLOlxA6RM43cyLv+QbcAWwJKLoUlI52fU0NezGRuKcs0A
Z4PElm5LJeIgsiwZVVmraDSf+p/YU1xfFKfOi9HiumA4bPryBxXUO3hO8UtS+76DxOm2h8mDW8UW
DdDPNCS1sNbgJNHVy0VS5S4xFy32v3IWgIzIY048gpkucXbJS8aX3VdVS7W2pNOnWCFYoacQ1smg
dOo5LgWvCssUdaoOkaTSC5RrSftfmpK0xh4E0h2VhKfsBrrIJdaGBkJALXvlpFjQrja0Emw8QmfN
Zi19vWe3cDS8cvCneI1UDS5Nxs0IcyuLNq9+DhUm2yTB8aO2R3gYrylcbKukF1aYqDg6BdYNKcnW
jQX22cOY/Q1TOJao65MLIFckcCieIqIAFcfAMHcdFQg95Su8e1LfrCSMT+TGNPY+FOzVJNaWSAjf
1tzKgj9+6BRzOMzeLjA/ng8UbUpLzo8ir3hDzmLyibhuUqn0U4rGGNiXHJ1PePtg3q6JSM48CkJH
x7ou3ZMJsk3v6GUD2YEJufo4y0dw1TEtlDGUTlbQ7BhnvIZLU+qhePxeofrWGP/kMYxz7qBTTBRH
sgW0rWlIdzH8DZrF1OkoEARUwvX2O9pqW3l8ZP4+0HCm3vAK2RF1k712nNlqmdLy+cKyUFNLSVK3
qlqPFgQWv5o/pq8szCiina0oTweh6QnxWiBlWL1nze/0PyzlUCtBVb5DtefzSIeKgpF6+c3oRN26
h/4uLl8gW1k/TaQmBMV3BMzAEgUeixmv77pmteC8dVhp/QtQs1gHcFXh7tCbadv84w2nGUxgnq0e
yt3p2xrDDOpaqIa9oCjhJTP7JLb7UcWIajxgne/K1vXFdpavK551gI7qRGavfY20j6alQxB2cXdk
izsxSS2T96RQFyZTiQW7hmiyhVPyrjxygXS6kDSKxwn9Dy7JK/MehScw2NRmNj5DESkQ72YH3Hfm
gjb45UqYqipoGxjG4J7+5d2UEhRIGFKVobHsyqTEQp1Ren07x30m+Q3lJjXCHV+bqEnklqnJs2Eb
sk1cC5nuGKF184cYjGGl31nPVNwh3f0dO5ytnzM2+wAZrro1f0aXYt/t728n5tzl11Lq+AcjtVaC
sPL+GZndI+HjuUZ2YLrBIFh7YFO/NjvSIwOtIR1abNGRMLdWS8r/uzDJmagBfhAFk2ZtT1IQlPws
MS5+WIfcdt0p8MFyqtPA0cKwMcMs/ein475anSjVKpLCc1uSqcb7NA0xNRm1wvgmzIGV2jJn3xdi
tlKPG2nXnDJNjdm23iqBeLfBossYmoUdvh+3XcrJqQplQzfogjg3XeOBgFVyiIUH+ptdwcVcYtsB
OnCBzcCj9efWvQWsdPUWPioJtj4ALS6DpGROnGRj8hgaprXz031d11XHDT2Gz6digW4KnTbP1jqH
eseU3vJYZYx7UOd2O7k3zn1gzaX3T2uQVucl4uT6kdUz0FRWZtoBz23PgeHFd/Myp9Ffnjh5xcIL
hDyW5hXcktqw54KdWYhSDUQy4jCXUtnUQmJdntxfn2CsMxph+nIGCojJfRlRH0jKjPnu8R006ViL
137EWttB4vYN7i3NMYQMV/IX9bCR2UnV3yA7i6fwtfaMeT0xb93n21icaZErg2LMtl2rrYHQMm56
58/zZtcvhpRafNOtlCU/YDso5tpDMT6jkGL/AZGrAv9/4QKnmVmDYllMdx2pd5wxlziqoBAF24Ku
tyW8Pru1/KYohcKu6V5WWPJzAOXqLdCsg6tGCpPhByeyCHhkjCN3C1fMBOL4OBUMk7FndRxBpa7o
LtPM3+pk/N22Qsafhw/mJaI1DhGGkdKk/7KOIDHtdr9Zqv21NL89DkLjjprAQoN4Ng6ESIECzNRt
xM8lauCXtQEIzfp0hOBnPMFzEjdKBo6Pt3CHFQV8H7y5E5jLPMaRbMoXQGaScxhiifX9D+gzuL4z
2c/4kDA6GJWkR6L3y9kzON65sGL8VNjM14ru+tbT8ISKM8RFhi8Qe4gM7G4/SgyAntqUxNHuWYk4
cGkPzGdB4mAfZV//25FNDot7HpfgT/kBLsHqQv+zjvt0IWNUBUnSaRYENndFFklPP1OI442Lp8Vz
bMVgGNteYaoudQYCuAGOjgOlpZo/sNyMqtW+gm4UhEvvvc/pan56zdce2+eONai/ZdMj+34q4U4q
RnKZ6pSSkfcX17pK4aPMWwPcIR8hojuPtogcbAlG9C/GTev5U4Y8vNnFTjmzqwMWbKRl0yr/ZFN/
cT/Mo1VAxFe4Rt66MlmJuYJg9q220GdFfrfS43LKqlJCcVD18Oe+M6zPCZ5owaYu9518e9SrF87q
y4x1Bh1gqxq/nYdob+feG9C6kwLKSxELGdD9lUl4oDB6csxryizZnJbMfCD5Mv9PlH1/MgN6ulIE
/QCs4kr7blgSUcN4mo2ld2qNA3rMbL3Q8a7ExrFrQ1BHPrJN2EMKd4dv8i4dp/wflPEJLjMzR679
3sbRI56bB0doCEc3AbqquIUPEq0SoeH2lr/8Pa/vwNT+cv42qwEaRj68sLeIZpfCaS2FyzWorzrF
GfcWGYSSttYPOPXP61KnqlGQeMpHDaAi1Z0Iue0kdRhyU1TRuqCPRdDOEcATX5flArpSOrjWZbkQ
WBn9lVKCDHLg4UTa8Kjyl3EYEoXWyNEcMeuuAMmZqWwrpIlXC+WF5O8HzrWSk+YsHQ75CiEh0LfO
kx6CyEK1cMZeYAnl6keKB7Q15NtvvbZHdwTy/RX+i9zWOQMfA4LLGxOPupYroVFRYPF+2ysXKyK6
pnHTZFJgXWzCj28ujgir6q+c6CW3oJ5CEX81ZosdOJOy3vZ/ZOWODoL+ibS1OVquTDwu5rNf1la1
ctSZnVHwWmBBUDdHzuhkDZZbvH2IxCeQeMhxrnxZT1PUFcdFwdMfvCDAc6ufHUymmkr7mJiy9WsC
aH5EMzxaFFN9YsPa4Jf/R0/UDXBe/lKmJ+JbyxSErsiVAsBQzshy7mf71a66kzT/xELbTbDr61EJ
r2IqgugwckBR2NTeK4sJbbCe5VuOoqmvrMmd5rlYoBcyRpqHi+uairy8Qz4ZGmyaRj2f/fHETHz6
gofS95lceMzAjcKl5y1LUH1VHpWA3NUvpZmD+cjl91v83Gibzr7mSBTM3RIbwbiS/ftuKPoQHr2D
wT+dCVd7bJo7ZO715T6SbsibgeTy/bjzzaC5w8WeDcpDk0nBzrTydV/O9hCXsarjXAOEjQrEeHlU
tJ1J+pXpD8w1HKfSDYMyXSyYiDPKdkLhgFshESbSkU5GvPyQ/EcqtKghSHf+Ex7nM1dAHjyUiw3K
BWlg0IPRQbOdG1HKA8v5QQ7QCkTZ8VsrLAXtzYsGJIAK1l4dflHqXsfZxOFZM4LmY1V6IgTV14Ts
NSdMSKep++opdxqFEHD9gWu3GurWaz2jyyKQq9FdNU3WA5088d7O9bXSPkvUicTu7ybtccW6zxxt
/4LCBi7ZtTG4OxhwULr+XNHM5ry/cdoPm4v7NKJBKT0/mJzSpqozmlkSifNazL7gowOeHxxSYESE
CxiSY7YKCIT2VX8jdCvORnmPMraf2/uHgfX4VGvBGqxhqF+NuOGi2lRA++DSwIn/MitNNL8HEOPw
G4XjXiHrIxNPf/R73sgBwwyyQanbY2CLKRcX/PpzitVmwdwxzoX8BhDSaJVjrQ4Jw3T+/kNACOFN
933z7RzxQOePzlIGfeKiuuNc1HG95STlGAAgO4CmSc2X5uharzHYo6sjaeH0L5RbgnXySW4EQhLn
qqFnfWCJXi30OEaguGVcotHLsaJ+KM47F6l6APB4hDR8Q8SjrLb+cRPMJBqykHzHkLK+x6/mQ5b1
albYYMHZTzMY711eSA4Bm77dxdNxsTnNzXeI3+taZWXqN6Y5yZWmQO9sfnDbYQm2I/kqH2dFTGdi
6RoS0V1xBoGuL1Pd0Nb6NQnRvt8Cmj3nNnVGb/fmFIoS4HCZhzhfHsmJzn/W6l1inviSEA7XK4ww
oCwRGqiHPyZitLeTkO0OTse+sq99SW8hDeLFvt0mofTb+ixMK+cvMfqTqkJSXNVQneqAthMFAUzY
U3Xor752cC/B9L5+UC0qLdosiPE9x/bVEQ5La7bh0r529SNBaJiFSVm1FybiO6IVpxoHIQGyoIvG
TdwDzO8XfIZxMjXyU5E/MuJrvxmdE0kh+HaOjwmNxdkEzhm6j/ScpPQtixL6cf5V2oU9wFC6fVe4
KYq5Wqu0jDLKdO2IBAQMzJPNUN0WsMtmUYkUACtX+ktpIut9cSYoRRioph+QHbeUPzwjzk9UjEwV
gFbVeRdh2dzIgAIGR7SnV0bcl31Tpdq3x0jkEDVXB6IZIy8qB/hUpqKX6OSC3dbpkapKMvVCjajf
hUKBzY+6+kYp5434veKJ4ohC3ITpAZMOemXq3WEZQkt5wOOYC2ulmlrdbhzIbKMS8iwHCExW6GPM
KXjbJQP8A0qEjmzrCY5a7LW1ZprsR5no8v5IHjGs906FQ62/eUFIpysod9ZLbJBPhokNBf2G0biM
NoOG2+/NJyhqz4Ud0CVyCT6WLScsygUxWVs2Dcxe4iFRS6DV6UO6xVtOtLYg2p7lxi5SahSiceBl
gnGLnZmJAhZb2ZhqnJLdCNzUecRFmN7orX9eL3IuYCO0iFOZRvBOZU54c8V/9izvikLgKnmszqyX
jcgWjDWGAVnRFvQJr1MuNkzeLs335lfvwZAcv6OTVAjZ5U8JSsc30Ufvd78bVGVY3PqD4nLUDnR5
V2/Pv0OVbyV9aH3/xrRBvR3jEc2Y6mXxO3QKpIeLkbOFn0/Ydobn19e70AMAXIPpvz081TBlqz8W
sJQT0xXHW/teuYbWN1O+7TgI6EBg5LIDsv7Z2JY2zHdEa6hIpLhEC3ausf6y/k2WkP8zfZsquAA2
xZFLfbX6lFn8B4bAoWVFTc2DFJLwYZJAUZSKhZcJeIEdjEdUtN+OucNwYch64J0wq+EBbpzAWDV7
vb6GYsCIb9Y0yG6SPgdWgYGfiqX37oEo0s30TRQnZLjMUZAjUOc67bNnrmV63whAOvqNuEoGz2va
2Yn29d/20QcBAz+4svOsTEEHOaSE/CVdimDK2mnIJn7C0jlwezaFn2F7mwLzRl5IC+8jEmEs0EOo
gCl5vrPq2K5IvOkzRokTdsdx+v03q6y72IH/zLCOllqQxDed5rQeJA8SvY9ErkmvSACMDMcTtc79
Go/Ffot+2Pb4zmiK4Teinqq6gfDSE3jFtprRHiOEnY6BOL4a0S2WuXqbkvJakcowtyZnrHV41tra
PQNi8PbWpZ1iz5eswZQPKv4h6QXU1IjtvAdn7DhjvB/0FqqKE78J7ckJuOojF8q8r/DN80rgo3ew
j5AaQ2fZWofNpxxu9S6yF4uKboXCjcf1QPa0n/NSrc++1puD0wMirL1OA8ajshxDrvXieGPRhUEn
ct8ojpMulTvwwLTQgrgqO3ETzdRp46Bla9T+8JOLS/Ads85WJ0ucxrE+9EWOrsyHkT3zLQqbGAoC
1ez+xYno3Hms09B4fTAJw5QsCv86BVd8uZtYpQJrRhuUsD6eZLs20KIdKNM+qk3SI5mMnc2ghz9p
Gv6cMuHBUOiJRVTc9KukTiTvYFmkChSvFxiVdmITCazmMpITDwHy5mrzObRQPUuHqY74mVVkbzgv
EYeugazuRiXgT0Y48R3Jt6ajdZhR2uwj7F7yGHt047D432rP5s9DAGSBOeHYb1rHrtcBZ3Me42QJ
LXSsXuIK1fY2n3m3WbM1vz58izD+LmIhjXFYwGrjV0K2vbtGYyTkb8424OyxASBMvLfq5PExOXEL
CnCS0Jrco+WIyuekCALN7+XAw2YO8uxM7qgrVs35fgrpDonY1PpOSGNEl2B6R+MxTUL0vgV2xTzp
+v3jIS6VpLW9YCQ0EvH/vd5wT/pI6TtH303PXRi3AtLTaAp2GvQgz7aggzbLs7jmT44PAnIy9Og+
yKb4yDDraed67L/uIaysJPeMTRKuZgSbEC1NCDFbCsoAVYWyOZgj33sf647/6F0T92nr7ygcLRL6
aOVCpaAEAqAgSlFPJvyNOLVArsqfPamUvsmGDBnDMk5ZS04GEjltLAo62zYkq4efxm+KSphGc5+R
q8pJKPhiyTSDaUMmdBd05wzzn0tgVzi7l34BGRFVEe258w/oCFtDbmTCJbdhNm7ehqf9OVb7/W9e
HQP61Tziewr1WYuPzzWFIFn6tqgmH8ezIwxNtfhuBTLE1ZGn62GMPVqbYOOnsq57thT1rSQODDYM
xpdlg9jMGBp2iLlK3CuDvrWJcy2EmMr9EGQMwTpPo2lP1jD4W2zVTGED8wdoO8MiOs9fL/x+J+sR
xPatfpAbNQ5T1QTndy6jrvNX4RpbRRv874ynvTE5luYw1pWVFoz82RTs9n0Kor8C382WuEZDs8xJ
l8JXOkhG5DNwMrAjy0ptVTRxqC40UB36/KaFXxZfoFEBBsP2z4ic6BbEeGgbyodl7ZvfFS17aaYR
mqyoZkZXs1EOQkFeeRcpohr5IvNAouNncEVbKAFk2Ka9m9XIhmTIwsT/mV0oXCRvxcLYHrYlzuK0
85aWNAZm1YBYS3PDYqUylh+UYa2U3ONS8qmOvS/POGPc28c7bah9QI3vQ1OCDgf6lpGW0+CnRNk2
J78eNkhtEAi95ceewnM9zbuuw4hRZJwy+6Bb13BRDRpfLwfV7mt65NZbYGB5QbqdEmf983j1X+2A
fLUSdhrBctKfo6VBKyYdeIYdeKYVZsuUbSFZtTGw6ShtPHWnX2sLI7YC5Fb4GnGdrnYcaz0sJJ6I
sX7CpssCnYos7M6DKhk/c5dD3koCPh4LIT3nncn1sDveCe5cYLXxpgCkBCcAPs6AFsF4DfI0PKGN
lTlXtZRUz8bCBaz8oWwn2zVdB8btc20oKo+waHHiZXqWnsdSbc3SZOXvdVxkP5YZoYJHlnRBMkXi
Hp7MdVjOlN+cqgJnJbEzaY+fP9HrRGMag6rzS1JbvUb2qM2Guc4t1pHcO0373BBoqMUYIL+7cju5
pBSt103igc6R6zUSRFqZCneLvP8zpaIBeVW0Mmk+aUHLgR7v80T7mm1qMDupAOvQDG0q3Y+fdmW5
tOcqc8B5EqrIhyhRoxi7e7ylqVBCJD8gX+rnTBiWOY6j3aTgmWUv3GfLQGnuUWm+XFsBq/ROIhS2
YYRwydjG47zD6nseo6GMXKJgrz4E0zo/jpaIgWkb5muXi/lteDHAajX0zOenL6dLMU9xbVVqQ2JJ
fLdzZywI/hkOJlwMdmFbIzmdT54c0jDw85ap/8Ef3nSTu/UzdAMsT3Lw+JQ1r5WsUurriyDgh8W0
kPJI9ABDneJEVd3d+moS1bEyrTD3LEvZ7haYhvz34mVc4sF/eivpQMmCTQU6eHYCaTIBhIuHa42d
SsTbjFDIyoccZpdhF6Zw3WOScYRXWYZ+qHHrxWmMNe3PoINgOnX8fpxwY9DrFOmQ/E882aHtlikr
4tqgiuW0udjnvLyqiGc36NRz2aNuALts+UhnbAINZsUgE8YJWvWUJaMBMLsrGnieY71IOYPshz0F
FCDP7rXE0FLFuuTRMwIF3qm40Zg04mPfuLoVVdt4NNrfSitJjK+coO+vrtFTHQgVUK8hNMB6OuFG
Cp7cjCdNAFs2nehSu3mvC0dVoH0HidDEG+XllSVDCf5ffyYwtyDFg6WYexih9sRDKeS82upZepL4
y5jltUyIlXgnTGaH4XoyLMJl65IMfmVl/MQ8D4m3acpPh8rN5B+PhDMqONrN7NzGM+iwO+9H6SXu
ByjaAet22wus5PcYCykJPQ1aTuarFemIIuF4KZ4DpnPSP+e3QyiRd9QpKEsXd4lhKZcrP4Lzl9vp
CS4Ela/4gSvr/aZWlUfGuo4N5nGGrzepyMQw58LrBe7WZg6qlfGk8OsRkqDuxiv3WOgV87U8wEZc
PgeIbrcs8MlJkznZ2GV2z4jNhHTS18EizTjgzpQBnCotOp7HnKxFc4j4BSONq8Z/kW9UFdZfz/e9
2ofgonzEmKNFGGIwI495wj5Zdy6eeTF8wrKN3p7tIQcS+HedbQZzugWYjDRP0zs2R2T4ChTjCpeh
8meyMHJ0t3MnSWzVkICf8jNo8SZu6+N39q4ItVbqv72itZYxGDWLzcipwMifsdqUKeHsaozPaN/D
4sFoqfCqg0bkfS/BeV6ileWCgAoiI00TMF2n870MXMn+CmazmMSnc9/sAPmvw4YUneKbtqp1HUE0
3+2iynsU4m3qnLVXUC6/YCCrRkPie5/MvTuDYLrlfpONX6qdwKAnSJ5j9cqLNwbeDrk+wsqVKMYx
+mSyIcS3o6SOX4N0FLKDwBuUxG8lSxbrQQaY9dUeGITRmwNLmAXfsEEt31H01yN4PqJVqce9Y8HJ
ccEuCpBt1pGySvpgqEzZhFR6wBP71BSKHKArIbEp0NrL1tB8cryQsIqvenx8r0DkWF3QgZzol8p7
3tcS6KRwpkhTctKXqyPA1Pe7W5UrXYB6eCaxl/SYvoumy5JXqWu/Ydnsag9yEWgtT7EhfVrKlEPP
mX/SXbgxXIW43M8ejS4K0fiU3rFt8HZOGkbM8cdQUB7stRBv8Rh7gM+v+9AwnbIHGh+GTi5Crzib
UW180GMk5ekfaSHrP8UDiYa9/CFmHd9kD3h1rKValJJBNsfaaYzTTS9jpNhgrW3Wlhd90DPtbmuc
dZwc5tBpstMXvtSqbANAYpKeCGzLRYrg9oL54aHO701U6z7F1G3RE1pzH6X2GOHovR3UylSC2I7k
FuwiNLdIDngdHrOXO94lgoYQTjBQxuqUIFpMXGAX5nNyvP90onJKKZ5bmgmI/wyyhbcLeU/gvgge
7k8QSH6YZ5BDuzmDfLQ8LgGLIJTQGgMAmfssVYhxwqE4bIj2DtBkmaktcLQlZjN/7ko5hdjcZgz2
eHMIoa4l43vIaiwUnSxbJBj8ty8ECr765K/s4ZmZlIeVS7De69NLsbz5Jv9zQAeFB1+ea4tH3hU2
n1xTTs+k0m/aw+Txc5pE4X9oe95WGMTq8O11VB8mPwUHFdmv/R0jma919+CPX/UCDrfU3Luwoo2P
0nGYT9DZsGrRtZi+1bynSuF7gvl10HGCUYVXyQguN1SRpTxD9X3gDVzllX3tl1xeDbdGyHK9mxpv
EACnGP4P/YS1+pwvkdfuY4PhKg249DVVfw+eo7qiBEhlxl2n6g+dNNo7Aob/nt96BO6aiDT7F8TK
OdRxfnHijB9h92+d84XUoe6Gr9yp3gEsweCUW5KdrDsCkuu8bNNN7wkKeJedvyfDowW/vl6EmxqN
4IMuPKGsV4tEpoGsorNrW7Qu76BRMrLXkloh9iF86NFJpp7rVXklwLS0LyK/KKtXqNDmvESqTynv
7BdNP/M4WbNjn5AtlxngW/bdVtoCYncv95iAtcwR/RvpWJqf7PY9v14iboqesrSUTCL/fq+0Sv7U
CtwwRFtzTVF6cxMqSqACoGhAbsfTbRZxGIJw9jSqJIeoMWauckI9csdDWNduBd1qR66a38vs9dmm
M18gsvMi6uCKryuXfILOmFcEHAiPrEcMsA8v3PrOL43gtvi17+v3VY/O6sfX53/VcVQCITV5xzbm
TwbJLPQB797qm72jFxpSOE73oI9eBtwMc/y6Q8hrkf+9020uZQbcIu2yv/9MTDxHbI1Tvb9Oedg7
7EP8g4rDiFe0OnuLck+AKxbybWlmOJM1v4u3vgFjmSXZK2rTBll4i3P/8nHzAfap8lYC9Gib4VV9
ohDHQGgDVuN5gNK/5hEcnY2drxHDYsWziYDLgqExkuF+Bfc0pD5ZKqoQ34RaB/e/HJQ1TXXQ88EU
xh8bMpECAIryBOqwXbZd0wW1S3d9riR4Mbl1Am9dQ3Ygn6YvPVu2kb2XtZqnuvURGGs+nm8i90se
9s6F+uFKyIxC1dx9SNO6CvKTp0oa8cZGLUHRYCwW+KEDner70b2DiJMIe1tFHSNJtCWxdt/p9pzK
Wv3EQIcd3OPnzkJ20NIVO5USFCtnRqKgFYfSksG4BNaVauRoaYhz7xEEaio6opxcjb/t/AqvZyEl
00umt2+c5CGRERnGSpK4hhZsJYor+PWdqJ2PQJOHzyHcjJ1cSpt6o/AXyPSjbhBUFpRhL+6/G7cm
VIbXtQB2U/MDBjaEqsSBEmStRLK1B5hTldPD/KO92Gc5xTZ/6GeqkmaW+VOrCT/yOhSdp+TrVXmb
9lCjQAGVOoaVI1t3f538xbCYeDTm5su194ScD4SF4CgBOoUm5qLFhHf49pvD/7Fvp2xWpfK+L1C0
5jmMGbpqRk6w3nctMVqz4VzIsrnnHjYOkF/FONFHhjwbkqNE2vwrPQYDhG5ZBVMSExu0A8nc9EBH
7nf9V4JGYh/hKnVxEo7MUFTiWzF6xWPcm8eYCSPDGJsVAa/ggvafN48VbXmZoRNlYoJcnsbSDQ5h
M952YpC3IRilA1KnGQOB+fWauIsklJF4P7pBzsIwxNKZDCps9Zj2BcwZx3uEw5xvAX+lce4IS2nC
rabTEBZiTWKkO/fl5PyEa2g3tOemztL6BVK5JS1k70poYvU8uyOgFK5loQ68ggW70slwTt22HT16
BvdF0uoASoSy76oO2C8R4w7VJCC7lEUv9oMsXdtoflE5F1dqsY3mzvTxl9ljbFtpDRCdFkOt3wRG
MxRfVbR3qjDs2ElRsU1QWDeRZuPH34xozjC8bDmDc61cZOr0kbT/+72BFdCupY5oeUyVl8KiE4yd
66R6HIBXsIs2EmnRh9DyK3pfeAb/7UjFscg+JNFp0J5n4eyU+ToXsQkHhZqy2Cir/H75Q5K3Dyxx
zIVZIrzmaI6K2rInSc4SS0jpQwpEpQnFKc4lhUnK2jcWz4lH+47NCiYFC3OQzpfNOzyV/kZVLIfV
89lJ8xIScPx5RCL60QvB91JU7i157s+oVnWKVoLv6aZHgxi6+060eFjdLrEz1rMIH8Qb94Pg5fs6
aKEpQ0hDFvuE3kvGhWGtRIthZgB9jw2DFDdhQrIdx8ryj+IO3I17Zrg1WbgRFq6JCeeANwEPydzl
S+xFXqinXFg3brjnqyaWKp+3LQP7K2pVsPM3GyiH3rf0Z0mx/Tt+imnkws20F9FBJmpHFRGyLe4E
YdXMG2eG1mu6A0AxXxDiTvm+3JCtVQZ0MWLJJiTm2DSdWv3UJYjqH4zqNZveJ3+NM58XqeyuI7iu
hlQEDkUAPPQyZrfBF3OiSUDVO+kZ9YkpdcVmhpiCGjq0OcCxMWze5LoGTl0UzN1tUUKqaTl3Qd0y
uHYOk8BMWXGgajTA53PzxkRyLZbI0Xo38T6tfQPDivpjvyQhvN2lCJhSHVIB7nsacUvaEd0TLlVk
xKIpg+vhPF4lcRPPagkP3vEffgMs1KrODyOMEYmMKDXB7inc8fsgGtjd6qd9W5qA1TQ5rfVOgZvr
7HDzE4AeoaTE47TVocNXtBHef102D6Ldf4PPuYb4/NHCW3QbM0rvjatSfNDI7UGh7NPDjjqqbSBs
5D7PqXZkTP2MN+7UegYxyNJfvxecDIHkxTVD5g23+RJDAAd/rJN8qtl14W5kAekPQh6iH5LVdLzb
jIJ97IOZ/VGkBR34QQFfumhgDQtfVZuGL698OqqhHrz7osie02A2zbtF9C/NHm0Njb2LLNDiSxPB
G1wvuqRR2PtxO2bKLuXmu1T2e6VGEr1zKVQbU983JK5LZ0KVDPYwCXDRr/R1RY1R568xhfqoxTwR
SsIdgdnn6k82sdDSLzgwygsJJXw4WVQxXEqM8y/zIDEGItUnQNneuWAS7zZ/z301DsMPDGvIV02W
eb+O524wPOU2Cw1DDalHPbC8B/Z9Sv0DRVSBcHKCEMasfbuWkVftPd4wZ2Kpgr5tcpP+heYKlyS2
bNSSjoeAJGMVZUZY3u32Es5HpbfALGBPAM3iHvA75n9lEoH6X9vdq4+UsmTjVgkUymTND6QMvE0Y
tCer2qTuJDMffkl8ysjgaPKftJpbfAnbP6STan1D56AAomeuc75JsQUBF/t9Cw0WkHOnp6YQtwSG
oWiEmkw1IwxaYK140gRMpiOv6LSbXfFxmoTvQh2xGvvwI/UZMKzogEooNPghbTCnVXPCxTiZ6EkV
Bvd2LamLViCcuApNooc7ykutTUqq/UGRAqm8jJHlfg9GevkVk46h2wLQ+sguUdzNWNjGq5MfjGGY
KIhIAvCRXfiWEWOZnkSG77tV7iPySuxdQDdYVLxqoJQAVlVlIR7n9+iaLSo4Qf7QCBvPlU9bDo3S
h1iCLvy9Trr2R4kvqRmpvwM7ToO5yeGywJG9bm9LtLtrw6sqPBaMG2Maz+bmRJvKIAqibGqrqb6S
tv1EKa1AQnYxClxuqM2ky4pwzfOE5qEs44U/LS9bNIgwwml5iTDbbJlNz/w1UAchq9AJ0I96RU27
QXTmzbUVFPaynd52l9e/7CELWM5tS6+JvL/RYK9/PU/p80RhgE3rWkAM/SEBz7tOWZOZZHqZc6BS
Hp2ifblxUc4Z1r/s6+V9vN069zwZ4CKnK7V12+Rq0IdbjAGz2REB0Uv3Ekv5nVoQ1A9Ux789Krcu
H7UxfqAF5a7iFTVTK2JbXP+Ju4OyKza3RzblWiw3HVCvvV2YbdKPVg8kkBvnJbsOp+cOj+DjSnUy
n5VliYQuke+rTut/USC6FIM48FvlsZWChAgEwpXvQ3PeUGnuECPkafShxNJ0tvPSN9zq8e3cWVLq
SmaXhLjGIdKwl53BkFMiMoqP6UiQdzUjNbJ0abqhTMbqDTUUoubLyAYb8fhdNH2jN7N0WAatq5H6
a7pvdS/HcMjCw5RJ5O1EcMEPQ9P4afIbrN9BklN5YZiK4BnS6fhFNaLotMEtNm3etOCsKMlnn2qA
rzjEJDGSbFblSjCWFdNm2CxVmy/7+bkYeW9PvfOhPVgQ7EKYF3KGnKLtt60CKLLp23o7ZffWe4eu
1D1TaR80ohh7rLVLEKonYxcb7bA2iQP5rXwf3LrqlWE872pzk8lmF0MTjI6pCY1DhRwXCdEEtRgt
HZDMGd1b408WNROjACONefmbP8fL/8NhEqZLT0h6vb9BxJOhQOg+dAsaIdwAK0/raGCC3KJypZSW
h90L8sbYFRZ/87RUYBDetn1ZXUmt+e5mvBh8rNOTNcD6r4Gcb/xxbmMakl22rgDPYYkn1uln/Nqp
avgv2szYQ8TEztrz2qvtOqPzJsp+he3DMHEfZ2/KpW8w2jFibeYzgWt3ZdNJbWUN/FVXwMm4DrdF
SJ6/VYmR148jBBdYDAOo9j14B4Qi64BvXY+awUH4WaxK45xFAXDVY9x2esEjL1jd/Jy+NL8gszFp
BvvtSqIvirFBsrgM9sQQytG8u/Z8+McpFy16OkmA49mWmDJdlI2q9L68OYNbr0+SJ8iGV1nY9JWA
srlrJZXoUAkYaJFye+iu9HGuNPcJxiZNFOqt8pZvxX62JMmVFsFNS2uXvq9jzCFfn9KLx1RNBlDX
E1AaWrSbY1gOZlOXH2B+l0JW/cF6nTjtY8vv9dSIaC5sP5Kh9zB/qPZm/gJUsDtWycpFPc7PcwRz
0hlyz1qFts1x+HHGSqUUkEuED0hFIlFQz5iZm+5vN7xZIiGGVM77i/Ig3Sp9YbX7y44MhlDX3t8X
zFhwXVn5zruohSgmg1/LEVrP6jvSHPMssWaQrnq0f1ATU7uzVlkyCgbUz48nmh/IS4AQYFiSJM5T
EDzBiYFd9RgbJvywBN/8tSgN5nz+sO5c3Rjr+cxi2l/teYu6qJtRoczchm4203SPF/q1I6WJuPkE
5zhWzF8WwpOKkQLe3YNhCOUigUa1KWlJ2se7aYh8/eTI9kyvjDSsvjUmMNw/ecO8m8hm0/gRxMvB
2r7WJj2OfEJQ+3PsrFaQNFT7FjBiGD3KB6zWoYcCmiDUTG0fYOiB9JzSLF4hrsYzGs/FsrdXUlz5
QsJPad+iofQRPszEg5yJ9+Uj+/rG2iABzs8HX/37cbhx8IMrj+68n/c1TMQSOe7F70eM/ia9Ddak
ze45CXhhzW9cWM73hpGyfOk89F0kJVEt6luAvMQDwBzr7XOvV4vgfug1KYika+CKNjWboR47uPjR
X/xp2bT0jpG+y7DBpTPBSaobbHwBnWs4SMhxo+aFAiosF2ItblvwgdFDCZr3JlaSkkLCt5EBkVNp
sOEPnmiQVyUFlumK60DyZw/LpRGPGC2lQWv4zND5KpDSIU1SyTB1lUZIePaWqZvKsNhyNDXQK23g
c3wMMA0794MUT1E4co/myKE7KKVjrTuOZmwICEPz1n3cbPlPewy9SixU6vGwk8DJlrtxZoav2jfM
EwNNJxWKIaMlrW+/VbZkACXQy/ZJLvKeRxn2fhYyvq1cpUEwJHjPpfFPeo9OMid/Gj4eqiAPvTuv
VP/qsgRB8jn5+XKxGN0YEHQumtwRBEj708Wr2R8fiAmnUEXtJnpW5zisPekBCnsThje0lVuvOw/h
p/3dM+UqSuA38mDbN4kiNOIwaBVaB0eRxm2ZEBjya1B+4AZXnO6PwP3HRR8uT+bNMPqEwDKB+qci
BTSqvjxzdVeIkb9Fcr2qxm4fVZeD7vvuC+LSKOgNrrDRLmH1xDbFL+SApXfNjF5mv8F0nZmThwrG
tMsJiRmeqvXEvSvFxeIwQ20L/e7YpMkxi4PGaEjYyzhevXFYQ3/lNosV+EDh+2vA83dAuD/+HW7y
rG9W4LIOHhLCOvV5sFU/jZDK4mMjQEDHgRlat1049A7QIFZxxyEBBu6za3/371+0EpyuJ6IdQ9wS
K6ke8IUuU8Ku+GGkcOVtsRdZPLpLwRKFbpwCng67q0ccTdiQdqmUq6lyjnara3YeQJ1412kPOUei
vsJTu+W+jDkWf52w+RMQLC4cNPQ5rPWo1PUf4QeEenRZ/BjkPWTjOr7NG+3uIJz8+CWnd/i3q9hJ
W5Z4m6T1w4D2qOP/UJvHWWLc9ykrptIxvN1X0CqAYmc/+Uwf8iwNGBCK5ZP50702FSSY0v6BU2cP
yERMrntJUpQSiYMcSVqtKHysocviPT+PGSDwDSQClvPxIoAfOW3ijm6pk3qNtOgsLks1MhVYDXDS
IkIn+EQ/bZFckjA9TwV2qMw3+hGGKC4rUhmAuT+V5eQnOD7MaOleEsjeDI2bh1W1kr94ePFTToiJ
5hvagao2MoU/5UNO/Kq6mA3PogVJRRkVkc9bn9t5i1FgnhvQwAA+KtjDuqSHikYH5io2hPXlA6AP
UIEVDkxAEehC9zpFeXnUBV495nSz9zSI7SXv6i8sfAd2jHRBLDJST62Kbv+4xLzbr7m6flyWotTV
N3YqNN00t2Y1+MEO7RGks4BvgV16kc3q2SJhaminZOzGwvzScU9EjkZsEIKpQMfD3fO2rTb2Ult6
nUjgrgblK6X0xpOU2FH31Z5QLUe3r3DvjXirvjxKecYpZF0tJtowgs0aMqkzRtJ6PYR4uzCbxvQa
MRHLaBvkz7hL669iCe2AeouQEFEaqsV0EsuBAI879N0XQqoJaE9ms8UgiZ0LdjVWUjiIcNSVBBMx
Ml43VXm6qxb6LSHuSbBIRIgFUD+uJ0L0GcTIP0yL+uUDlHFZavNSs18LAPOJT7bqLsTrkhe9aMgS
dk0/sRpIUxMFX5kdF74ue86TyAH/XvIY/gAsHKVbRENNHzD6sjBEg5VEC2o0EVD/l9GwDludlRGq
YY8qt9TUbWFhZY5gGJII3B+es1xqlmQkgmtwo+dD2O2V+97RrVIqnq7d08nJcIZpa5mp+b4g+TSj
skGH2YhDGNE4uZnfYD0P0skNMoxhZxb/LnJKw9JOebCPl95wnZT3LVD77Afxtqteq2SyWcAoQhag
gIKuO21VAsX3dQfzf6Nc6eMIX2IQupwDkdbZ/O9J69vwxjMUgigxBmePYmE2rCjgpq5tQBnNmnBR
54/IHVf6M0sdgvTmZplhlO1Uy0ROo+IecHJi3xb3mR4hhS0nL+UJf7ug8bhTpq+cB/bk8QdzU7FW
KowOTxaZj/PHxaAwiL82v+Qjn+Ll9WEreVSGEqvWNKNwKsjJXEUo2+rf8nJ/XQ4vSVJ4Z4lbFhpi
hQsjnvF4OhJQmwDAl55jac+0p+HuTyb2snM9fRhS31TwiHtmqvnCGlr/IjtPQ3jfmHSMfLJBXkXZ
VOFPadi50IeAQ94ZrZX0621QXURVw10sEZtnTuaj66U5CtcecxfMvwRHLY8Yp3ODNAxO0LzZGYw5
kyTBmJWAWS6SLQhlgvS3MA1QnptUJKVmMM+lSHn5giYlbSowiGf0vzpRifF6ZK5y7Iu9wUO/UHst
97HwtgnFRgFzfjxR8VdsdeZR5lNp+JjXjXRBHGUwYOrJevmHeGyBRNeyUe+iihuCei/VxUyzcGC6
kMYHreM9QWvRQgqTyKbS/vU87PjZ4XYmxwWbx/NvbOfOpJdYwqlmBhhDFhqUXMRLntvgORHrkczI
cvajtYF7a1W1bK18tIw/T75Y2+QDNddoMNKGIfCb3g2MZiOQiESXD21dTtynKXZQ0K9xV3qVTcmf
4wV/1zcNl5OFbs1Sexq52wAo8eg38DYAdatOZtkCyns+Z5TUj1ZOEPo1t8+h97MJz6d85NzQUbgG
5WcyOQou9W3TwgE8Ugwuk0t6SbOialaJSwFdtJDbTKeJ2zWCvNCnfKF1Us1g9rS+djdm0RW1WlFc
iztCqBoKMULjPK2JhzZ+b2M2xNIvMmZYhEA/Ji82nHWL/rOxS5jowsDfuG3PIGQqqqJ7XrvvOa9Z
hmDTzI7Jzlaa9Ss3us2c0UhO+zNVG23iVvV0i8RVaSo8BpDOCNuoSkZyqkkMwVF5bnbSTSa+Bklt
fk89SUkq7COyhD5jwalsjtvGOPfKK04SPzim7kVpdcs8G/foN8cTseijROWL6UkapWY7Oz6arVdp
ps3m6IwcOEEJEYaj0JS9YwhjxPcKzKOhkHh0hjaEUe2FAYxT+pY59B6JJo3W976ytFgbdCMkdYg4
N4wzfRF2msgdsoXOm7ZPdHTRLX66o2d9XiPLxm6sHRu1Z3vTMMn3jc9rTYenPcKO0fOsYZPy5n0d
HS3cavRVM+/poH7Tqalms0UWT1e+Xn0GGlbU3awpNg2YtMFPCLANqynA67YQhRhCmkveTQUwJ2Yy
zYCknY2YUe+uKo/YBPqjFa8OJvEJet7aJqbnXam5fNA0PdUegUTd11L1RYb/8t8gi06Pu9JRI6Yh
MZMpSqAuKRIgAr4yuit5UcIqqx3MWa03w16gBWrQ1SWjAUHD+U/PzzL9DLcj0DzJ81cflssEUETs
M5FCQyokC3sg0JPfh0B8oQmD8YXH5NAE7ip0rjnu6Sb8ojYOEoL7Tnv+UFtYNjUcYzvvsJghfiEQ
o5RhEfNRcSai/rQdaiea2JvdfMCNvZdrbJknY33jMtdu/RCDt/sJ2qe7/4yToVURxk6rOVcfU/jS
a+Me/vdKDHe/zH0hCpUtDVQKEAJGvrUslVR5MEyX3vCcDCpq18tJ8ahvN9GuMmarsWooHWtVmV7S
dbeoziAZpDK6lkym1Dazf+L/i+JKPY51uOIuos19QpmPQhTqFj42Qk5JiHqt8aWvsUkpOlGYxgKo
XJiBfhCsKG28q2+CkdOkaCsAky3X6Dokb0xfxMhq0RfGeLpcdxHQ6q9N0mHbN1QaaNTWshqe1F43
tr+QTjON3LT2rLGzOkzOwlg6eovEfFxgUBBWtHVZlGxXr2lghnXDKCDh77pMd5JacwdDXL0eUZHf
FDj05WTmhNu5ybc/g6fCHuWWBfaQMeb7AH1+GBO+bPABVFOVXGWGsTj/GruUV50uHzsLLS2Fkrxg
wdUQFvmqOJy23laOjELkKI/50eHu1RaroBbL9EQWnO+tPt8ivpYDzsE+JYNFRj8+tsqnhLUSTG+J
odnU1H2ftraXBz+/VK4Xnca4WXtgjqgEMMEKWpmwfwwayvnip7lBYh5AqGIlxmBSApCgxHoE1Lvw
b01rnK3/abpYxbKvOkRLZJd2Ta0Bv4cicxMF3PzMK+qKQFqjdA6XyllGYF7OGBfLpttQtEx72HUN
fzq5OHQz1hJgdiDEn7alorAl2wawYBYBkLiQb4DjyNBVkbzeoDTx9SDH5DhKyg1MTcrg1N8Hy/Wl
pMFcWMOK06D2nQqEoWvKNR4TjPLrLMIPof2hAFS0SUoCwczB7ey6aTKS6RTne0tAbuJVDPUWcooS
dbaBUrHdJsfwF8PkCC0S/kVBG6CsGFhNR7trq70b1N3WzJZe9AKisFwFp/dPiKKR1vF1HzPNhFGW
sQp3G8RTSis5rGnfUJ5fF+PRKRqsSUR7awhOLu8cdpk9++zzGyVOjmXL/XyDP/1/bAmK4FSAM0hF
mirdlupj0U+8oCN2GEWZf2H+IHW+O5CRdZS27ACQ6ysjXsGpcj3Rx5TzI8stP55Eyz7l4vCHGkwl
rON2kzq5jv71OcEtYRVqklqlbQFFOygY7mTqtNOpYxf0KZ0w+SeDvB/dHp+gyjaFk0BbCjf/sD4Z
s9bmFY1KkvLVHCeAkvL/9u+ZmGkbit8IB7e9wMe5BuhnTQp/4bYy9e+h7H8F4UwfKOebDTlp9mJi
+ehthrveK6XeLgepTT/GHsWTiQlzz2r86905ybEaXN0r+EQtqaTCs614EgdPcN1EtRTPbpndsMzn
JCU5jCW05sFB47CHjKH/IrJNGe82cRtTnVGduCHxAUtyLDcODKysMIBI/i9BKOdcaeQX3NFbdIX4
B3+G/nkLmtswcOnrfIflxn2rkmi+mIRJkcpyJcgKCGRYjYV7hOmy5ZgBKrFP3fceGWPiuYGwFPQr
bunBBUZeJ6DRPwvci3TFLOn26Yhx4Jc16OReZtNBbT4bWvvnSkeJh/Q3KPh9Q4JTJXLg9ttBX9sM
8QSOy5a0YhbDpDprd5xziIiTK+CQ2GbtbW7pLZ0Kup7/ojnhFhaDneCXlMXbIo+uJ3i6SQ7ZQedg
Iuddiv8XpCQkLggElCfCuiFkFEVgaIEhvMju6KJXFe2suluWDtmraD9NYIuTwTNJOAsO7Lv0Yl7O
NycRqMDmvT9OGZrdO+I1lU7niXRg6HAASqgFN7zKBl38FckwedC2rGi8JhISH/flpt/2vxewHydP
JCI6PwtU/OrFuxaUquJdxZEFDCTlDyYdZArbPpsbsbEnpeRW1jgrBK3ajZ20039JBCOZyNamTVVT
RmwhmCdbS10bMPOSKwg6MjYEJrFxJwh/2q9ucINv8KpKODi8+GBdglFwWqDDAzGyg2deZL1ZLTUp
+JG45EDopYFOG89b/cCTovd/6k866P4BLbbAE1EXML/KL0o30+4mMDfaDFxeL5ZRQFJ2d5yoGqtq
6CsPIyX644j8zT2WelR8GyW4rwUht9CmV41ZKK+yNsb+0vNvF3OltBTxPmrGbR9w9R6xaOfTSSvK
R8u8sNLiySJSyrK1s4t4RJ4irZf5pV/KXD7SeOUPqrVjFuVDVZ3REESNRndFiY4hUcpk/3cP/hOk
cZ4NHMn11Mhk5b1GKKXW2Rv/WHyyx5KgsSqN9qumu+RAAPO+626/++g/Xi+Gj40nQz63uvTKGEZ1
6dIiO+rJVFJzKZmWwE1uxsmA4bBkawR+QHCVF5LXShDOSSapkYp9HAsTchPeWZboGTEh9E4NcmIH
+Sa2PIThPxUTnBhNL29eo3z5Fw0uieAIAlSk9HhLS9N7FfwKwCLKS5Atl6/5l3lbtz2BGeRzhHDK
P37wbocuzeB6EgPvOHomJaAsWlKU64Ow46LP/u22rgKN0YyvienFoNxtUo8pv3TD7XzDYNLi0kwB
euYXIkzRDdkSygFwd+eMqutOzsg4kH3GLYcg1UaLts1PkLeh1AFppStFGjZKD9xCmxlPDKJ+L4vm
BenK/sZHgDX+7dIoBmoVOJ1dgF3j/tOGtCp22uvuwfEjz/Y0r0vQIeR+jVAwDkHclip+9M18EgQB
DkZlImYabok1hyNzMxtnYS0EohRGEncv5CA7x7VaW4b0gHuzMWTNu5ba1NbaqT8Wb2PO0YpwwSHx
XJRVeUhUssmtUY6i8Eq/CBHnQfjNxNbzIuOIbiRlww9PGk9k1pE4l3pSi2gV7pYs218+ISDlih+K
MQjYY3hP2bbwbnOxAIFGQe9rJEJhsykJGJMKuGUWJkJ5g31uA/XL16KDmw3PGWHLK7TgnrPIQRxP
/auMluGRxguj9TyBObMuZCVGcWtLQ3iNnHeZrJAJTbnE+onH9YZDELuwX2MH0AbdBj10zrF+xFkA
tkGc4dj26jP+SkKsS+jHa1AT8PCaaga3DnT/9R3YxpP65OftoCDOZHOisjyWud4MPmRE0UqFdBRD
IW37KoI4BEt2g9zczBRYsTnR3Yy0Jx2g4UoF7vuT8jNv7RNF1mcbJenQYqOrUnX6zupZlxO9puZW
2gAz3Yme77v4ZfHVC9CpZ7FKi9lYqPR9d1U2OEM+CCqbUUPMdnw63yHZ8tatCYl4Cu7JP8U0+7Iu
jENl90Y0hiWUiqnHbFCiNOmoLS4pDmivxhVyO0JnEgahUCDt0cXKqDJPwY1CC9hq5y7jreDrzSEK
KLRsmPXpq2/xmf393QvwAQSkBAvMF7QJOdbJOxFzBGcpsr2GjV8EbbO5O54Mw/MUFIPALWjj2ZxT
PMY3YDCJQFXTiwUTeT18beiauYJX2flgQl1RHx/511FIxtz+7Uf4cfhZVBzXqyfxhQ3lsiDlg758
dhv+iqpOMvOHQ+PPFJRaZDboceCZq/6DRbeBvYmfrVaY6APp/ySV3+4OI4dafk7h9Ni/t1gZaf8p
kyClFG4DdjMOe2hLbDExay9oyiaq65iMOZ8ZsfeF+Qs75JQoX2l73PsXvXUZ0dSrJZNerjpgEwQx
jbB6NJo3oLSOYDFzQFAupuNuCc9AZ9wDpmJ5yOz5w4QBkoJQPXWSdbuGIdekHhTEzIZ7fqipjqGC
79nmD/AjZ6I8eCF7LGUHA/Ygb70Msne+TaKOMzUrHheftDCd0KKA47jm6zQrltvyB1u0FPZN4UZQ
Kz474+cu0NP7zY9qgoXVaz+enHk9Pk9bkQ6t1k3kKXOqE1T2zmKqsdvDPhs3mcWUOuVHfzRFSaQm
2XHBXoNIov3fmDnPp+CTLhveCGjbc+CGsXdAnucu7zYQcV0sBlgbB+UXNrUevHLKpCkn3/SrLy6j
3aNQC96jSCL8VcGBFOLLbxFKbf9aJM74roGfJso1XItwfHkV8WJ20SMdEfMOhWt8B8h+MZwq86dd
xtNFRXzTPF2Hhty0MVblNmDa5CIGAaIwmpGjMugk5tQE87EAyzs6W6TLSVokBTJ+XsZcQp2gmnQX
xj7rxzL+aNdLsSY0Kcl4PJkSL6dtC1nTA8Pi8BZ9ixn9/UoWcYYHqYa5yPI7/GR8CjuyavFV0B6P
JdEInmlNLsFeMW5dGxeJ0j3zn2mofQCFbEk33+DP8MvhtZdDD+0CUo2acfKJdB+smMzEyjlayyj2
ElTEDSRo9x5g9pbrq7i4/3y0JVq/+g41qEE6emBQ1HCWrSCMTpDB9Cjq0rJOztHRvdMafLshIeNn
K9fQYFEeKxszOGGoZitDHd5EV0XAEhJJA4unvbt8TfVp+g1RNyKqfGl98ye8V1Y7Yhz4MQYNZ/x+
9NzQDreQPmafNUpzYBYyyzTkhgbzaRRxLSRm7JX8JGWKWwZPEHOzilwK40w1nQXJe8tdG3hvvc0c
3zo6xqNUUjyDMY+r8JY+yukZ4T2OfHhO6965a9kKSz1DfivlIrGusvtxxuTtSjhFK81nbts+GGUU
uaBOcgJb756nYripxkZtKE2LCmAd0MC2v6Q88x2omkAnIzHTMLoe4w6/PUhRpsjASQrZp7hJs61H
ZWPSncUGZs4HUhrh8ah8R46lOp1tsNgBZMdux4ziFHKY8T2BDeIhsVCmgeXMB8BZQwggMRyOAR2B
/Or74j3hpR9jKjKIyGIg4AWEWIURpqsOO6lexWAyZw4Y7UPvBl0aqSoth5Iweu6cH9oUWpsJjEsW
6EdM3RA6o49hMzjkFoQBEKDZa/n1kwZK0CX8e0Aya0dr2uoTCXxVIBZ2tSNGC+ag7oetzmdQZC7l
gECYy3Qf89bYlL0Tq3xTWiiHxYXzjCZPpeDnGV6/s88i7LxrUSx7W1UxvO3Zyi0qUBTthVWWZO5x
RuiO7aLRgzLRc3T+yPLmUmkz0vZ1Q3ILNI0Ud0gcO4+NdQURyY4DXQpawz6oiaH3kx9KHN1zuZ8o
E2tfiKiAimEvu6nVvmfdgKZEaZWBbYpVc+4MUocgkTx82gFvEdpx8Yips1yAYKOYHVY3qhzQJDou
94fiCBZMEW5IJGhx7UMC/2HrLQuucM25OxLSBCWtOiej9z56FYxqoDRw/giG2kwdOi6z6bhzlsBh
bVpV8ri9vUW2KNKkWdFYW9NBA1D0ooM9mJtZFKITo6/O3p4FyNCrwbuIlWq3D+ZwOKdXF5X1T5Ll
fSAQjZCi4gjk7U1QpoyaC+eNmGJAJB07Y8eSWSXpqMcZcFd2j4FPe53+LiHhYuX+GwObXjGIdl5D
nbQRy8w/pSxrBWJLqLK0EB2wl1ReiLqqRTBIl50NEXghqJ3j0v3VOfPCL1X+1GC24ess6cyWYffw
ZaPPD8nDnbcRoQfEmwu1rL3v3A8/wE0fvglslxhWmxOL4Wfzn0ju5rHzMCHeGFTVGen9I2f24E8P
WVNA7GJ8Jo7FBoCUdPW9ilMsr1D7PbGExJr8TuHp5Kny/mrXzcsbRKlJEGVNv6rQKJ1/YnkGpneZ
fDIYto0NuyQmjPChngFjbuPdirpaE3nhAgJfaYCAt52qtiPAaqAh9pTWkPVGwWoFJ7hBUxkAob36
Exm8bgwDjIULA+sPkRI60+Ce7HD2Z8Vb3OvAA7wWMWG3mW39hUTQnTR32T6ALfUsXk6ibyyVxGId
R6GhuZ+AM7bHebSvT5fAHmsNQHk9BAcDIae2GdO6Mqe7n28mEY2rVpenY7V56p140A4DK3sweLm9
GYtVPsjcDhyBlPBAu4DRw0/ypiPHfCrgtAz5GAFJDWL3+RaLh20iGCMrQSVchxO3T39Rs0UxIVTu
V8WoPchOQFb2GJ5oWPRWpHO0yxLNUjW7LarLKq+OGN9ssCXrw/fAaffHoZ3hW3yMlLzDYNVpX718
DnczN7XJTGCr37vh8Gbs8VpIdH9mfdUcJ2RJrbRXNupvmMThVZ5xPO1zIqnSaGfJNDN+o2gvDBT/
yY/WYezj8xpyRJSlkd/Vs5J73/w9L0xKsMv21B5sC6VhhNGjSsi4WP6vf+XE27DyAcoNFuZ2ZQDh
mGpawuYOBu+BEshkXz3wz5Rvd+fPKLjznSjbjrjFQHD5Rb+XBn7FcUFgktlQyS2LOMvEn+lbY4mU
gLzMCxDp69F6wJL22BYXI41S0PrSJH7VPg0Kuzwt4nDCugm/XULl0Mt+3CFkKkGxqN6WJvret/Sl
z/iMsyfY3GlwJqcV0X7BGoEhRCJDqg/eNX3IxdRvPr7/xwx1TbGxXxjq01YPzqvl5BHsEUaoCgU7
30N2aehUgnE9H4gOqKbdHstNlhnNgpNRziHDJzjk32fYFPdqT3nuUUDm6EUe+vN6qC2sAo1NpLeX
ofb65auxk+bVTvrfYEZRrTQqVqMuql5zeHkz2dkY4pk9SCQmNecWwMD7GPfOReMq/AFOzkSMDMcQ
s8YyATpV2YmN46QU2prX49dfV0Tm9YHw5284GwUXTh2h7yHN0+8MP06kYAbg5wPOiM61Jkfdbxbb
fT8xGgBE5y0Jkg+Z2GFVabpz2VBmALjRd7IVWxClCzaOB/VDtH/e6nPSPyvV7w5iImgMIcCUXId3
cLgWlm6/2/bNOppNE8ju+gwHOxC7iOVVJQm3Vzo4/5RvuxSHSf7NBfubY7hd9uMzL1C40Ee9+Y2D
//J/FelBf9fBI5FNIYxAgF7+QGRIF2i6YEh8hGSeTG/bAasKViXfmdw+ID24msHVpnUnahgdIKUF
XIdbNf/gtp18rX4nyMMtEcFkkqBpONJnpdNSk1y7WgmA0ww9Gploo9QE09yUGeWr3cWQIh7ttxjF
oYVoWGtBmJHBQw2K3f/R1s3EmoDh8dyOPz+lm3Fka2hEoI3O833nS1HoiIrnZ1g5j82+eYc+Qwuq
P3uqTgWRi//mmXItau48jhQRwO9C/1T/5g1huu+ltY21Q7YG0QHOIU++uZSb3GIaHUgsntEs605h
G9+uWTlrn98G8hpvB5d/eCoUeYOtWLrg1KEOwBSNyPLw3vZxb2nRn3MI2YsRusiQh1gIfiejt4YD
kfpJH3Zv4QaNcBD7Kln6DHWLUS4icKOhh6R8I0AydOtgUIP53QJsKYTWazgzOFHYJGKtbmzWfNbj
C7uO0+8LR4H+ct8seG4McZaTIS/Nsh8DVx+7Hd+Pg5DtRgve9Mx0j/TOMw4YvEKhz+KkULWj33ps
MIcHcutjU36M+ru1llFCq2WBgmBaXBupyfZ1ksgWIbwCwRZoPUcNM3Bar4XyuG6TDQA0rlWojHEg
dAnCgV+6Ukyahk3ow1m3W70eeAqshlvTaBpj5invgSXjGualItkuXJER55inwvD0SqKxUQhchtyY
Fk5cAz5ljrnfXWVyIJ3jgr8qTXerN4dwrAnvSM2F08VKh15i6TNepWxBhWGmYNIb87awNGL7E6mg
JlysO58ZJWE6NuskgWUi1HpqNZQXeEoAILIkZg1vYe9kOKS39hN1CYitVqcPrMrYsBzr678wZwdO
N1z9Kj6M5ENnCsp9DYKDeTHV2HLbNpKqREPuUyAHa2vZ6Dq1fq+sJ52Vjz6OiCO9tAEsHapSwA5X
qXZPdtFLN4VvopOeG94EEGBHkZ47KHNNk/DEaOr/K9OTBTCI3QBgImhCpRadGR6X3O4PTYubF/x4
3H1ZUUvEY9WNQrUWqUDZDPnammQxHvWYpwgQAYjfVEiUPMm2SnyMSoAhsrV34rEGJMrcCDqf2+R6
B9fFyvr0CHtvJj1xk+EjY5GgUamIiLGYYNP4LbJbulOEvbjjqlYyn5bnFxzPWnNRAfHqVW5bMgde
Xd4CzQI+pZn1nHygyveVx67Gi0DeWM9pp9Uo0exmWwQqVey3oYimA5MmLfte2C7PT2CZXf1cWJqF
2FrGcD4JT6wLBq9rStgpv42ujWKrE2zjeketBlZ9hzdgas0CBQUHTv17NFTepRK4D5lqNU5O8zdd
4sUw4T6kvhP6p9PI8+UJ+qRrZjX7l+xv7TP51CUYpYdj0Vk2FMa5fpJuDnfXTeTiR9YTELAG1WmI
ssZZluaHCXYxEoFqTBTBg7BP/4tAa6AmoJrr9SWTKRY7uFcH9O8tQYD73KzqJlpUyznF70pJsntU
/J23dkf+Kpa23bR8PhcHIb0fOGSq6SPoD/CwJMpnMCvBPOcYwHRuSA7hzxYAD366wiOgrfvSuWV5
DWA4nqXTaq60pO+EssbHUicxS6zkNGKSM1jZClhPDJOJvZfUO9/lIlbzC5QjNzz1x9+mGzDO/f2r
KTcHhnafJCM5WlXACO7EtaESoyoW2dOIOs1sRA8j0PgFEDhmqgWPTOOm8QcRnPTAi9gc0sfd+mJ5
GqjHg1K1I6SV8H8c6qjORMlfhA7Pb/WlS2ZoaS2U0OBrSI8n+0WzITkWfTVoWnV3QxQbspkvG2SW
FhfNsinX3yMUfExhJa+0KEknnk7+64If1ZAFVCwNiBUxxvrps3/OVI35KaSgH7LegOSsMFrd/qyb
0sFfiCriKL65RBkns1QD5WWBOzuBRRSAvPejbolZtDPNFCjnI2GDRnpJ46Yuemm4LI+TfQby0HPQ
pEGksytIGGLRGPkKlaStAxnCzOUlp3B26iga5bmU9Hc1YXSn2MGCyLE4fiAj/QxgxhNhwuZxXcjs
lFiHJ5+zBigIA/sls15a0g6ZAWlMN1AxxoZzwO4Fvd40LJAKgede51kyxr+QYnUfsaJ0F0LHcIOM
wpTYwtojXRkDnI79xLOdLyeRjDDYDi6yf3QKjh1Y6RaW1Ouhj+27DlpJ/KouCiUb8Q+DjXK8apvn
ImjHidNdb6WiLAR5sFDI0MSuiRBQWaewpscxB0rllNaPDZVc9l+U3JX8m738Icaue6wnlb6PSD1q
0z5ch7j2e5P53DmItKXVp8Dw1h58JD1oOhASvDsPSwiz8pdXXi9z+3weFj4QMJ6yWs+qX/7ZMfMV
TX2KtcwPgUGLs1xEOPboylwiU3EI6d8hIL1DjnR9DQSXKlUpuuHl0PtsJ0/qylKRnqZJAnLtowJ2
Ru3N7BVXn1og9xTAxpMcYH6tj0X1hNKFsswGSO1MpU/3Jtan4/paw9tqmOkM/l5/0aiH3eoRZowm
dqpJfLNf9hiBV5OZwBo92fLyoFOIWB5vn4JOnzOXSb0lMktrRSl1Dovae70POR0kKZhvZptbAGTW
YpdxKN75tNeoZl5/Z2KLbU9zZqXcCjaB5/84pj830JENtQPUSbKVmq2UvKGNcH8yq4INhHIahtND
GiMxoCp7XanZsN559CmlYBgXQNn025/ORmflQKMdR47R6t1RaNlY4LUHz3GYTUcNMdPTdeu+7MQW
tpsjNT6BUqbIlf92JCbMLesXbtS9HcSyEd4ZmOaqAdM6NjDVlx2suDgsjPE7tzuRZCYoBHDcJNOM
swVIKd8KeuMoNQPLPVjZPtXAs5QM0HTZFF/2QjtzWCAT1Psi3/ID/78g8R/TBKlVHn1KTb1dBSPT
edkK1j3QgcYCmzIGTZghMy/iI2CTb8iJukU2kWqPF4BKNEay2hAdpSMib5cB+i+AP64nQ39HJY0K
6WFoyNeGupw7dcqJYOFr9SDXxX7FprmZsIOlQRFWqW5rYW6w/ZCBDAEFZAcpW9bXHXO4801mRnSB
fheUrJU9k+FRR2kx8MzfYXY+yNhH1TCkjqHU//r0dn2SI1BfrEwBZ/mWe+0R1/afbih0+JkZCw2q
nVTunkVtbv+pTsLFl7UkFRJqIVDuuRKd1vI45sRtkSW2Uglym5EnqS6QyWUxWagAjdRnqkZUItp3
34qMEaOqtY0j1LzJxEZfdevmJ1Rgwj1zES92DzknugAX8dTCYAy45riovQoIGKwJYDCWlC0j5dnI
//o8fEs8ibNtQlq2jH6rpaw8TnXTdnwFJ7C1XrnIl1YctDCELdnOOou1h8k10ckpOgrcFsvipC2N
YX+wNZ5dJyaCtvWJmyb2PeBIl2Rhez6mvpiNFE6I0Yca/gusYM0DDFWfiBz/I8R5a+ztEQlqNZAk
CJe0jcqAjK1TF0yR7JZm7C8wGtugem8rInsjg5QK54LKvAXXLf2+gsLmc85KmrKl4bqNxtlnwLC5
/pFQTQEdJZDeUqB2SKQRjwAuwa3X5SJqnn+7aOomBOuyZgoNHN9Icm/2BgLag6/pf0CzTt7qbgku
TNQ9GSG5zL59AregOPGxK2tWczdRQQTf2emOymBnBHa0NdHVqNfp6BkWS4D6rFH/0AsKwEfzCmu8
08g3dXa4XV/m0hYRvwMr35i777ztaJzvtNr48zC7VmhGj3j3noIVQXBKKxQKfNQHfObnUthoAUlz
agd13HFKlpF8PZiFjPbVos65L6fAUXn0yXvbApR02LtPZkVdxfwzOycWuOdHnaV1/Uray0zxCs03
zIvlHse2trIhZ1ue6ZPEUqpRfTLbnAm8Q33x4vzIhPB5m1CF/hmO+RQb78Hg0WW07QdFQp9eYvuk
DDZYJwkZzed2xixEA+sTRlb4ueb1jtKaoBZA+q/p9BODh/VgqHBD6hMJcyG/kMTJHbQH7XiLquae
sXrskwJJkjboBgvhXxJAfbGIXWWERBT/cPDEAZni+55YTe/oz/geyW6vBSBkYCLydpQ4YQpsw45O
Xa13zMNOXlZtpgxGAMnmHzXtgStWkrdccQxrQV5UhN0QQduh41LgbgQS0IEX/SestF8NnBwIZpq8
1efavksx+M0kwIYFX8yBh6XBcGSSLTcL50DYUrHZh4KWo9diCHWZTpzxyRTdADsKEE7irYjO6RZd
KxR1+Zs+4xum3QM5YNIZDf23+HduA4j42SX7NyB7ZQ1iWZ5XHbsBYBMuvXLwtDi2c/rhnHclXapt
yhs/zpjrNUcfnCep15J3ZqmwRQ2hoKxPbjAgTZDkDHBFGRioJ42mVGq1ugXKWXNw7suHuFohrUnU
zYtK1GaJvUFXTmWNB1NhMtc3e4dWJ71wGdHZFdKUyVHdeX+sgVTxy+ECoYIwzckFFAbs66R2ofx0
FdZAARO7OF0ClAqQfaqclAZfDApJ2lk2LSJofV1oXi7OlmBe0Ll4CuJmDYxW/lOMGjcaFOM2L67y
HvkHld3/YahptFMd7Oexjq/BvndIAkvA3u3Iu31lok27myRE8/I4iBghcmTYnQWXRv87+p9GwZd9
utd9Zh/PRAL+0yfNIF171V3cu9EwXH/K/mshfDpqGkjqK9glCRmwdSDVKLT20DeelSTsVL57tmqT
Zp5S8M0BwxSQD0OuWtT7+YBfDuL7qn41ZF/W0/7tL2pjVR7A7GaSqoZ6eAtnGLA/pc15KIVRqo+r
9blNhWSQZt8alKXsGQenuZZdFAEmscoWHsaTdZMvaTiTByOhMSJMH1qO/VukO7qC+bq0ctS92m27
dqDozsu2J3IG1wlQk6ufzLU8a6X/36euhdX1HvDagggW8us4m+acDhf5ZvQtTtex7XR47xvYYhBK
QKs7CfjaSOBhp7QcdvHeXEcPvwBRAJIR68uvugNdGOu+kirbKpRXbYgsaIbXmeG2O+qeDCPbJFMK
eQKRVvOxKB3o/4HcVTIavFgF5TfOx2ysA8MT9Vz+9Ybir4Yaz0kKisCL2UfrDzPmelS5aRY7v3Pn
uEJhzcl5NW9jzbJTaUf8+KD1HPwCqM9LNHOFgVn8KoeyT1QrL7taN3zhS7VxHmPyK8YlQZxKYpNt
3vLvhSrxTHtj+1gAcLI9lA8IrGRVfoGoYDz8rJEsndIFK8vhTXOqyVGekIwjKxtNSZcF/qIHY91h
ei0Rnuw74VCUE7vz46uVKN24Tt47J2TgmwzQJolTfMzHbl0GO8P0mcZVMgGuHt2NUPjQ8cKpeYb3
mzVSWjnHGydN24LYYthQA5GyIc3s7ezrBqE4HYEBtQzrTbJbLA3q08aeuvVsZVLVzresnJm+iC0P
Yk6zdK0DSy00ctZpNoUHyqm8SDV5LBvbO34Ar3rgDLtO9M4PV5j9idSGpmFtkq2hBhU6773O49Pw
2EoQjRo0EhQHE6ixf6MOnDeX5wie2QO2b08YlKVuuOLfY5t2nxOO02T2AeU8G1e0T8dl4Eb/UCPq
7aQUgrlNNE8yabmlZ8lrsV9TnKpNCN0/TwqP9GsHU8Lc1bnwYIsYFs4dcARn+kfXotJ06TYZiksW
m5JB/pwwENcq3gUCdbE4UG3VXsTCXn/RAeqiy4N4uZaW1ecYItKt91BrgPxxEkk4e8RbBlJCe9VG
rvHg2B4XNyl20n9dsADKPwmnGA/9BLUo03ZoMreVdhRsQVkYzJVbJ/X4BXfKDL8oIf7wSabSGweM
Huc0T+qjKgyjtQNUvw/NW6/EqGZAUkAMNsyKHFnQsk2PasIF8Mp00l884W+VtnHBhUva8pUeCTxx
wBVgKMZZZswINKZVPzQg8pvbiYkOdDcFNpwhmArE/c4+JvSi/xrnazz8cEOK2xmVf2K2WD9MAR1E
bw0X2A/Ypx7ilWm90r8QMvZobczn+6uYIYfj85VMAJzMWuIIOChZyFjo2WdmAr4DS5K53f5AuP7r
As3E5i9iz2N3JsSFe13S/vov6HdZZlG74jpep5mR+iXOr8jL2+5pmJb/jONjQlhxR8/55hkPmZPC
P6kq/q4OGxDwuyBG1BvpyFW9U/ypDOS7SoD5GrEl/Fm2TU40dAU98DzdmVzZYLKq+Lnya4kgQ76q
3WfD33wCQqIrAIo5+DFqkVSUW5r9dB9yCvmcTafM53iGocbd04oRcFx3QeihnHm7tpYirDTpxaxI
phjRVxUlfsOaLT1s2dlyXPgz00yenOtCEUyImYKb3+7jXx47Z5PRee1rI22wNvxEt96f1CQmH1cG
HaERUTvRWSOk7ZaZZdvy0fyEb0CBapTgpXmweaU+BHyolTAUPIOY6mHoGrNys8RH7B1CGQTNkQV0
cqGcKcsJAQk3UNNwkTmHO7r2qq19Rb1xgevzuYMK77zHMwAjE9uH/3T78phiBq38yraUj2QF3iS+
4JtrZAKNenv3+kmszSIVQ7j3Nwg1u4RJxS5Oa1zgnAA3B0iSiToYqczVQ5e1m8qxuM/h4h0LZOC6
Iak3hPnUO3P3PqvK2ZtEpJWuo1c+3GXQEv/E6WXgKSy5PTjCsm4A5O66RWyHvR279ipAmBZbUUP4
aYfwih0ifM8vorrfQfBtZxGJFay2auU3Kn30LFyF90YfEsSyWDLhqq0eGGKS90HAOVX822zFTDO0
KaBTxiy1Bj0O5R9zy1QJ4Ix9boMBwsOemSYAfHnIuBzjHOrx5yAaKiCLwzFeYdLabPeJRBGEELkb
sMTbBPv76N7ATAwYryZtAvMvf3ahn/Xi15fynuBZxFedR58HiQhApZuDT5ljSsAqSTgj53OUcp8G
vCrJAMWXuVT6ixSsZYfDJa6at5WOsZxutO3Jb4/llI3dgATcHmNswRb1oSZPn2ji5dMDEVg3CCLo
8JCZXiXoWnC0AAz3GWkCGwvlBPdzNMjVoR5nspPAlmRES7l7u8jo00rW+w3ih/CU08z4NO86xymf
mpH5GCB/zrMnUdYp+7PQ7wVXXj3qzb61Uwlek1bEQ+bJL5DCDbSOg/z4AI8VYXrdsRpV6bbnF1MV
H8ioh+UQfw1/ud17md3DhF/jUZtbXCli97sN3XWLGw4TCMVlrmq1VbOx7T0CQcdAJ8FwgM2EHXqk
/TGArl949fyrqBJyuTZJF2FLrpJDtQOJ01z6FgzNi39y8rgRwCe/TZClMB0uA5mbB8XGvK6QQu40
o4Z7Nu0CIWFzTbGq5J9iaquBZKJ2VObZeif8WQc+4b6p+8FzFdiVduPMb5OsMTPDyyIjv+e6jxXz
AzQEwnGBaPG4u0hgfgQvusJ6pNXMyJlcVFfApwsqluHabr15cx68JK+0GHLGCsJ68imLQR85eXrC
PUvgsWlqh0yn4hHqsfkXcYzNtq+eSCAzILsTEujphkF8gSLpWOumQpHmBa3D6sXSU96OFWT/Flkf
gXyQVpvUsrDp2d3VAkD2+wvy8kVRfrlrap8TVHGWgzSDmpQVNrFIm7TKhjs578g0rBD+00Khjq69
tk8+L1vbjyZWlqBypA9E1wBYjoTZ31Zxy+rpIVqmF05Io8A8uaXb2bPhyKReZDZok5BekVAspLvV
RbRg8kjlVJvKokVU7lVwLMwB+yNKRxsqpMNo8PzetXqBrOxPaV96eWyZTOpy+z5lvTiz2dgY1JaU
4taNxW510tKg8/wlSpxWGfocY9NHUHZ6mw1VmpaNPO7bloLDiHQiz0E2xIHvMVZqgdS9Sp8g29Xo
DKz7QpVBvXMEG8NQnKhzY37/AI43Ccqo2F3GpkuLqQ6V280AQ2m1Sx1+wHh+gksnEwEqej2NEsui
8c6av3Zfpf5j9QsGkpICB6gN0mExseZyPeJkRnoS55ogOXz0TMOND32ygEqPnQJ4+9tbEYsBF4kV
rTjAeRdVWRw5fGXG/Ruvt6JJbEevmn5YLYCybALP93e3f4/2Hp+Duw4H7Ppwi+OtSGzSUEBGjL4L
RObcvLEIX0wdCbVWrpD5AoWqtXORk40MbRPH2msTPnmFueM7x0nVzjQuoF+kn0A3VDWGErGrg+wn
fjBq1dWnUCNvbYo8mMPnAoAco4D/1/aGxgmVdQNx5DSJRhR4xVLqqJ/mk+YJzAp4i9xg/e6UFJEs
v3GvAejo8QhUoQ7MNlXBlbgDn03GqXA0NzfT3XwfAyW8Z6JqBToMrEq/zpCxJGz9oSrJKcL38ZIJ
UU5PFAW+cbtrXI0GUE5KB/SmflsJ1qzuk9pFWZ0qxFZBgcipgqdODo6s2H+sUhMKOhMDjGB/4IAW
HzvbKZUF65b3VdJwe6w9PVcEJ87Y96JRmBHjS9UvIwxASVnHH+lc1MBs1d5lqKgXaJyjVCsIMQhy
CRMWH7Mq88lmcCAruo6w6Hgne/ApvezQaBwmLBJKc2+IgE4dWnwusR1d3OU4+3iRCteEvwpgl/NG
ML7DZXYBHTlKAx25yA3uu50mNVMo7P4qxzh5631ZLYwb8efreRzD3Rev2fPJlMrPiZAf2HcIDGwD
i+ftvDaIirle17HorXFVw6sGK/xOCJW4XZIR7b34MlBYvPg7mZphis7osAT7nUytfifQQxB5YD9j
VtyT6RHQwFmxVSm6jDAWHttZwkZn+Q0Z3kWU60u4MKpiqmNr6dKJHOpAcpgg7lHJBL44Fh9O1aRI
6CZqtk610ldwxc+qyqVlP+bmPPsoKzP8gTG+UZ0XS8oOogqOcqOYI1lyD6NaxP1PT6jDrUVJJaml
b4k6Lz6VsEpNT5mEBI8XoI96L5PgfLAiWg7TBeZkITe0XDeowt1GjrntDidyna2NG3Vd6yuMxPGq
Z7TP8KCP3sp14LQVMIiv2DSmhh0CNMdrIQxpSR7YmHiW8AMKVWF0OCSJcOfGNn87iJaU4F1QBHlP
n5NlxWQGwnDopIRHcAVD+QjCkKeo8HGSYl3d4E154z2Bk1PZw3wR6F9xCP2OMVF+Q8gJ4P4mOR80
Ph8oGJxQ3IL9FomWDkW4SMdUYZb6No5DVJtymzFmpMnMNedyb/f95nz9buB5CrouIi6sNpSjpOdf
XxAvejvJiiif4W6Ge7oCb56vPUHUxWZ21R7SOhkF5Ns1nwWkHDUORE/YyV6RQG7mgdseJnSy+Kef
TFF+2bO4Bo8JLkwyM998AQ0Goys7bOzmkuvWo9u7KMupvChSyV72yNFA5RUwd/M/o2GNfXQBcM0N
CymHs2+h0HnINC4sut3pABNnYQqIgfRDPRiX1TOUIV37DHs7LZMJrVHeUnvPwPyTWRlVnI2nimib
smJYdIate9NN98Rm5WVRHzUaZUP/kXhH4Tdn7Zp7LD21TRgECak9UDrggled+CdEUC19adc2sBnA
3N2UX9/yQG7P3H7gONJlyVKGW9nZfKV5HYGfmZ+O78b02U/4yz9Fkiw17PLMu7VPVm4iVZEF8cJ6
GbYL4JYeeoAfZMUpRHRySslF+FhdjLn1rwUnboSEZfJYv8OqAyMQ9uUg46EM/ts0RzB2B6WQg4b5
4+R/7C4FHMJ0A1YzQDx4g7CzsoLSUZorFpwrfM1LgyGv9koLPRhLPRJo6ya0al10mam6b0C/lbDV
HcIW75UXHXPE3zLkrkozT4erPawPSdNaB9g9krdoYuIZS9aHI2P+TI6Uy5FlYx/f3t7149d0+Xzm
xcOAoJb7vyKGSblyZGMfWT5oaXEtH0iJ+ewHi5fCRlkMYvTujSiLXLwTCjCivEub6CFADeK1RVr4
zLzFrpozj+YGda2QrOpczJ0v1VGiv+saXF64W4/roJyK/FQFdrl0vYvjgOj3/iQUT7L9AFaO2tX3
T6gEiSyoFLL9b0laBGov0ubvwx8Sqf9dRukfHmSstvCpkXxwD6uyS+r3NCm+x7xIEzIklc/NrcWo
B2x0l2Hf3C1VOrFpuJz/+WPfdoybKGsewjplJZ49rJDd3KcXPS2bay05QKPij1FZBnIQEPFdLK8H
dKztiL9cVBpI4ZAEQoIXjjFQh/uOZ4lMEqDC1ck5FQVMn8oBu6i5bso6AZ4XWUNTMkdKp4u8E8nY
daYEZ2PG++lVjOd0xb+73lzc/SnZk2UORLOI4RcH3Smu3cTHAc2D0MPV4dKLPHt9kZgfMZNRdWym
GPQAfEEFh4qPe9p+j4BPuqYB1vn2EpJcRVh78MJwZI0RvN2/81fEYpRN+nNjQPT7oe7IXn46dB6y
BGyNsNEsGT7Fq0T0Ac+NANedkRR55NJ/aUHb1sD9ld5mMf4GDf7Iktm0ILFlsT2XdTy5pggC1DR+
Xa2Mx/FwjStGsopQse9pxYi6e96RdPD7ssVOfhvq5TmQ+XYMfHoW1gDYaNdZVzDja9FGYeKGTBkS
djuXtCX+VJcftJiN79BJ2RX/j+O7GCwik1txYUJcQKJwu2kDN6xm1eEta/8vPWoC0DdYzQpOuvjM
M5exOAHhydNjOj46vxP5a1/cLFn8tj6/nVn8FsoEdn5SKJupfAxCaeF7f+kLuY7EO0AzsJbd4dyl
FZeP/XPg+uEm3fcsJPA7GlBhClepd4CypKNdBZ5Zf9eI519wCGlq7uqZcy9AoW+OpcjXK6VNAqBo
mMTaLITr8sQZelWQogEMu2GmSFiXHifJnz3NUWC3zuRK39dFGvdNOa+AcrhA+Sa8fsU/3pkC3BvG
0xdxU0nUySWmTVw4YfpuE8rpNVo+/F7wOm5cUabifob8J/fVrxokho/g9WCm8V+7ZjqYfSBuAGiM
YJSgIQndTf5c2sm5iYT978PZeQJrEVLb46l683s5pUY6VMvLjILsKcPxuEY9BXZ1xcdYTtezutSg
WqeUFqs5O+FzKS6VspzlIxqvi9JD8vjtG5FUvCaK29p2yPtQ3Nc9cgYIBpoSYLcx8zFqHtoY97Ms
gYkXOHGU6cXQbeRx/pScjycIxWXTPsw2tnRj0EV3OubRdvMOVX+eqA1YHTZv5P2wuj/T0kysy/EC
xsHCplv1JLvnDOaMwtRBMuBYklsYEGYk+tIiSqIa6grfGuNR2fyynBS2dWRT2Rf0nV7bb/UkDHzm
VZE5WqEpIl93NM06xTE0p6CAkzX5mgW723I5GNrDgA23dCyH2zLj02TSYKPEX/KS0UiDD1CzdZ/4
jg2uLENDDVpTK8jVVvKukEl0TM7kXkxntTcDAfQUw1TTuJPNNTzRQELXGerfaxCRTm6uecEYHX06
rw7ECKktu4oQbX/DnGl+K2ZCBQINrPAnpI8RWzc0a+f9ZKwvywrIyXNtWD5f4TK25vk2yNgGh/Dt
8OZ51YgxMtuF9haCZq8yFHqsrBAZPZ+2aDH5T0nHyNw3UzRS+PqwmtGEVvGD4B0a1KmCvZMs1wit
pFm/dOWIBiOHk/ujU4M7HYYpU53wIyZA46TpaiM8CAkt4mqEzMVMgmAFJmpPovM0KflnZtdBS+uJ
hRzuvc2+mpILO2lIx/gkABnkD9c2i71BnHxHrf9QI6B0zvRh1IHoJYXMkUbMMZNeZtCFSVk0WF1P
irka1efxjBf9OZiBx86eR9w0LKcu+KTnJ+iuxQV31H/cTi2Ew6A3b+BS3yGFYMqvlj++Iw50DX3X
OrARdsctPwVcXVDEspXiuuCRfxZJOEYdgo5Xfyc79B4BLeDggVpAaOafUkgUzg9SYcbBhS1roTrc
UprKfg6gxr/S02q2oCniq6WPTvUgwjZYuKljeqj6/Mb2nraU6MH2tjojF7Ztgl2Z3bzyayPei1ea
D3H3/mc+sddEnSizrW4/FK6PD2CZ33pIrkPZwH4r9H2gtuLFd8SOkuzYFKFLd5NtF+/JhMYMFVqU
gRX7BpLumepH0tpWeVhEQfLOIpqcUHQuKmI0uVZDoczjjvAnWzhe7fC2ncLBo+c+JR1ZuiNb1RtV
bsYROrSl2w1sMscc3oWhWELgloaGQE4IzpQJfhfTZRkDlfZjGK5Z5ZNZN6A3QHeRE4cxdKaIFPnu
9roOKVe81Sjd8Bi6jx6eLIto3JXFjHsmpFZ8ues4uwlCijTaEV3HbuFl1v+Scf7GI3WSTkhlU6rU
FPeD3KZmM5Hnrb5QWdHxTtssCSQboDDxEhcbVB/JQ2XTMAQKQkYAnalxLTTWvUGgYynwmXTSDzkT
ka1FvCCX44rLW0zzW98Ej843LPCZzXrXb5YTjhVWbU9GmbBWsX80B0ci3cBk7D/gItG4yLWiMD/f
wo6YVbhXoplhNMqMP/P5Ik6z2cZI+yp1EyUDCjk+VBMxR5qjaWZaphhXtcBlLqjaVSy5yjrGPbwN
cqD1a8uhHFTyYesSuG/U84eqdt4QIkzm11n+p5Zi8P1s+wxx1nrQpqdT4AGWbUpOM45AVuf5L/lR
I/8sQFQNZiF2XTHctX7IQ0rkB8TNsFSWk8dIWHY4Hp50XUmiwpb98r5uJFL+QfRvh1UwaG/wSc6h
KsNIow94k6vgUUHxC6tjIYYPfWSTYSZMU2oEIZtQR/xP2PC/GfE5+cu11E1VPJU77Bc8GnCT0yCA
qLvqf14r1yV3zE0rZ5E84DzXJekZRaCDHr7RDIfkvZGJFugYLjOirP99njv6/iI2bMy035QN59r1
wwK2D3EayC9kjSyGyP3WyTF5rrndEardCy3OpIOT7JsoAqkfEkOYhw2p/mpJ9ItSiHm5zJHqYiVf
i3sVFswDAAhwqctyGoavIoLzAhgzt1uj7XO582TvpqDx1g6MprpB+wxXN29oAJsD0w9KKjnOm9rc
lgb5i+xXBitj/qAjtAupLW3P8fQTIw544/e0Pl6B0R4gOcfm3jH7tYFbGMcsyX+kHp2+xguoFmCU
p49+dOSZN7E6eS5iP7Bsk7pyBVoHfzfSVUAqylWdutSNyRUiPKJMDW35uvZ1IDee1A9YRopkIY8p
LaikOWED3cwCok1qT2YjVXicrw840t8RWSlUreTaDfSqmHudaf1x54rEiLYRuapA8K6jehMzD0Cb
kEpnpj+9AdORh7/9qVelWalkOaElHIRTOEZHSUZlgGho5xaJS5+wXrq6c0UrJLEMhUJ6/+NYXd9G
2yGjdveZvuh/Ak2knnHnrjAdfKiVgz4t1ChBwUQYD8gcj9MIMffc8eb20+vhQQWhqOUwsBLSB7cA
4S4ON+4iBV9nTL3QtDl8pFzPfxohti9NcXeZs7XMxltPfr0Ad9NyCm6oFD+Xc6bLo3AY75sPk8/t
RdgiZl4yqe8Fl8hQrmMTxXIarl8h/bHcsAnaCEoJwVPwIF0+Vys9osNu/4KErrVYq2ZIaUwu2jNh
4eEEo9GaA6XCq7MKWUEWFyPtM6BfFf8keqpVsRPLIN5buCImT140E6Dp1MH58rw2LQ56nnbZH1uX
kiZQtxqKVdMfcsSJw8bQtpP1SSQ9rsGdx4swhgUSLzhmEsTX1ad4lanXhWLHLDVCPiCg84D+xxks
L5yzgB+g6nw0i6uFoBovLJqBjccDHFS3QiHdTWJHO7xHlxo7VMpabpZBemvlEGKg5nvW3vB/SLSn
e65HwBFtpEpBUurPi4jGzUpsb5ZMXvmLaDvi8qAIa147J7iYtcQeK3tbqCp86CviiedTdFpCYbAQ
tTHyFVbLNzaRaDoosCfZ50axV/PbXJ4lXZxJQOdIaK2QBcfl5Jhqd11fVKLLM9i8EN52JgD0JDMh
rQALhcF76v1dgu1IZnWqIG0o4tSOaZpD8fwHBSHEE7d5YnAPelobhFrPkf547hmPnPgbZ5oMO4PL
U8m4a2Kqdn+Wmy+oQN82Es2OQsUF5Pi3QC4gCpsYZUa1QwPfQP3lfZJYUqC5tUplTTMX3ayPv7Ny
EomR6Y/jK8L/jiIysVIlyds+z4oUBKLukzTI7GOtYc18yDvEUcHa9ISTJBqZXrld9z/TJ/VCvJqx
nLQD5i53yHZ7WqRxVLQus+TL30gwjN3ytmKzWIJSDcu5yPKFExRnDOIiHrLVLeOkOsuqId4ugXwQ
3aHtk7OiuXYez6k7o2VxPfOEviz9NMLUtcU33c05tvqgdHcU4EcUKANwlUcH6Mph6PoCio1fmFcj
Lnrekl0COItX2qKCvueGOR3qfq8opL9xq5Fh/4MFLb2uKbcs9uOZrcWxQImDw5z5hIU9XnUZe80p
5qU8HEesF7wQajjKX/bOGbVs8bOYEhj0lnff3NGtW52wO99OxKKKOeeu4/FeuPUFhpxxP1IqVg8+
oeW8YaS+RZFu51PkZUbCPxtDTY4RVmYFOFskluV9Tw+gF+igDcfqlsrfX+5CMn6FLdGfehmaz/Ur
OiLnCEQV5NMmZj9rG+GZIELg5zyqoj2oFUNMCNGj4c5uCLAgoGK7GQv2EhNM10Ma0hIzCz3Lindk
UvD3hrbVAe4sZ+QA9Rv5KxMohKr1m855pKCRpjt6CeItblw7FpXa6bFCl1Ka4LGJKc01fjLlcCJV
cViZFW+apgEej8YdQQiH/d2CzkAqpIGJix0w534IWk9Gq0nxtkCaMz8/QAT6IOcFb44gKb7cRasL
cpAkwXaekMyUMAceUlMVifG19R1QonGCpiiCN6LGVI8wsEBwXAf2Leegzj6mvS1ykaC/dPtk9s8g
K5MPyG9e+hTEiHke4vRGPqRIZXMB0+PtQhYaeFgJXXc5w2edU/gTYufQsMxLAkuxxtnft+/3y5s0
2z06aToYBApyVlVs8UycUtY1ImXyLxBsloUjB6ia3avgvt0IPJ+3IGD2chUJ5IWiOuUqoWs6uZ/Z
vYn90i4bpkZqmHlvsr5F0Uukh6dnwQTQ8TQCJSrRJOEX2JuldfKNrYiS4hAng0Pb2kC3zqyaWpUc
uQRNui388P10dTRrJkXQrrhKV6iY3zogU2bXQtnl48BXhH2CKy86ea4BTij2ylJwdQRviIQLQ7I1
AWiBBSMk0ycst72bVDdQbtngalff78cmkuR4BYTGoR68ILLD6tl7S1C5+ETt9L2W7/0knPHGL74Z
NlJNS81PkQ0bAaX09mVQzI7BlesupQWTA/D2EIg1huVCVDb02eqimH25ptJehcxxTzUoqt6cuAb/
J+xDznq1DGB40aJnTAa5KWqK2ukKbtzFdVTKxAsky6yYGTYIjdhyzvYnAPDAm/xGJQRbBWZz+69H
1k/c5Aza19VXUw6wJleCaqHZ3hhYFYgM7XKkYDDgb4OSh2sKlvDC5nuaY1wfUR54krDi+P2tpvCz
3WE5PYnBhc6eWQEJgo8jt99v2ZYuTpYHqCRCImtEjA9y86yVJ7MYA9GmVLoZ8P1VZw5BMi+nlQFv
OAc7hiWu9zfxZdzcYc/GgaAwftdEMOMZ8IzkwFJx6zhRW92wrt87zZuRljycL3bJXRXsZxmQwjjZ
xWEA0YYbvdRr8S6J8M5upyFuG/kqB1EQXHHgLCkqFaGQRUyqwLfBuWydyleOD/jvSyE6whTgCurv
8ZrS0GcwF//YKuXzgOVEUQ3JNAzOlaBaGrAU4EGNrmMTZzpyMZinXFg/8uiOVKp0IfECgVpfteo2
MQD9ejRut9SsAsPsuEy5UstekEtrO9vXDRIlKXh38LP4WABof/0GlaaujorzYvJRfqcY83ciP78d
euQRUSIAJ/w7ewtq+i1nunyDCm2+CC6er8Oi5/e27MEbJuVL4BtSU6l34LJLYQhzjiKO0AnMRh59
FcbfYzBx7cbdxMlWheJRPFNIfu4uwaK3rWTOOcGjJe0EBK4AFoWLyRAN/P3/uRZ6Dr/n0S+DPDtX
LRp7VlUTRnbxSzi7vv0wledsVGSYqkQ1BfYprLN+vqLkjpUCDwd1BnnAVxQjE15+ZDJ5vbCuoHS+
DbXNF+YRFhWBm43ewcGZgmxM0NrBba7jQ7lTdTzVOejYqJ+Piz3/vrm8pIKsmHWuiGAluwn4abPy
Y7jtstodjRSiZw3EdU8UZs5wXt46uN2Pz+hkko3xr0xojTGaO7n7E19QEZ84rA91nw1dgbYsTVXf
flKG9YVqhTxDwsyAmnQKVW8UnY5P+WGjyIQP2itBiOYoWZzwGx6Fuh0czTm5zbEenEsPJvFlNBSu
eqgRMykYHH5+52ksw5Z3rFUIhtnoG4xdNesbe4f27ryIhv4+TlQVbKTDyGh2R7GzboGPh5guO1xN
ktfPly3B+4f9L6NGQHOn5qbncnCZUeuPe7vM9cG8tGFJ9dMoAj7Opr4h3e0UOEVxQxX+rPQBs/Ng
Hb96p2ENYxvPtUcw/bXx7Uz+buhWo7Lk0jFQ8tN4W9il03xea0A0wod45o8vgQ7WLiN7d7M1Jx+t
JY/HmAKWpuIJiAKQgdCAwCY0htdPG6+n3cNtIjyNjmM/dma/eXjBVCG3SWTzS3QWr3okZ3Z/X7L4
1Ga+Z5IAm2T8FKlWFhXtkcXuw6vzzEFXMR+oNUZgaD30apoT4RDs3lK4No1m0nnl6E9MzYuiT3BP
5jazucXmLIMN+vcT418gIPqz9Aquh7SYYtWiTK8373VQ9NB0SXGLIZ8sBXESGk6kgW6+PnNHSIf4
EvtVecNcFDbVoLsrYhQilVPrANHXY+WW0NCLbFMa+4s78MIxOSOgrFpxnH1YP+O/9zt7WaeBZKUx
50NxKqUcSYY90BYQipMLPEmmkwHZ9m5nZK8Q6HZKNAOLDN5JlnrzUj/tKjuzNvHHkAGiorHPzlNJ
K9qxQuyQFf2Rk0puOBLjKfPTbnhoOgTXjxuDhY4xhYH8HaWpRDNcqw8VIA0/fIdv701hkAe0cFFn
Tw7SqK1SQwpkgmpqULH2tRFe54BVZ1eOLkXEgCIxbQ3CPdrhGgd2eVZhcqnmlq0aqpigGHyVg0zo
RcCEmHROuNIFLrCrfsV+HyS6vvmvwyIJEQE2fJAR2IyS/gUKwxKjL2BDbedIljEwXV9fkU/Ed8Ed
JqLyb9dzGtTQRhoprb/PL30io6wxUuUPgxIhG3hdFP1TEKEh39JUlDPZtzrCQPXTX0qOgaqKVT3m
X9PVig++1aBqnBMn/p+iz+I8PoYhoJGNZTL3wMrIPrgQ8KaI4fW/PDYSMRSTmK1dRwsVPE39S5OZ
2wo5I1Mg4NL0EdPTQxg1sar2J9/SI0NuDecj4rXAeZklNto3MqfsyhWXZwCf6XbgtWX3LdNViI3h
Qec9xVZUrWZtrElhPS9pxQ2ltzK/lZg2YRkbRoHApQj7T4gekf7eLk7tjnY2kwHucMO35Ai/TuPg
NmZ1eDDG0PpMSFpbIBZ2IX0ZGYDdeZsmjr2Jr3kwmRp3eutQvm9ju4/Ey7esjQbwxEudMuZTywn3
BofM8L8MwXETvQ5ec756DMcNXPaASAk4ue62RLGVZ3FteGhzvrSQdvy/szH5kSTgQUArbw1hCPEd
1/rTyxv95JusVLEz1qs7KE42O9tVOP2ymX5ivL0lCNGmQR8l9NLsAuAiuuzOne5plh2pjv1/mwn1
Sk7Fxx2zvpe4I/BKt2Y5hm/AE6dln0kbTGELXI+HmMRvrM4I/1zTm7oKgcXcM4jL1cu/ZBYAA2bQ
vAZV60X7s24g4KMceYKokF1ueJC7aPCCc1AImNaMQ48mumlvpL511on6KuAdiYHiiEiczonZlvSl
jsRfx/ncJoaLaHHXJ36h55wNcq/4jmlIEYTmwqQAfhcqouSwZsTpPMC2xictLh6l3o7L6Mpdauek
R/EGhDe+dRV9Me9Tfaf0XDoH1+QSZM1+gX0BMBUTRVRelf/3u1Zg1nM33daKYzlMXOXaQzGYDh3u
qJWFJ7LTZHHu1LtMRuTeG/rei8QuRnS5h/T90vp4+ED4ng/7K4skBjxWiLdfYbvM+4TmDPTHo6XK
1/wg0TabrC7aBhVEwEPUU3bgWqOZ1ud9UJWKiTAxR51RMQfQM3R1Cpbp0cAaKu3p/jNBSicSyXj8
v7sTx5UC3nDku60RCbBMseKKF1RQ3MopoLnH5oYdDGJ51A01/rhiPLMX9iqDYrdyQy5tKNp2Gr7i
NgOa3rdmcDS1i1Zq2mW3KQlcPUsAGom9HefjdYFc1e48uVr9ajWD2wEqfx/tdvMNcgMqEI+tAmJA
3PfeFi/UgUFktWQUyk279MJ8XzEW29jU4CdG/lNJEeDlS/JHPFgE/ha6RGKLPkrZl8kAEbS2kKdX
UsaubkHhmxovkpUCxOGN3z+jEpLcQVutCCzLvZY4v2UEdQKW/rrgLRWgyBad0NwNEGib0oG/ehH7
5SoIxtfu0NvpGgqlqau0dyFI+9epj4QUEZo5Mpv/B3dxm8SHMywJ6GXD02VSa/cBnbJTWLejVjdz
PH1cBMh48XZdj1pr8LTn3jeVlIA9PQEjQOOyZOadVt1onapbdYPPJRMnz1K4Lt4OXKJDZ+vJ/hlz
gBGH/BUGNJufW3hbvXBD+Iz2bnDs7zX6JXJ6j6fLTS+v+jBfPlDuqnZ8ZIt6OdiUrxykeJvDQkiN
CI9uBEEoKjux+09fJ+X8DARg1VcWORHaelODWCi33z+SPgFaKfqEXNc2wzGwROpij9oSLwhv48Na
DikAHayXZmzA5ab7Sjh0gqHbI4YkhaKEX+TKjsKVGBzuZfnuPfIUiXNY0YbHjstwLAUS73k02obk
VoLQ3ZMcsXRxkPxV8pb3IwOaUAI9XWrws1W8Be0Gi9IrqK1cmKhAiFDSGyymvNh/xPMsYz5KDgVO
QxcIYGPJ0bYW2whj5Km84AxvLOa6o6mjv0Nn+Vm+TchKT27YW/Vd0OIhsXAB5OaR8Slrmkt9CSFo
NyFA32I5Sv8MKTmzlqUYeNr8wMbMzvglB6Bx3WGr1nc0bOQFzTFihkCz/aWXEoQVyemtZvpH4NXx
0eB2cEVk8nm8pyb7mTNTkAMrfJiKAcpD/x71uKB2ZHNgg07IRGqMB3H/c3jjOlMNsZeLcRIZ7sN5
mCNDFG6ZWB65WJePv7C8y+pthSgNP32t/twUahjGge4Dc4gnCONf1naVRcxsyZtdrHDxV3hfxMuS
e3NwaUSl8bZgEzoxUmymufj4+D14bAhHxAGJfPRODpUiBdcJokjgxIZYcOI+TB+RhTcWe5vr33B5
Her/+fKqWtNd3qeqM9h7LXiLCUNBJiVVNZQqAths7D5Hu/WNXs7ph73wr4wFtlFZpeizUkR7eeWG
HwRvhMh5bM6U8T1Fl+R8VWn5O5I6bArZnUzENngzma+c3qgwF2ysEuyKgVee3VS4s39gSU7Vfgp6
f48Z4/Kunm0VRNcY75kBPOMTUu04wM1fL7iK3LGO4yXdLOHV2QdOwCDGyyBYVn4Wv8xeNGIy5ZnG
DcUfExfgCrQ2fwDzDULLb0eCmbvDTP8XJTgmHZooyLNtD/ndfcmguuncvNMOOTxXAYMSwuKshJSy
8xixikdrzA0zqDZpqeu3WGcpM4Pq4HjaqmvR6oXxxUwiEUOMC+F9kiguczQ95L2KONKHnljzhfEM
+PXoF4VWcKNQsP1/fR2ioG74fWb592H44RYo6873hxj9vpVAAZ1tLXL7YRjEizAIXr2FcesrWgVt
aiGu7ezLqqgfOmP8tHNRu9dAf8Izzv3E4LzdpMVZSjyOdzkWk7l8g7f/elaL8J16DK2fzF1VuvQi
C6nyO7cRsiGt80sg94rvekqLYd5KVJgoJPyIJmvN0GlpLdsEMkbMXs7BBNap6hKFLB7M5iKeTL/J
zw4xONQhNETFXYOKw2xe7vZBC2n41MKbYi+toKvaabZjWzwqEyoGPAvZzTm3TZrio/6i/ajbXaWK
rtYXW3xt6b7kpSQZm+Nx1h2pzvbhNI7kend5xbtzPJelT4zwEmBxSOOUSCWjLRRBb8CkeWAhH4VV
KMzmronOewBHwDDfcxE4cNVE6cNSdbyqJFtoNufI9NRxdZxxo9G8ctUYuUsi2UKPxEpsJfOSjwyN
i5vVQPAOB1pf+yBwgxBqbNe5c8nNAQqjfxuBWPlcfOoQ9LHSNGUGQDPSYmQEdHBtS+ys89dCfBja
ukMSDyi8xo5HWIOd0T2Kma7s2iJbrvjUPckWNxDevUPZtuwai96z+HvIPJf/V19q9bf6IFWgVo0Z
NR5u4pxOdjkzbytxnQukcJOn7DcH0Uuw4LXFfl6yHn6Sq0RyIgthvnjZKDe2mIwlUZrohAbOr8sV
43TPm1zbXl7Muo1FWYQh11Of+K1Jh/kNLOqiJpa6U+7NilY4yNlPO8mfijNkhpG90ceLBTnpvGW+
zbkpXKAuyPzosBEbDsKZ84f3nCLfgm3he7ZJEe1axPPzyZCfpX0NGl/Hp6jjJKlmOx/P9Pdg1YY4
qFxISxdx0NzeVaQEqCsj4ff87WJFtGXurjlG/UDKgLPamTBgcmh5SgWre8+oOj0aSlQsnSsUN6dP
hS9qRXdbYiuTnED17xsvQjfwM8mm0Te16SIovqfFUBag45bTGkqflYjXp5hEgblVh8EsmdiM8sXo
llNMszrj3hSsUmfVRERe5Ac+mDyFdejPwXt+GWAVDxi2i+9Bj1tUobHxcpIoySJsY2NcDZikvDTg
BE/Z13RPQm3D1aPu41LhNtqfK240ZAeiwUds3glrhtFgCQ2Ph740pl604qP3Xlt7Q84w6JY7lMXB
LzyS2kcEkDv4bVb1Xw7Sy69u0/isgvkM1H767dO1DIxZj0bmq67mLqXipTmPrIN8zEVwsfWg/fmI
+VW6VaEq7hdIHCJW/xOF7FdkMHuR+MCd+Hif3mKVhfnbMffGclXbY7GybNKhU6KblXGausmQpaJi
NqZqfXCz8xr38uXhvQqklWhu1LGJ02W61w4Y5PkOS8qXucLrmNjxGNHPow6JFmKCKM5QTVRqlZ1B
y32u+IgvoXHECixi60e67bgfu9d3NaEwPHsFNDQj1XQ9j0QoPGngdIgUUtkCDudPZVUkkQOERExO
KxI4xXCC2+140ijV0xdS3bcq6E+c21uNaj2BeTdOuhngLeiREYds75rtEY5YgzoQIz9Buopw0pac
6xgCCO4X13tn6GoQXMUMGexStPVK5zKH+fUV4mw4ll31BouMr2A56AMhpX8GJZIpKWBCvUqPjl7A
7rkmtVF20eYpdMKkvFob7k4/9a5Q1x00gCckHNCbT0ar4HTKFTIjgBxfdwM1WsIIN3AzDOrgZZeO
6pRv1Vt9a6KCB6rEDNqfd25A/CBqCflDLI8QlR+crV+TRYmTTRqpiMf7n5Ps3Jt5MBiHOw3cswo0
zHOfZ7qGm5pfCfJqjjzfsZMW3/4zbwejBYrAly31/zJCPokDCLZ5ci819S4+TIC5FugKC52hfzFV
9PSjmnLq0PLyJ5FX0ldOBWiJpynHuwwuBx74XjNizHowBYzFC5Whv+9Zq8rfmyt29epJTWDq9YCw
+dlHSe1Vu3RQc3i3jWXuZi2bLmJ8aDASB1tMYAhMv3pnyuO7WMkMRtDfbfgjlxmU3ol1nhoD3zyo
YCQmoX9seVAmAIYkSXFxN6MOjl7yc2XVoQM2FhKBUpEUT7IbgfZhJ6frT+pmbPwsCRFDsJ2BMUv4
aGMQI+VxNhTJOnM4LMIRW/wElbPlqMVIRh15D0lH1J5NVWA1uNPnELNSb0YTWJkGNzlUDsaVhxGb
jsVykAdts+ai5wC7uZQiYZq1mWt3tIb3VrTa1bxilBGWD778cOOOZPyKf+3p+cQBtjwDKZ6uXElP
YaRg1wtO7Mbbw2dMbf5jIyt4U7FW/o9iHAkZlyVfiGuvWktX0H5xrbPU+e5aWTEXn0NWHz+8G398
DIOnk9cPqatJq7UNClH0g/G2XWOUPJU1ORshT7p35BtodixqQZQKD4JMEECFpMbgVNFoxxoxFbhJ
eK5FfnjF0S0r0TOWEUmq4BpqLF/+OhluB3q4916nwLgUw6EVi2INTKHLkJN/79n/57p20vPAOfN4
Zjz8SMoWjqXpuglOWhOUpvbQqnwkN4bEZvLasU2Hg+sRu186qEV4lytu+Naq4dVLRcsSlCgqmuLs
ma+IUzMIfte4/mB/KUKyAfKcl1cd3kOu89kw9APgJOHsuOJAu2YKKRFkoIxGwpjsezrsdHwdhQWS
PasSkLMi+JQEUdJ82VbpHNw9u5+JpTy+6HOI0pPrTRvlwPJ7mxuNS9bOeXjsCYBVHw2/KA8Bpanl
ODS9Z45WckUuaVQ/zb+IdZ9OauaA+R3+7SI4k6Xc+j0BYfFS5tBeZLrFjfvubV2bERiIDXzJQR8l
aaWQ6VOuuMiUnPgQ3tm7XEaO/oD3la9+spwAbUijkhS9SLRyCzj9DvRMRwKIXs60y/hPJNn4fTkt
JXZAV47LnqQ09EIPir1pIt0JiI0N85dBo+dg4ZOjXZHtyqMfvHOxMJACDtD6GD36QCAO7v4208ou
nDfU9FuoZA2D0AJMZZdcdcrofrSt82b5ZZa5Igjb15MOIyHFqYTFo1MiKknNmT5+6TedAgkBtwDe
lZ8lHmh5vSgA7/ui4EeWf3V0lw1et2JxbX8f5HrWgttkyRHcEVnlr1eD9JT1N/SSwNFrRoLkxudR
L4Fc4dkq+hW3oJFVhX6xtb1h+ZrsLBAn/9+HPesxe1wtY0AGxWYmTMVclY/YnInfUtAsoz5GraUl
jpBzNTh+c7G7vulvG/jQreGeUf+SFe0cRF8uU4M7lTS1bUkJ+Mf0YvPdnj/ZL/D17oQdB+4PPzxV
ph7h24Bih0B0o/H/4HedKl85UyFzeVvv7Cqxm1dusVU5rR1XoVIg7LMJAHsILjihkS5CsX/r6e3V
9Y3AcyKskyiDR3fmopiaL+1BtNRnt8EjipiXffs7XnKjUQxu0FNUWlnnqREnNxhasOckeiBey7Jn
LAySILHn/qdtqORT1tkJyM0lC5MhamN0Uaew+979xVIbOjd5EfaSegRnMQ756EwJrd7yfG3YzuZ9
q91a4N17aSw8WDqZqiB6ZDtekVBMncQHlzuLFvpxWZeH3dn/oG5HfS4L0edNmaN12gSeqOr/uf1A
SMoBpN0wD6DwJ6J9LAu7a2HAk+iebEmXqY8KUgGyWJFmpp4mSVK0tYmxeVjcmilyWk+utKKLbZrw
gQfJaFPBuBCkLI6s58Vp+CACLMbscF54RwTsCAmHEPqpZJZcO+lQOdkKNslpHSPfJFMgjBbTJ0wW
/8yPkduExhXSZ1v7FT0oXb3YuCB84S3uW5Ndoeamhhn72OOQYI1DhFzvqX5OyrDsH8SP4kT7f3cA
g11pCQn+fStLon/8KJj3V9y2++uBqrneKsSKrxKzPWPKlgCVRmvoWHl6Ec5tMpZwoLMMWmDeZnH9
tRkmoWFKEJcbznF19vIeYiXpGp3anp/3nbE7a37L5dF9QxpDyaESqcGDt2Pe2P50+PXjT5YY51eM
eLv8LGLMgqoOmIAnxJRsGCpUMkxoKxWv6XnMuAdzIin5dk2ITFTiCq0sihop2iJ+bI84n0BuGOfs
jQ5Sdl2ayNJtpzyUKwYHS9cMvqER2gV358XkxV8O8KVRtBWAMoy56tROX9EQKFszDXHA0MpUO4g2
M0V8/wuS7uEFmV1cZD3LpCUglHKu50jk0cpZzQOCp3xrwLdk+UW75vEjTN/pjxP7QDzQLHlHHnG/
jZqkacKrwzyn1tM8ZdqXT7bQdcQJxG14rImSEOANAvvRKZDn7n8cXiBffxnVFQijaD5kNVy4n9mz
AM9yBdMY9fy4jDrneSgsC7YHi0vXZ7OF6nglhNvQj8YFWqb2WyBeBx7ycLAm2VXwN4hnp2C1g+Wh
8opTCyr9vQP9H0nYeF0FoaOf8UZKrTBxFUzM96wPY/Qv3urfwbB7hZvo4uPaDNZSQIatJ2fFUjml
1mQMH4yXvEjFy8QIXo9WweUz3LiplQi2swmx10QQKll/3aEZXk6GYg+fxBGsp97Q4GRENp1y+zZI
d5nR0g3AbKE9czxeKQcktvj5hLu0eAN7YA5Pm9ebesRv5NynCun222ZaHxkv+CKXB3gyHRYtv+8p
6qkEiIv4FMzMaFqRhYYaPQ0QTNUAAUwDHwxuYIUziYzL1aFIwaFTZCd4V+zdq6dwmnj1ryCm3UYu
FHshkRhryQcDTuTvXfNI8CRy4GurHC3+4VaTVI3mPec6hjvsu3c6ftGKcU16eUiBZuRCItH6JdSr
1an83CYwA7mcKapwZfwHwvgghXI+DF+Jlk6jAeefn/937NAPnkhOi6sLs1VKLWE2KRCsIqPaxc+O
VsjbtjWpRPuXTtFD9xPovikZXp6tH0tSslgRAhBNx+kYK+a6MbOUN+Vez1u0L0MISHkSLDGTRBzg
Ed1pYulI5HzPUg/sVc1IBfIarflcAwwEIgqKLQGDAawXy154rrw0DzOtojfMneriUnXv8JKbPulf
SJ2ZMp14+WnShUoS8e6akO+T/2XIOHY4XcW0XZbq6o41MToXhfzkAWKfTZvhus+qlXXF/GHYe1Zi
DmFTr/Q7ylr/iMC/AF8tTN8q3hV8YjAtz5wFgW/MBEEET07S7ATTirrAXO7MJmonoLvSFqEp8/D2
5zfwWgUBt1JQvT4Oaz4NOjgsMb/RJd0WbXfL/PvY9HvUa6G3qmNPpOaQUhFaTqDwsNQ7FpaBu9jp
aFu37m8R8+xe1XGyBCGP5Mih9qP/nPPH2U+L9Vy1ET4RgWHva+wuX2bETMzrlLJSzm8Lcide+HvH
6xxubChbykcUDa3K5fbcB4aNWXmuXTTOLKVe10WlUqR3mvaB0737YR0OyX+Eq/8R1DRIOM+o5svZ
km2+CQX9hDvu4O+I/DdLkpYW8NltjiXt7s4Oo30ZDMT4YkvDjNBxXU8c6FL7xw4rAv8Mu2fQ+xYW
8OAWc1qnE27IbUZMiZfwNvY7YH8NyUKlpXyk8zNXWFmqhENzpgYw//gRMfcg5RHk9L5aaxMoWTm6
++jojVfYWqr+6c88T85VcPYS25IXkBlZh2Gwow3zQBSpwGoV+wG8ygJh5lrGxpK0BCvTNipA7HFf
IeLKhyW569BXEU0TI5nuW8iRNtER1YWJfxp4IzhYzJVoDGLq5TdjOLX3Wi6oJoecOzhGadsdDuTI
sYEccR7SUI645V7P4i4qJohzG4pR1HuNrsPdCAvPcH4VRq5HdSVo9YRSvoqyRugsaErqkpuW207G
t+ltKmZEfmii48fZvkyiuEGpUbFT4CQf7nOHzPHrQvZCjOjAnx39leJTiFTEcdisfcRa/gopwPl0
1sINoIkHgT3LJ5LbJFanPE+bmS9nx/2RSszsQFxCG7J5+SmxVE8Sva83B0iyF3ktsrupX6XLSkrw
BwMcLm9yov884tWZionfjiXYp5S0cn9dULTGo8oDJu9BmpTsyo6qEmvVTqXlAHmOUE2XEsOzcuwo
bofQbB2asgaqC7TWsw6SthZLc/1+umEIsm/REO0uGVVGGPLiQ8gUd8gZtyy7fueSYyi5seX+RUSF
0WlDsJKwLjoRx8zdkgc/0TwWI28DT0cweYp7URwVg4aiRB6JQUqZEC25efHfROQ3UErrGcWnyiI4
AkW0yTPk3Gd90KgjxUPLxQtQlkYidH98GMpNZfaGVb64kNd1cPaZY3jbPYfUBQMr41VzYt/7774U
yOA2sbq0EA7Yoa/0OhpIZw6cjVRN/gb/jaQRAN0jWUYAfIs5ls1oO24bxRyT+f28UW11O4uD1C5z
7N/AQ2iLUtNqmA1cYlBdnKqPqqcQmdfO0qEHf3CSl5epzu6W+lxuLg5AiE8PUCCxM+HvqFXtV0L6
n2LOzH2/ylRUynuzaQjjbmb+mGD7DYvzhS08vEqTnDM6IHz9JpWF2TEHAnvA6kX0tTcuA4tl4lM3
aBbtTpq0KfAVymKLKNeRZBHsIG+E9DSsiR+M+bINlhQcIqZPGl75+lYFIhI5v0b3LdbRTV7r62hI
1zLbwub50vqwfEiy77YIpN6ElBf6vnl3eMVwMroG4uE23avKVrMk0olIHvqMucsapp+ltFPa0HC4
M8ayOtFMNXcDGPfhihtXEs0i5F9oNjDte3kfMQJwCc5Iv1ioNVsezMy/zgghAXiBzwHw/tiIotQz
MCHDJ458w/w/zYXGwhOfzlgSBROsGdUXbrqLbVAddY5pzmWk+fw1W2PmLq9wYASrgM0yWfncZi/y
aYLdurgYFxmdaN2mxNBbsmZeWg5RnTZ8/yKTQY4tL7jdwPYK78oKSF+BDqlQToNCoCcAXkkPS7lv
rQKXN6fbjjk1gypO0tgAsa7x9QBsRZ3Euhu2NG7YJfpzMAjbcdcfDqGXe3Rh2HtB8RSxTPR4OOIj
2FP5MvsT30KvSnTjR7U1EhSYYYlYRjFRxr0WhVFa7FaibhRHkrifvyn/LYSaFgJ/GnDTH52O8M3U
L4hi6tLdYAULxFrd1cn9MhwULbEkhbWiDXTwHiopeCYzAbqBPNnGqimIqrfrcxMKz+xS7CPyD2+Y
LSfGZwi0Fdnaul9jpJkLE9WW4pFFNMFSjCchEm0bttlMIXFJzJdXLPQ5hRtuL9W/Vb/mA2gXWU+5
+LEDJ/Qq5ejUx/7VAc0BJSRX7hutrSXK/Q+C4Al9pIarE/w1YxTSbddVEgPQxNjm+cwD+jyMNHCw
xWFPqJIbcdG/CzFdY5Qi0bIrcy2my8g/TTuQv8wDzBU5UAMW4+eML9q/mngSZDEpNp8gA6C/d4W2
+JzZsqyRjUfLju0cbElHwIT7ej73phuUjGhhBD/PfSeiL4k/n+DHMdDduutz6Ulg+uZLGp7hTiWG
zpjIB7NOseVSkeyq+i/+D0SpQWsEe09OFbu3GbE0Wil5AKZf1ObloQngkIDphieCIhk7yJD1bODg
OBMl4LDp0iXhQcSACq8rC8qgx+o8O0V4PRlSf9mHVvDRkyAvC0xbR37d4jJEb/Bqr74E90OjHKJW
UdHD5nYNqTGxiRZ7qPMIXqNVkDHv99hRfnaUfxttwjHexiOiM71yUmVln1tBQJI1KMK0j1HIsB2N
GU67KoSqaurG3si+FEB6zBnl8GWVzvNyH+z3oC4Ne+L4hKHaVZkHfbkj082YpXmH3pOWb5Vel4nM
5q4yaneEdJ5+uSr3qCD1gihAOhOMkBzlAxiFNcfUzUg1DwsqkGktisp2/0/2Mxj8DaI7I2YPixUm
AoFvGc/vegTuFG4r0cyN53Q0JKZIJMZgjEDmX4BGulibrV95nm1xHGlcUbKaqAsUxJf/5MPHTPOI
pCTvX1wQR9Mie7S4KLIa09pY2DCRE7hlxkwu2Dw8o4aCHPpPvJ3GQgE4L2wMVp3m21c3FfLB4lxQ
WvefYNDBAM7vgeCZO6yllxVobPpvWB3A3hjrWrJx79CXLmvo9qHh+1HS3effjoTA4fYNqrG4+Bnk
oe0T2Clvf/3g/lpEw9zzYfrjFr/KIBLhncm2ys9CX2Q1+yOVq5F7XSLTxDBfFmuf3GjmAJIaDBVv
xpF3XDt679PBS0a4qQus7VeDxGXKiCnxK1lwqQl+upvxmi7falqwlaypYmPGuQcr7Iniupe0KZkC
iS/NA74JJ5TqrykiHrMEFLTbLRg+22g8cOjs92hLWaObp2xuwdbElAEbm0y3uGkqEU0QQA4esFRw
GFd+6uLz65CqNF6PpfrjzGMAblRAsPwHrjcjQEeoBZ8DgI1AQbFKc+0eZBx9JvyFE9u1RIj3EpJd
uJKB9SuVAx2ub7qYQh7YB88VrGQIjSHGdbfwZ0ld1nZyWG74XbeB8h6yfvcu1AJxL6RAV9GYkKEc
Lp9shMSvxm+5i+Bjxo7p5R6wBnH/wZIAjMp5s3zmwLtf+Nu5EkY0PE77t0tyryGqwu0d0oBdQ4D7
TTk2fLMLosMdpfMNxyHseGWUo2rOvDiGjJz70ObxPYOIHoXwBElx6YE8CiLgtgtfoXn4oC1eJ6X8
sVEzXlLBSObRQuXWpb9dp3gTNwMIlqQQAIWe7dCZW53pB4Gz+wQiOkhGMfkcfcj9das0nHPljH/3
LNlxZFRCXWj2OSN8BmJ5VgcvScQnNh54cxr7yH+B10XSeH2ueDfBHxBLykzIBd0EVPkzXRiV8Mre
PZyBx3rYPRhPXGHeGf9gWlBCa3lQs17LHvJYd5XYePrhj82C4dI3NYnUPuJxpn3XhbiiAOS8QTJR
hTJXym/dFmSA8MdQEHISoEEnqtwrwuVXsD2EJWdyKss7mj+q9GZttVZc9rxEdsbbCwQjGuni2Cbr
GtCG68f05/hxmjwOkbOYhVddVdla/mEiHXvadKpp6ShqbiATtvIqLSY6JNL+Fv+DVsso/TDl9Z8c
Qu4yR2BehFkdR6sOWccGLztlNA8GPqmxsToCSn1T8KCKZP/ZPS+w3BFgG3uejzMsWVSsowh0QvpX
Jv4zHvjmlOdF3S9oRnJXe3SBiK1hdtJtQklvFaWhMwjqPWWJ060bWmI/yoNmRTNwMyHo0W8rRW3d
L5Wh87fc3T6Qv+Cgy5Blqr0DbryDHhiojT2pXavzYuBnA/dN5r6X7gcz67l+bjEjFkdvXyOs9lcH
JPmpMPGe2onjVldJICSdfn9qrOr7SjYYqz/vx3ZzCgbThpbvGLHYUte744ugl2VeoOUaQgDYAOen
dhdLujNtT5byW/5+do+EvoF0oMSeJCTQmY76wCHJq86eZzPKacaj2FeXo6HPe/Ca22iXBdbqsApN
sTNb0eU6pEJfs9ZpulSsemv+p2sZzsdJTY/EqJdTfNHbClRT2//jVIhENIQuOJ1yPIj9TwGHQmgv
k1WBgTfpLEbsQcq0Lv1ocYnvscvSzGV34AiuBOS8QxPE/2aAebxXa2XHX2nCh7IbpgOdjzZCLnxa
sI8vsv3eAxfRddo4mVQi0IqAZhnqz1TmsPj0dut4bzem9mCGY0hVA8yog0YKWlMzpJh5DeZ4I9cw
KQYtrIJi6c/9RtaPq5DaWWtSnJxXprhfHGH0lgfeVfh+6UXbZ7vTUbieihBZlHUq9XBr6zqCqQrD
PcVH6wAWxfXdm3a+N64ucqWMmm+5pLeOk5bEHq2CfMVyEGRrhsaYC0hyVbm2U/YNlE+xwIskXkpS
iP+98aiNnVgj9n9wA8xBWJI1xKiH068AVxYIJa/kIK7JoAmrb/Luxc5xxeH3eEiE8Pa/WaI6wGsU
mKC6i5cFR5ZMESOUyEd1UngH+tjSbDosuWGm2d8afxjS7nbzukx/m5NuBFZVwGniA6ei5wDPz9YS
bTaAOnHg381rOsJ7debcVqEZDlLymW/CWNKuVKbuwY5TqBVsRrbKtcGjj2j05yxaBARj/iiNkYTG
nLO5fRtmj+a0gTYQuPsDJ/YTa4ji5PQ24SO1mkR60M/LbxdfQi6GcEwmh73Lw0Z7rBiFV1G1q88f
1IzIQVgXba7A8OIHfSLfYdeB9k2lmNmSLUyUm2y9sqVzXocTxL2I31SH7BWEv1ckYFi8J9f6+Meb
JMC96UiVFcKYxuYfIQvWo1e2TdgXuvYsw6+acpw00zC6poalRQyVXQ4ueABfuYrPcPe8F1huIglK
fUkzcsu6nGZUN6SeXQDDIH33GY1d3HMVZ8sSqpMaLXIJfUwP8YtaWUNWu/gyi6NkucYvtn/ttGBX
eadzpMr2otYimRd1XGekXq0CmowOTGmRgaJ5sU5BaW/jmv3e1kAvj+CyKXD0lmRyskVAGPT9+raz
fCmOVyd4VMzsp94V8PZ/bvsSQmYO01KTnOSCVY4NOpJ7CT37vabuxZp6p7jVNjCbegyWCaqoIoRS
q9pX6vXt0OvG6Hfy2xk2i8LO7o559e/A/w/E7u/dPVvE+siBBunccJ0XvsaVKGVkia2gB2hxIizJ
u0EocGGBVvBX7mnozDsEWk0gAtwsUX2Il65f6myHTrb+Q581AsVfyahCjYuXFn1mnCUKv4mUE9Ks
VVt020p1MCN9NL2brE8vubm7au+ndYLlzcHx89lIb9SfyG6Y/jKRLUY0wUdvwNxg7q72eeAc6rsU
gB5ZOL1/zNIkcuh/MpXBKk+qKrRLm39vFtN5KjPvi47aJTCpiAQeOnjLa58emA08KL9AlRW9Xvyk
bgGMsN3BhSQhBFbDNJvrg58HLFuxZUaS0ixdBGGZAALCT6JFMhmBFTEyg+NTYFyGUzpAY7/Jq0CS
3LgLpo+hs7M+KyY0TDwYbI0IFSRk5JXkgkgVTV9ShjVa5QxS5c3fXF4FtXi0jNXqgbRn+HMnKRn3
/CEjYXYPqNY8TEeMWcvey+Sp6xsuemqZx0DN/qOjJx4cUxhb8moCYfRHihwG0C8SmtTNYEVBg6hJ
O78/af/Lek6Ss3yFgoBMrxBrruW3at2ZT33k+syxjp435BtuPPD3eDCjIvuaH5V7r0cQyTQI/8N7
myf+7n52WBEYKzTeRHYmf4FAKCk6MAYegMunriDJzyvpxIV3wpXaRXclYBCRgCI00a6W6447q0i3
fxlrCIvRftK44RMuuqkCRgPSl2ZKrk3zH1K+RZt+nazmWyFyaEkx3Iwrd0YgwQeCRbJG5EN4vM6W
cQS756rmz9nKfdlU6a/vyw3XNVA/LSnm9ZIC0bw8K5kPk+w0YH8N0Jg/foOhg2YjdUYjcVyOM3S0
eGKK9Lgsa0dw1QS34s0RLI2heZnwvDygkT/1OUW5RpBK8hnUbj0wCT+nL6EJWasfSQtThQYADXOU
45CR0wjAG8Iid6WiXpun3bub5IRo/8g24GhNTkDuTcZ3a9dMQEhaZ5aID5YIk7T03m0cj/Eit+07
nur0uiJ/p4zpTWXHQln0JkrVYvPu1mk+A7usgRnXlkG6DhIgG+l4Vb9frQyGTft8/GPHxTGi8qCN
4xmRHWHx8i5Cx3vVziZqzt6y9UygZMaM5V3qC3hxzf2oPCm6lNJQQZ91D0CUOIlW0UhZipKJrab+
ku8621+I6fpGKM2xI3Y+pZ69R4pVonBFaFm9R07YEN81B1m1ba3tbUb3N+5CmEC0xIQ/Pq+l2BFX
EuaOG0UcRM68ZUVfBlZO3ge0hC9BXvz4L253Uhjdbdp1bRWuPU8VJ/4RPhEP0LpqW0+pnKik6XzM
8LAysEZWKbx80amDlXrEBUoa2vSO/7ku47Jw9lfYjvcce3AKc/PYEA404gi8mzzL800f8AvoPi89
qF3uuT137liPGgI62fURVtOSmQwbfxht5AnIz0i0or1ugF1lVfoi417MTkHAqv21ie8WDPaQFZVA
xYpwdBsrcb5s8d5k/q7+yJVNLi8pK4DDROSpgqGO1LARv0vEAVSs0h2ms2xsIwZLgHe3JJ0risa5
TIx03tW8VjBcMy2knavqWP3LzQBPYlaTjkOk8MEr+hhiMXwJ84tzj45vIKZfK4lThZqc90LdBaes
tmt1lAkMcBAqL6Gdbr4vDoiY5PvnHZA4RgqNR5zXEb2jfPaUviWebvKl9hYTIwviDRYXA2b1OMc8
iwEEV31vEyEUR2kMCL9tJLFKsX/vA+Ji8/rtf9pmwNshJ7pRZV+jJoZhb+8EkgeMapTeLtAerqoO
8TapE4OfaR0J5jCiUCGTOpf8kBADCvU/VrW80cuEX4fGOXnVi9+eWpAYjQiNwx1PA5PfXM9Gy9bj
3knIcc8H5/KxBVdOB7kpE96nSmw2UV0uYmB1xxEUgCyYLZo/2LiY6peBaHASklT/pJZdaFD9AtJb
/JFl9OMD1iXjWuMj9UTMGAK++A/PEcmZI5ip7vK9Z5TebaGoHrxrNQHmatK++aKNLGn+GN7lzDZ8
gToAOfGWpnV4eKP+OSVAPYbwew5Mh0ZESM55gyayDwK09D9mVMb1gZCH6xLcBcR2BmGg2C2Ev1zy
KaEL4IAFcUJsH57GkoMEGVBRfKKnPycCM5dNcZBUuoRh5vEtS8EL9TXRIsrqhAfy44OH/u0o7/Kv
CIVBR4ml5qvpfo31hR7R0Ghbl1GXEM7M9Tn6XVAfsWCBav3I5162LS9lfisZ3tpVzFvILzF+Xz8F
hhVzMomJbMhVEsk56HKHuPdJsVclysTO3Em1RwzR7O3ydeQUSo/pjNJxPU+pL4iUusjb1LhzE7xh
HzsJIRIxcj+dFDWaN0jxqLXvm4iGe9DyxVB2eO2QFfRJwN6O/95cXMcebaKAXZv1H3LyTWooxaN6
cXGLZzWW3MC6UDTWMWyWKz8LLdj7QQmdKuJG1kUwVN3hpTCbuS2JUBR91sKmS9xMSB+ydKAgi+mI
ITvHZBEaSggP9hx1PmwBi+e2hEV78n+sL0IlVVPBODBKZ/BhMxE5T/3DXk2nVNoJhd5vD1fm/BZJ
Snu22g03YW9WVVEjpNdFjuLRnuNBE6I7qdHZhzb3UjTYLskFUQIgTBNK3VkFV5q0zEryqlT+ntKl
6euIU0vYgA8gIFLUQnSxmPHopLKEXH/IlP+F3SwgnNN9IIiGStEv29mpbNz89L4K2VTBKEfz8j3r
MVci0AmWteHYbDYdzbRaw7n1VY32p1BdNAsSCEl3krRtswO80EigOgMkbRu/Opnm+m4xXcj2outl
t8ZWP/sIAHRjuYrm9SBtt1IaTCGRdEK3kV8sPNnS7vqgxBV1wNub9Bx+2t9wFgc+VrQIpLgAYXp+
/tHe+EMDLfL6OMztxo+Pi3wQ1+Gnntrivh7+RkJsZ2zPw2G4GLxIORYyImRP2OhscHF7x/0T/X8p
OX6cncZuMdCAYLEXiwxRxXltxNBaI4NPZe026wB0eZ6b3muQeFNRoSeJT7saSlW7GKVQrgCXpkfT
r+8RHMlJqMNgQ+F4qBR5qkwrXxMCWjlhEdq7Gprqu8ppJKNS5Sj5FB+u+sTNiumdlaiMdxdOkzeQ
TJNTvqWJnlKqArWnSGs5NVMFxwW4yePOpvqaFWlHPdHf4iuNqZcu+cUh3vk9uLz+ChDh4D+1Wgc2
VucI2K/gzZaxmsB3TXZu/UpwiB/5u2IN29HxcmXoBNuE1PSxCnYUiTS7KTSjXDH77146dkQjqNUA
YGRBpVjpKPEB5befGOPQoOTxGB8H/eNtm/D2VTQXYZdtY4TMZm+P76ZkrQXqtu6zx/sPKMIVDihp
/H6Ai+07ZyvCG9SQIPty8BF8YayIY/uVqxyPwMR+kogyNvCt261nsm5afnFtYYYbKwWHWfK9oE/G
7GQ1uvk2OzQRoMV8owSFyvz1VxiHHEDWafarBJth/FAtc47GAIwiXx6A5lhFlaoI2HAiJrEsCg4w
AEjdRsPvhtYaZZtvikMGkTEu6gnK4pm79EBEb6Y+5u4qdIr7P3bBQyyxV0uF2IhNHXVafim3ee5b
vawa0gawv8P6Im88HPdURJ7qLpV5bpu5AN0wo1IvryIivs3LMPUNYwe9KNNlKeWcL9dKVW6a1SSv
SNNh0icy5gNJQzdSZirbDoUA93IFhdiB/GQtXgiMjBb26h0Hw1iHifdl78F2AJmOZqAaCkiXIupG
MQp25hTKWxhjXejYignaaTt20FfkQlsUt0e/ziqeCrQ/QaP46hhbdPZQPEs1Ss5COYvylkrBJDwh
Xoz0X9HlJgkOTKjvMw7xe1XtGRIX8IGBp6zOV3E/ecDOdOXVLvGR8d07SCHXx2BLpP7asZUbBdfp
qAkleBurmiCvQ4OvO6D6xlNroKLKCCyilDAhJC9cSUB9P9lR3WfA4VvfwWjToTen7t+RTYFvD9Ut
Rpw2EIidJ/RgmjNTmEa5/uYzY0hC1fLHBps9H5+l9nK9P+mNBiXUSRi4BQF4wULJ2OuSffZ2JuQL
JUrTcOwaLmRZei5o6kGlzfoxCuUv+N8sJETL2FBQ7aw0Zwes3/n+423rZuPWk+fSDRPJVlsGM/OU
lGp8nmNUMXsl7vqXmYSbHNSthsV74NP9tdaquIE71pt9HRYMxyyarTUJ0qh0qKgwY6LiUsfl4w2o
FzqBJ4MJySaXeyme21Me/EcxCU5YTaH635OOBG17hEBs7iDkOLjN/+gYtlD/W9wxjrSXxhhNrTOO
fAY7Ujq+I3g8uw7kCu6Dot9uGX1hk3Qvvg5+tNPhjv/g+MFqbDN9OonCr0u2NxC52nUdOW4tjCpD
QrxRW1Zpew9IrlnI1JxIhyzSbnvy+Daxnt1bSE/Vbh6YvtZYsx49cWLUw2320/c8yNhgvXr0mFn3
2wdMPINGUkhffbQ5h7e79EUI7c6omuYrb3/52rDARoJNX6FkFv7+r+Ku21uurHGqwQdgJuwAsbv5
iDzWfqtoXjxGlV+ixoQrGA5mkaO8TVIwfIPwVPiXfHHFWQ0+BiRN8tUPY8sNfjFIWp8aAtCiISUU
dKgJaSzIaTeaC/FXhZw2VdhIwgU36izFN5SL5VXVO/ClnUJP3qN5u7E/i7covGBVhH83IhNTIqZw
drAazoc2nxPtPRJj1I7djv5V9Zgf23LIxarY9jZOJfkiB7cwSXMQpw4Wq8nBS91euV+wd9qLXkl6
mOOjZf7UE/pfWRklva2PNz6q1tV7VCNZFEvZQEaZCWvW7fY9i4v5CnHWGDnUjEWOIJUP4fnKfi+C
qvv/FHDtqi0fgsAa4YTclsEOvP6+BN3ndL02BD9toDi+6wlx/svLYDq4gRYXsODJYrqzFo41BU2Q
jROa9+36IY5jI8nFxW3xejv3qi6lGPtmNvF4V0qi4ZKx2pvTwtTVoLo6BRxTcKqDfQtBVKg4PBsw
RbpG4hFOZrTroH37+2aXXF9Yh2mghQIEAnekc9+n/YZMPENc5kADMDa+NBcVafKN3CK42mw2NnZu
RVrbOPVgW2Mau3w49fK+seGRYoqrrU2yUR6TR+m99ANqHTbFIVd+H1YceqCmRYRg4rVuVOMezdNg
k8PeJqJa6Aozp0sNtIm5ufpVv6cc42yhslbOoKmHji1CJeVoPqcxzld3R1MA0050NKmQFh9fDVPu
dTmFzDgtRx1eo5VNwAf3gVveqmEsnZLhkSSu+KaoViBN38UVIcmHhpITxsBs3shtuyL/mWG9d/0O
bUrUo91pC0mFft8kgPdw52XMTafBjRqtJZnzUNEnsayA4Hch80sL/4nx2n6kZxaMxmN5Dyd0iFHm
k7neG/9O7lj+7EPbbzcmfZ7YM1iiRdM9ua+5hcJB5ITRgs8e8V+ZlERk+L4V10pQ6DXWF3sWvQOp
YZv8EnpKBIjz56Q3jGBCwCiHFbUBPbS7DKiTKpJbjEWuHWiYjQTywkpujFfs3ZnZbN7i43oHuwLP
1eKqDUuA+kp1zRAEP1s0l+T+mqxTMSO1wvuR32HoaHJX2FgzhOvvYP2i5+56hR+JyZra2ygPa9AP
P7iNrgGwwLDVDe+q0uzB+SzR4H9+S6zaEXBy4HlEGYSTmtZ3uyLZPuAl9MyFX6RBf5eAS6OJFviJ
B7k7uU3gwtgd+BtPpiFHr9cXh+/qW2TYrjSdLaIJIxCsSypRjY0cg0e4K0VqY5LGZXYa8cRqRCQc
GH1Lyyuy9h/uIzqTXdFsr2K4iGPAj+uKFbo/T+4JISJyF890v51k6kxU99tUDZ/y6MKrqLJsql2r
zXOUKGJCJGwrFM3KEoOCH30AvrB99hy69n+IUExBLE8PzhLxlBAlW1CAWV6ew+xGdJv9F2Mn9nKu
qb4lAGXf/PVSe8fysndG84LUMEcVeIZ99nYXH/QrsATcXoHsi2j7zh7SO/oO3df/ZnBLMLjN9XlI
MtvnRC8LLYb+oxp/8E4Sg8sYNyJBLKf2JyCG88opTM7C3QH42RAYN7iI2d6ZB6dp/GUi4bSzmNXm
rH8ZWh2/7UXVbchmHDrk1T1a/Bq7z65AFr4E0134G99AVPsRFMA73/utmvaqY1JL4Q+rItO0AGkD
pqhLSrk6KdSae9Ysq7HXhMmllRBP5qaM/cGycq3EjysTnSnp1hkHyEivzTZQi/vbN2rlsP1mTR/C
/RZGv4vWBiyrSBI4HV8B8oodB+/VYkPmRbQRW+DsFnp8t7nO4IUe0NLOofnYn0MzBubqt2SMri+7
FK4OvdefJ5I+bgK7MhCob2jVysDfRNjwGSZ0CeqfxfnqUJPo1EOYGbW2SfivBfzNsawDC5bOhkw7
byFhXAoZsORld2AVhFW7KJ1CMXX5jfz9rwhpGwrtoWprovUvNi5WmcSYLxb+NloI3r3aRem5B2RN
TlefDZ6H0ZFeX/HaEIBHJ6YDjJCsbxcwaOEE1AQ6oT3iHP6Vw6mWItJfCAlZg3WWBQsi8bGTcKRx
C+EXkupKfhftb0UDDGwq8M4JbeJf2+UwZWdPMusKHvx+nbrbhy+QD0KVMNK537JVi9NnbYk77iJ4
X73VwF926nCHU7ZacojxnJkujI2djnXf6/Cr0YZ3AUfwrnpFY13ryDL3JFFuz6+33U+qrdcT3yHC
ruF3cHHSHsPbNunpjYgeaF0WkEwqyZx9w5RKlr+laAtyRqKsyhup8ed9x/bnDA8jHq9z4qt4KPQO
zqWVcZqInYlHO6W6d9Xm5aEP2bjbd4GTkeg3ldgdZi65NL3lrfKcrL9UzrUMB/wFeMLk9vWincVM
jRPfTbt3HFA4HWrY0zBdUnAH4foPzfEuXvcW95pc5iT239b70nI/3C5ooxEa176dR3rhIUm8ASiy
LpwczmqIBBRcHeuZ0N/7Ed0qy9e6SOxwzss0E5aU+g0MZVdbcS2Uz6icFzWTOnajR0UGaxJ6shuY
uguGk+YTofmfTY5/pIqWbvYd5DKS65opg9tDNieR5zogpltrFlB9hsIePkWCcAdO3UZnoZl7gmUA
2KvMCrOo64nXXPyfq0V8qQowLlggFLmjqzD2YVRqGSMGPT8nXNZB0GPzu+Q1yhGGXJqimlFB+XaA
EPBiGZxD6z2BzV9Dj3iZMT9f4OkQmmiVoL0XYmmdwP24ivcCx/0sLDXpC6+aIj4G70Nrca0i+UVV
elTpfnFJb1IWWc6c5a2h0p0VgHLL+s2C+2XQ5sgZrxEaHIlMfogQTO84zmHRL24K6G1HisBgTz7H
Ngz0npv8qNrWAx+0z37gBIE5REEryREvSCXOOKSXP+HcMrFLe9zsuAckQYpIq/2k5fzTkVZxdA0M
8DbpuVJRS0lsQFiPyNHYpyjorTVcYXzZP+qzU70v4YXPct0o4LdgVBthE1uEuzEd+Tgpcu2Z344i
I+1Hs5+nAjZnc9ltEfNH2w2+XZYBYC8ePBKKL2CbP7yj0N+HTBPvdgF7oyZYe58Lyu9nNiT+VUn3
zVn8zRtZG7OCPUFY1a0jLt0+Tio31JvI8b39J72PoFN4Jt/pOcda2Kjt9XqT4XjdHhwNaYj0hQcE
Vw7df2Cc0999CKM8dXuCXEBx8yJxd/KxZlt8cgJvV5BuHw4kHNLBBIs1yfd8BZH/37jeH7lZZoNt
g2jASjQ1tcfI0EYXr+ZCA0TU49vxWfkzih39tzB7hxgC8hWV8WINmyhGciFIpwc0AeP+r68Z/F+f
AD0uasillE7umvEX+Mqf74JTCGlJelodUOEuZaasY+vmA+YeL89IWeE+rIaFI6+PJUbgGITsr9r2
ckA7JhgRROo0RSsXrblVvaQD5oPC6LEeMcb3N2p86XeVtIf3IKsdAIZ7rI28AcwjlVDfAuvZnhze
fqxxSYtv3DjR7qrRpOygrvedoFqXWPPKxn+fi4wSzIFga78t8SgoTo/ooDgU8KY64dXpYh7l/Wjt
Gmy2Hk/wL/Fmd5RfFlKYHSREnPWAybROoCaqdpooIZqG5lM4nfWguqjuXVXi+T9WpGSDHc3Dm9tp
nVDmQ3Dq3bo2rKXp+R82o0+FT2XcAaGx3OsRlBUT8EjQkRsYf192Q8A19a6oi3Zq1n+5TqQTzo2O
R8fg+XBm3xHjJUBO+0KSIrG74Bxg1bGNj93HOOrYCxvZMH2OA9kCuVDiwbDF0zRZSjKQqVJY2LZU
B+m3gCHkdbH+jQFpuOvWz5KjIQ6AzoWDFIXpLKVRB3CAdjKquGs8oEr9JRqd03QnhVwWFPbLHAV4
9f2tdin2EHqwudpypopJdkckIfUVnqszOzVQjep5lFUew2WnZDXC+RaYUpreiuapoaS4E7KC5P9D
zYBUBSXIPXdGfLxG5iJmXPp5r4IS2mnhXFagMn+S51Od/xnNy9ZxicUdKiuM7dTv+I5rLh4xp+lG
h0QVKd1id1/ZUJ46rYZpbI0Ey3GS3Dx+oy0CtjR7iuHwUdamoT2XQEL18CWPpQfsjyc08u6LQXI+
8b+vX25j22Yx0IuCjreHd9zKzSE7r+wWqdLLIavFdRvlKb5Sl3cUO6/zlF7BSnnKLQw3SVBlhGI6
vDrKEcg9BuumFzWYw9hwD+Ivlfsew1k96Ze5mVMJ0nMLz6KPNx68PWzC+fomJe7b6jjIENmj9DCO
rbJasHkQ3k3F2PK3rijrX6MYn/0iqlU0jiFniHwg1alEpuU19wJt43x9ATM7fevH7hb/kolE5htq
J/Badwtx6B45mrH2iEOAeGyqkor6gP7+S6HBva3AX8/AJ9UuM0FCC+o5fFnc1IHJsosJIUb0jQqf
hAVkrTEZNtNCES+qH3/jRFJJArCmEF9G+7FdDqaT+qZceG+HGRnH+7tCTJhJGR+9R6pMYYttulwr
/DwGjS/+ufTMatavRs3A9cIZSQXolfMW9A23WjX060TSWHDLLvY5EdMovlXWMX2sK+XAsMZb4uW/
DYsjvlYQ+4MtvGIyJHW7FkoIW6s4MkBRQLH6e83bc3Z3J5y3JcWNI/RmY8SUiiYiZxQdOQeraTSy
nIlD6vMfqs0NpYXqat3027VAIom591jy6luENvuP7dnwo0wo4n6hcEsyMw7AdMXxJ69XunENKhFW
6MyD8yRJrlp/EOUr8450lGzP9QKnNQYiuFZnQtwqqkx6QITEmbpivb4k9VcYZSj6AVEmlr4MttD+
cKZrioR8mpH0gioDlRC5+VUD5yTU0EVRAM7Jl1roGZqCKv9qT5rLHy6dpZZbEg5SVf5HLfdaUuk7
677u7OyYIbIw94MHsaPmQunLdvM5S/bpcUHwElRhK5czMNnogiJqAbYbDLN+oChylpuVKeaUGfyX
+std2cyIm3BAnVOQB0+q4mOPodpl9zoe2bRha1LG2FtXJE4XwR3fmjC4HzjmWiOnpM9MVSPUwGiv
nd7VEG/5f+yDLIiSwiTdUDXjxmxT8RlLqxcbypXycHEzheNHhl8HVC1BaLuqofkZN9ChjOwESkxJ
9yFMiN0RogkbJBk8793wbSf5/FPg5KxS/aqEn3GtJgITeLxmKHvVt6SRMXs2Hm4ZME+jE6oDVrxC
uUvzy9pOWpj1Oet8Uduau0M7LSuUh4cfyL9sa0VuC7vWegCCPsHW7Ut40p2Fifd9AGkc9dZCSd02
ZhCASglg3TdpA6UBtgCjvbVxscrWXHo+Jln6Sg9eFRci2keTkI+CiTo6TaDqYbZmSKRNbscQN7ZP
LR9QJ5/rryHfWbDtuBW50ovMSswmQd1ngZaTLDxIGSHrnxzdRYDYmuvZ9b5FIIl9UMnkKnLW/MFn
Wl/w8tzZeiX43YOPDt2CGzDTi+k94eHsUBRbmxlqhWPnkyc6+RbLlX4r7i5DuG1S9h1zK7YYcszc
U6lYIq+MnHrjN6Awg2lKOwfmmzA26tLNPLxFlNAzimTXQzMUv07haXbZbEfzV/61/nQLUtg2dbW5
ImCE+gaPBye7iDEkhP8tKdpxSEPPTqGVUR9fn/me5Hb45lC19kW29IDQT2o7BCs6gk08jXUpz3UI
/0/fGvbFZN/tTwWaHJWv6W61RPMWQTX+nByKkG3G1W2xoRncP2ECYcy4meKIHbShP6qcQDFvnFiO
/gRXZwnX7S4qFblrEswRYk3+Z85zu9b4MrMcddyzICyrstTz4e4jhu2yzsxRnw/jsUR4c3ebGo1+
+3gvMZBdaeXSljNo/g4Wu6h+Wr2f03PXkRfbTtKgiF4ig5HZU4vep+G+fKNKHZhSct66608scRKT
1/eLxOpjlKKhnjmJbUMB7925HWAjAhaOBTMHn9O6CqCV3vz6hWM/3d9Gxlf7qgnqv4CImoY/slxW
xEmuNPXFQG6pYhm1JR4JfMbaXCoeGROzS5j3j9Vrrs7Ku2Ed5IVQMLXQ5nil/tqy+oGStlZRcBB4
y6ARQNzBQDY9G+xoQRI2Sisn5TvB8YWo1ncl6FuMl3fny62BlI3dXVy2TFD6QJrxfUPP4+6TDWPf
gsCG2TQMVWFJYaOFEXJPVnwZGZQ7WvbAlJ0X9j+YMlZZvLJIkflLAObhc+jKKyMaMZ8XGp/fjJ0k
GaSLCGEQyRFw+BZ/9wkgJ9xgRc9DcR6+6cWUPCMzUllvqzdkfq8UTm51nfdpQfGi+F8Le6DYkvQZ
ekq6ksVVIs++k5g5UzGrNVH0q89ftUt2V96BtjMij8U008MQBUeU7niAliC4SU9cpF91RMRGCyZQ
GoYQ22uTA7nkvhAYbhgpMKdjWPFBaUEiv8MVt7LUVAOk4RYG2rqVyLmIkbPBkf52ZBeHhGwFQvv+
/Sl0EWBVuNtDBjg7auxCuUs5InBubW/MIeK5biVU6v952R0jirq2aDxaCwAEI1eToElmMKdiURzV
dcOhZmYruPhPxh9EF7qJgurOdJAgGsc4Faz0GA6tMsAhOZF5aoOwlbW0A1dlpKDyHI2KwP8YOjUH
KKkdIZuR3WL6+wtu+DqrWCZ600+sxrUTmzPlv9LTUOgGL57wVZJf4cjCVxFVbjs0t4tjWrqPyKA5
MgXDXT6NqeF0JGoW720SLEZmQUp67QBZygdpUsSGYSms7KUR/6IVCoR6fazdV5JMNODjVNGDIK1Q
MmXpmOIOtSEL1KXKlAm+ApjJ0DLcCwSPDCByRpVsOG55toIxCs1yP+6PbHp3xgr45Pu0q2ZcMqNd
+UXMsFxU64MfKCNXsnVUnviBZ5yWFiH0rB7gqX5KUM68Jt5443C/TWvN9I76zhVZQTwkymum+ug6
4qKvNnuP5LW5P6yCEboxnXabwxtSLb1729J2r6jdOmIbFwEUV/zEoqt68RIxBBplzCEPBiaPEHGY
HKF1KHhZFMFRyhOAjvnp/BKi6HwTD9BN+yjf42qqNm6mypvzaocmuZV6/HiTSk2+lwe2bUgnIZsk
8eApDCTvcHtrrTYY5SLxyBbRAEjEWZhaJ9B89wxgntDwq3Dnp1lnRJPePfj1HJ4wwG3Bcim9ZgzI
PgSqPfe9eOKK1Dzfdps6v14Iu40qV2Or2vbTZtmDY7L4HMwm0yizDg4nIZoNOIiYEtmBCgbgYjXN
fnseCzcQ/N4ZM6E9IPg8M8SAdV738d0uaMpCKrdu+D4bDDBKCrdnAx7yx9n0GluybIUebuHwHGmA
Ba4cAxy6xGAO7KgPa+PHHIUdBnutCZITu6pm2l6g06NrKDZjmA545wZ7I8kiCw7Rnasm9X84fzel
gqS7P2XdTMrjQ10joc3amauuUedtKbhprwPDEBZrD4C5qkLDRx+tkzhGkxzXgjkr8EsZHkhrPiSP
padSCfi4Pvx1WKWvdWyD/7bJlINR9tEuP28QaqgitVrFTs+pmYQ3doRkRemGo27GS1J+aHKBIVig
IJvgYBA3ROJFI0hpVg0qsUIKSFizDEv+Rf7w6pI45e+gxfmQprLULryzobNfhYIbIYBRz31RNejY
8NMbSIzSQg4/hB0yseu0GscaAxm0oP7/m4apdAywTPthtjVias+sdQKa2uVRPaogZET8Q02Fi5I/
dSKLWmq4Ti3kJuk+fBZXda1JG23bjroB9qjCqk17XqQ1dSYLrqtgno3MfZZ2pd1dKoSCsjynn4bl
7At90Ns1IH0SJVhYfUlvcqrhenbEsumELi5qj/Ew5nt8BV2mn9bLcaYLsogE62ckholLiA2wMhrr
uE1qeIqakKv/0pTf5CHkMBcvjh8ITjx/zxmyHVOiGjG9MmKua4QG6s1jJCPRocaqU+Iak3lDHl5X
fFXkgdDUTqbq8MAyyKQOmxvLgGQJB99TddZgXKQJ+t+kIu/BJ6+FtZiyw1lQXGMecu207p3KadMi
AJAvjc6xcfSb1gNl75TuexoUys4EpMcnZrj5F5uIDIhEUQLSniT0V5STuasqHcUdbrfKvV/+oLKb
YZGLXkd96JgncAfz+JPYfIxieKGx2mWLUAqfqhIDQLLjNd7U92etP3oTxzxLR0i6lMm2IA43SNwe
Ip2u30HC/X5E8UGVhEQtsCwTRs9T7ppWU/hInkx0rcJwD48Tq2m3HeF25AvurD2eBenjC2TWBDNq
M0rN18Eax2aKQvXPQU/BT3vVp60oBXpo7RKBSAlBxEKP8MtdXPQ01Y02/T6vdvNo+0wOSJgA/M+8
+Wb0LNCoNnklGaqDvQ/eZE1hlWhMFhsxxWXfR0uBwa4w5OWFmx5zP3PH3P9NT/DCrRBPVWAIoDKT
kgOQPSc9XZJ3ZEjLkPbUoluaZncndvwVhdcgUJTiaFGW0LJkKk6TQKbBC8eVXlX6NQjOWNDKnECy
i6xFb46BC+0dQdLI4KdOhexRmgMCidhQZHULQGZKm+K3foWiud0d8erFybHZZQjOfJMIOEsRpTTB
lQnDz11/CgCzLhp3I4ehoyDN+OzfGTN5MRNQxE+kEaEzdp9DmnyAffPT2683JK8406zQlcEaV2fa
Lgkj1TEvpq7nBU/WQt7MkaaVt/rx9cOmVOUxApbymH0ol9dhH67PQ3SlfRIRlHsNyGl8q2zKIiJv
DjjRNwZ99XXO+MCUuY3MMDo3s75AI4W6gElsbvxjCkB4rvq0g7pRzpSIqiZIDJAeTiDyjjR1H/Fc
W2zekJFg5zgBbCmvnOmJauvxPtjZDonwofQuOIoBZNUpJmYxxbd8VyR0zgLhUCaUBjgx+v0M2hnk
ZGIRKO5dIMZA/xKhZJ5pKzVjCi/QF5TVgsNYG0foRfUxp/3br28l9q1Z3THiNMWkHN1+thqqSBj8
+tGFNvZvQI8Y3OrjD0PpkZOBG1yseuQlbWwXaEITJVQr+3rzpFFgJGBGjsPnqifzZLL1UAdodEhi
c8XdUn0t91MoHg3DAwdVad1TjgkBlbKHtj6t+ON+8zbSRNgTUxvGAsXX+LtBhZikzmHj/ISmGLyW
pnVQvcbqYy3gMhRaeil85niFKS5jobQIx/Po6dmKOhW67gNVGen/jlwx00d5tRE1zQN5cbQxq98R
K63jHQgayz5Y5ubQhlHJixQRq+RtwGL8Be3yX1DzXeFI8DqfquTkJrmrSqYu4LA+buLeCuPSpLm7
EtZkS5RyRsfkIbFXiVMPho+Fdanmjq1QfRfQva/Q2/ikLOeayKUUOT5EwACRogz+GnjORSnj2VQr
BgqGKCOq5OcFMnCrEqBZ0wKxPDTWYfWgienJk/tVZIW5dg8dspgYp0YpyNcx2xAlAOvhDezAD4CD
jjmyn1ajUuSPy8oSC4v3rui930BWtR+7FNT1tKZhC7dXJf/QRDA7GKOX1cBrkBChco7keOo6wt/l
TVtWmy8h0tFmJTBcOHNozm3nH36X5TREz64XPcA9v/Z1Y/u9ExAXrZr6V3dPEBI0bn20k86wDJSw
hGUA2Md/Ctxz05mOJQjKj49NwNdFBI4uqNU0wgoxaPX8/P1QbUKC0oisnxhgkyftAd4qXZAch6fV
wcz+adoxjBoTuK8cm7SDDggmeuuUrHQeBwQF/U2ZwlOWkgAYalzFLhqPH992q+Xb32BY9qsFJulQ
1N0KAtyrTCvn8xv8VK7P2k9ZupJ6iIOV8RS0+JJSUW1Bq6pWUDsI0XTbrsSFmexuQif3e+Z/wu+B
E+JxPVSkZwJqj/Kafv4TgquXiRwbkkV+Wi0HltIxn8LAmvw4LvCWq/pt6HprtTRibvJFF/frUfp3
DsaaWQ0u7oYxzv5mcG8q9T2x59w/yiC14ZitrWMKwvFitBCqmJoV1Y7p33age4mPsrgLmkyJX4Km
Amg1qvDOWn77AIWnzyNrkJJfG52d1Uwwy5y2hm3vs6z73uNOZC7jV/t/vYjVBGGB5ztL+l/Eq6O3
N1TeeeIjWnHpV9DtAe8SgZSfh4pCXC/S7dtijwPJ6mdDJ7bIAQxFVUILs8LRsgQpgJyS26Djolxo
vk8XCeFFkSW3vioh16Fppd3CdMULdslc4BjtLH+CErS8YZr74PyA3W97YASHVuXtUIJyxvrFEsiZ
xKebYVA+ywFAXNZr1vjrimadODSE5D9nt6ZC0GM9h6WZWPH6SZKHtUoznXWlzElOl1rWv7uYvBuH
8kJr+lkjIoKKrSwdi/y3t0b9B8Mc+9RidlDgdWklf15EuX4opuzDeiALRhzLKNfUIduaU/vFy7R9
HNCElRVlCBKFiJt04NZ7M6wYVDo640Q0vV8JmIFQZg7BrVBnfts/AwuE1NjPvMAQBUBLwqZ6HkL9
fqJERFcGsGZ2l1Tw/fBLJ8YeVO29fKlTGYA8Y+4g4azySDtQqVqLPQikKg7DFlzaywPjTXYylMbD
jlQUPVKIlLS1q3pZzlU26F/V5n3EHvg/1KATmi/kjbtF5/SkWla8sqSZaTaJxLVN8SqCrKDeLrqH
F0JVq3zu/y8D6+c0SbaajYyprik8RI2p8s++9BRIt4UlV+Gf4w8zukjaXeUnEW074Ocx2bwh0cqs
EVItrvqD1au2Jutg20PNHcs9TzHB+luCdf2LPGp9MdMFRcXzvPx20L4UfBYbfcBP+35ADOdaJ7V6
JouHzon69faXw/+i9ijJNDkGPKdE4RPDj7H62yF9pa+sxAxO/MwBrFi478srRXTT0fWxLJvc1ZU/
PLMgBcXRW7V3QsLagbqi8RXqNiN0oOLY4wwfLIW6cz/XjyROarv3Qz5NjA2Xyhq7xh3InfDk7uzA
Ki9038+G7z7p2YDcKl7ZydvM9Dc7Lm/e9pj1W/iQAOZgL0myMqVAlNgqhjj5lK2CCri3HpR01PHf
7mMMq2RZz7uJYtaU1cpy7QQfOnZWa2ks63cddadwsPN6LphhNUalH5mf+Nqj9wJ4XyXNZShKnbe3
KHx9oz9yAw/jdj66nfwecZ0pk4r4pR9ldFrihWs70xXfVSPPb7W1sgiOWknv4cwQT/f2EjvHaz04
TgpcOX0m5bfj49sOrAdELUBwGfcwaBDckp2K34XoQRK8bSmxE6pSLkqoIVgAuSB6oFmR91pqgJW8
8ZF4wapeEWnHZ/BYqn8qeMUsf1gKKpOc3+fvoxz4nLWzZ9cFN7zHiAWTNbmt7YKN2prxn7po26iC
WQ4VtZuR1NfG00lOx7CJEmMaPzHLGlUnGDQqMOp0Jc13xtouYGil9Lw0XDS09v4U3A5oaA+aGzZ3
i1knimU8zRRI7extJjK4Grc362ef0/y1mIrEy683t2TzC0xy5QpYahvRfjb2G7ZHfLxBHYj/1kDP
TU74FKfxBQ8ArP/CMoRLSXOcInOD4zuAElRIr0v696XJgiwqIHXIaUUcHjN0+1FvVeJhH9ego/xS
s9ObbssdyIq3KNwfxK2+WS52TJhvVzqr8vRdvB84OVECOW0SpYJ0nlvvOZqOWPJF6RvSbXdnL6lf
99U3IaqWjh5soBWEOqOoj0NmaDjccO2YnLIXLEWemrujMgMho1lJJwWSUVQplFhrvXPswEmTpo9R
CAzxDL2KQMoaiezJ4LWZY//rAj1DSnpXvNR6cCxkwb4UpYWdjc2u7ztHJIMA2cgOR2yHq+FEyn5F
Xq+2uJOBzP2216bhmFzsJ3yNMXye0/BPprrlU8n08AwgFiXUBRjtLg+Ca0w+thnuE6+ituqlB2Si
Qvg169IFG7uf6lN7J2g+Lub2xxchTZR/8w66d7A1KmAhSJXZ1sRbLRcLAjdKcQVUZurDgWlyFcnF
rDTPcXNJj9eTLSH0VjxUm+a8a/GKBofB2eS69Mk41ce5EPTBc2a3dH9o8ghRWSGg/SAshVFe7Cko
UKXQNg+2UuY0Gq387adWSAMxq29lxe/mY49SXLkEX80jrjpoU6bwABdiZjfsJdsOnzheJjJ9HY0h
AV2EUHr8dKXq6RNYPkPBWQVSD1zP2EIZ8gtkcZbu8HZ3TrQ+XEbLAWCQooUhGT/yr+T60wmvShC7
2DXNRRmlcu+SfkRAtrBrp2tiSvU2nAKgK+CCpF/XVcexCGQro2YAXBFnDNJh+1PAKvfXP2Sa7mTO
53YMyrpfsuDQRcN0/KwkcKRKpPccoekREEhbJszqWEGvpCz6eJEoumRmdRbuaIaqmjjOPI0v9BwF
z4UzwH988Vmwh/Hqz4prueHmVOyc2fRFtBrjo30nfzsFKksUPt80Ov2BOUxiLRhjpF6WwD0b4qdu
PpFfQETVFpDDrYv7m1eXoHCnPMbATi78meqMSu4+mKpL++Rp5Y825ZCG/MQTtyE+LfP+fczNYvtc
vXQcURMVPH0qdqv6QXHlr2qbyy0nhWShulmRwydw003aE9tf+TimMaA5lBYG6smBSF1brl+ptPUr
nbugHKufSaffXurXTcRC10ut5B+n5P74HWw3JqcHiyHc4qelIVJCw2xpL168TnwiuxYaKH3wLVyo
3vbdpZOcOAwSaScCWoPGlEXrvhvh8L4s8j+8bFS4mEkhr2RX9hjft93voQwcAxz9WWmEydZtzbU5
DJAJM/qePdm4s3jVTtuVU9aERnTqk1Qsc1EgAml2kNCb81q/Ie7RwulX/P8mctQrigJylI51LJus
Y1PLeqvfo91RsL8rjPGi3Sj7zGRodhbRQXeoz5TwH66Fita7RlowykRVNAQSWQwwK1D65lmz7s+q
vbKa7KMsReQfn3xLour5rBfNSiuyIzamcuRzze5BM+wxXUh1Q5wdt7upeBu9aUFtHACTHMlAkfCb
ilSIHog1QCHjWSby9LL++ifTe1O2wGhVKHz/bg4tJLzvBUWV7Ik9zW6BvMLBaZy77TAiG/dxDdU/
9xwEnM/6zAjQ2mtNWIKw0TI6oLvb8oPV3RWgfyeazTOhKuOUg6YHY4gNCQyyxmNr2zYjaSaih/J9
EcncIYUEMS372mEuFNnZUlgj1VCvFr91y1cH5CfGSGyS+rMRQ9+Q5mgSD0j0fpvgu35yPUVyMweL
RmuuYaZ6TKyUjteofWvv6yAIT1CUn3+Gbx1wpNoVH5YThCxQpH6PpQrOciYjC1WyarRVeqVhEpmy
zKveS6yW92WdGTfWCMvJJrUOViNAOJGGotsJTRF+yUbEgB4f6MqXUG49uC4mbqc+OSZ5mXI3ePOL
qxPfhPMM6K2waigq360m2eKJ1fnUS+G3Q6jimWVCicx8FFNP7D96lWxXR1u9YmZXSJo6PZKRZTU2
fVzdyhHlEbsUTQiEvjc4oYO4QqTyX7jjMf427CQau3nJxy7ODv2pG8d+h2UNIy+ovKO/LROLXZVJ
Zt31NIbV8FtALJIa3KCkZYMU5cUKPPIXJ9av0we4Bv46RH2iGRphIALH71COjf34uEMdwMfJ8qHf
dCJ9VSe28buq9imODoci9GbXTifzl3B7dPgZEI4kPEOVcxsGT0h5h/7NixCXrHcBBGCdQDOC7w1u
6NBETYkeBFMc4bun6Lies7WKN8BtxtdjK87Ztraw0pJ9CleCl9WK+aJTsuurIlB3m+IHih2oi3Ze
jkdWG9IPlVzhBfjgdLbqoWWKoeSFHT+4xUMm7vZ0ijRlHp/3WdRTPzl+qL8a/mXD4Ax9afUv/S9X
k5r7aR7qr6Oy9JPVgdff1OPnzWvsQNDBprcbvUQ4UC2MBK1N40NM7puc6CsHhsQBOKhwtuNgP43r
DrHepGr9g/mVIrNm1WVez8whNIcTrUxzSChDMPQOGrj/tYtoiNRx+tvSordaJZqfywMVp+eVvSMk
ppaM0/AcYYkAPvPOy66RVQ84TKKmVeR8syO/Z7gZoPFavAdHPrs04wlsIF0vbQIxApGwROZwN/3P
/whGHj1FoJI1Lfy0NcEVCTE7RPS45BF8qeY/q8QuPhJabPhjjZ56Zjz6jjGCIvB7N+ggQgg/H2Co
U6eJuRKS+8kotvx7zm+4m+Is2DeXIsg0F6/TCQVdhiaowoKqSQdU3Wbe582wDfSNi9RNMz+wx+US
ei8DLerY9UC2cOdRhV4d3ZDB3s2Nd+WBR5LOXEDY+HxUhA99D3nHcb6JYgV+VbacOyMH6lDaP9vw
WOpZzpWUTDvFy73ddJCVITclis+pGlOSx/+XzJlVVpYArxbdb1SrJOaATBxnTMZCkid5Z78OYNbK
U6QEtAeyrsiV5gqTRABuLGO5ewrJRrgSbTh3FoV8hrL3O8Lt78Y5zsSCE/u/xZQ7CN7nyh1cWfNj
insl4NFIQuxV7jxvPlMTRb52tSO/Gc5SIOOXc85tUox/Ftb7X6whUNfRdCOpxBGH/5Mh+1tV1a5M
ArHQdDlx3J/jgZkIBcjtQ+kv/mAj88x3+67rEm7oTp70aaWdOeSMykCmK9ejwbkZOt/z62Ovgjtx
fRhy2f9c96P39a0mNiRlRW94nKTsHGWZ9MefExn5CjzTFWt3/YYAUlbat0nW8Q9ppVuh4rjPi5dr
MjeOC8M0DXM549Za2MjygEnlaO1cwQuhrdNkWmJA595GiQuLAd3x4aJLGUShAgKmXxqxhYONlHOE
WYHFsjmdBfHEFllXIifEL1N14uQq5UvAo5jlVRyCWXPmoQ7UvL8A5PUpVWlN4KZfwXxRU1wthSfR
4+xGZrV84JyZ2w7eCvDVu0o1a9WdxpPAAsgK0ZMJE53Sf8eGregkxTZsnTTvjVlLcM6ew/m0IMRA
PCAYd5rhHDq8iTPKhKvzcwX81jbZJAi/N4t1xVh9eiYca3wsGUTBnErBfXYCbd0JUPineeFo/wGY
+RJa4FpCbWwDa21vmCkC+He1wGKu/VX6CII8avfPHjYYSirBoRY8WwCHO8KamWkvIo1OW8TWbmPL
DJyQYUVsMD8V4JBySoRq1xqIEPcvwRYgpTAAYShpRlLF3uFBmVPQahL+rU04+Wc155Efbv95v8Bq
9CxK7YlTWwArL8tga+hMpvaUNW/9eXdySYTCSTVRkZF6nPC66ucdGUkCkkr5x1+sNY35H4hXbMSk
D4IkXAm6813SPIbXn/pGiYX5PiTFO/z/4Ne+Z6uE51LjjxDszsQOOUm5gmjRoTjfVUvIvw5vhvBJ
i7mkDE8/14VoB/kOfuDFM3E50MaOoFWlAbXymH4BXi/meu5s6dZzNfSYQZOdJx0Wb279c3KLytZ/
rlYWKwVq4KA7Txpru2JB1r/onyU7pJtsgbs0Uq/wp9Nu4s8ZHMmBsNzHBvnpu+LnlCCstY6JFuYX
oYkTfYEr1muPtokWQPDiMEqEBxMxJX0AnU1r3yJE29/DZv763xUNLbsZoMrQ/sBHZKHiSe2+HHJq
ePpFM9AgoGpeZ++sfbSN6Q67X5kjVMUBjHsAviV7X++d5yrLdxVowjOXE44w0ti9QG0rlZ64sZxU
1D4MjG7Rshbb7/INfSu1hih+NrmlPo+3iXLcvjpwIvuKa00M/VcIcFvBmyla2nvC+FnrL9PfYZ3f
LNVIvggc6eN2zGhSPzblXuRwn4WXUbAPsTVay1WlQERNvsVd9iI1ToIqbucEXlqJBSIaVl2ITNth
KuCdlg/3TvmjZHIOU1SZPSLiSDsWOenjr5O9a+PyfsMYFFqyjNZrctmJ+Lz7iQ8ZdGlbu8KHn5Ss
3jyxiCEUpruqIV//O8rEgQdoAmnuO8WXFgttV4j7rJoCae+s34PIgKQQdbpxFm9rL63hj4h3M57t
5qdYAhOUhqOcy4KkYvKEzxsFk6F1H6lhCVMv7YIyICksfsbkX/PBxFpHTE8r1rtKJ1loZTbuiuWN
Q1uUZ07YrI9taAMAth1kMG3hm8Upcv8V92VR4XMMHNEZ3bLZ6Bf3dFzuC75Li/HD973ssncWOPKP
mxbtzVV5CDHrYGgd9ixmyD5E6JdzUwfTfDuz+WeAKb6ihszJFXTN3qCa9HE7+oXqjKq8YFn9G6Sd
mObdes8ckjGZyMtkIVidbvrfPm7iHI/UA+2ipZGdwJMHWLfEcU9dGiixcjpw2cbw9TOmcBDUlwG3
oG5l4FG2hCEoNyYpldJ+Y2xju6CQFbH7Cc+l+TauwvZlu1MttW96JRC/Gs/z/wyrkB7+app5NoT1
W8WvhVPCGrnF1dNKTHjff9YC/6awlmuS7GK4NVERujve4X8mBpkEqAHcMdW2WC579zUfUMKQ035n
jJI1cwLnh0qpd5DiHAJgJYlIYG10Qbtb2OjMlp0A4e1JjO7NfS5THdWaXU//M1x8Kzk02u35Pzat
ejl89QGPqXGAgRt9tM3Z+yclrZEtQNxfaVZH1g+PvZDsg0DvLW+nZHrmrjPXkFTDX2z0Wkt3McUk
Om1ycL4ItwImt2mci4BJ2uQTY6Py/qaQJowlNumtsL/MckQmPFeIrk9M5czql2VERcmCCRmmPEjK
wz8/sQKEaztDxaKZT+Mb+/Ncng5CmngeUCHBu6WbnQXX971tBHl7x0biZl6EKljWwrOWv3j0lZyo
z/mdb7pOyf0dXriDkRLVd8SuUd6/3UvgU3sH3D4JjGe2ONJV5intuV7DsFDQnTclU2zX+OEQ4WyC
kHDDrr1G9hSLp2Z3KNu2KFyjz9mIfgQhVooirPe9PBTXI6+nY7GPSu6T8xvimMqxU5SkBAdQdM5N
+m/FwhwgXrHh1+YBnNJaMkTg3tpTCkqX3maXCZQ5Ht9HULqB6WKBVJnbOfYOKBAjrgxnmGU9TMFg
dvFvUvEFPUR9lDJr3b3nQR5SJiiUxJaEoMphZX5zvuJAYDUQ5oXvvWseasflY6NPltnU8PWl8pMA
vpGMqTuuYLcRNRXam/gQW3VX5FrF6XIQkjJJU80GXoifeCstwz54vnEKXbo5pR5AoKerlv4zQOuQ
xUFx5bDKNzRGM7atYoxtgc4jgFDiUdCeAsmtimCmKedgEmbIREDbP+Uyh2j9nIhGe91gKawHXkGJ
0coYFF3r/je9n+OZ4wlOrHbpcFyArCmdcy83rH/ANQpWs4u2HlK+4++vSvUeoZa9FT7aul+uJL5Z
jbKR9+vZ51MWNDBcw8XTBgKlq51hB08wknvcvsN7VAqwvPdrrB+0nwo4mGizwIMHCfwyQJtzZtdG
upYkHYxZQp+ccU7fG23nTpa2pHCHSRyQkA1/CssZ1UWhCW9S3r4olB7IP+IyDz3gk4V6xxH2mLDT
Rbn4w0JgXRcSJ03HVNHIoez2v92euDxJppr/8uhSznOdS593ficRWSlCPggqBOL862/3orZDhIKZ
u7HK95UySCI+St0g0UlA/60HfO9CslQ1GXXlKhS2dEf9dqhE63bKxYNLzeQ+zAQFYsMdrQPjUf8c
NpAUUd3jWvp4/5S7LFVvP+fcXm7dhCQKlBVPPsApjLOS0ZUzuSImOLfyDO6awruBG/yfFLHD14xF
YvRMFe+ZoYZe9iEFwYsFZR6yTNdY3Ttl+s/OInFD3xmqLhBcCd8Ps80HyqljD6XtnQSxfHS1s33h
evZaZ4KBDC5ZDsPFyP9vkf40qMeWqAQATOpiIUTVJNBQLcvhkXkn+EgnAup9sEyvhYQ4L/cwdxCQ
FoWSHDaMV+/0bYNoVrJiXb09hII3/g9Nq9yCkBOV9vByTKQKEkEBZj4lAG6lzZYqtGKUuSxCZe/p
I9YuxNDs5gJqcfeFJlwbB/+3z6H+i8XMpYIxQAyJjz7nwCpYEqKVioEXyYLu3snqNvuS0hhpQDJn
XNTA+mK33hj2FOdtMy38tc2v8GD37ULQ/0en8OvG0PxBwy6iYTayqfLB4Dm/zNantJ2g3GFRl2jL
cbXPZs9l072Js3IHYPneqgwF+ijHaDt2gmrYPcAnTTtLI/8oGrhydPESvMoKmpE69PGmPJTm0hi1
HpsGLI4Z6Aa61+d8UCYneKehL4YYgN4B/hVoC98B2kMKk6frMFduixDdISbFwIU2TUmdKzdu9OqQ
ew1Kuy46gofwOJmaOvTeXoRRRAsWJvLzx0e8pSHMesKTWghGzrDWRyZ2K47R4jD3nVaaVqHM1lGc
OzY6V0Um/+1cGNnda2enWJ9UoEsZPPqBdN4tIRt0a3tuoW+kMGof2DDNSHUSuN+PUJrKy1mnfrC5
D/aBQmcyj0Jdo6+P6Ep2enEqeDo+wxoDp5SlV1l6kbVYmn1EDjZasie6NSYSNZ4813M9GjG444Pg
0+XJNY/HDaXqlDoyO7zO30NqPFf3tMLFpRA3ea16y0AONE+8ZFySG5FyLaFWT/z7ArS8ZyAahn02
p8rxF83GrVJlgDTzAlFWA/GE1D8Poq9iX7NSY9dPKA//Kpdcu5g0JZDFXjL6znAkVMRNOS9/QF4M
wmTkxw7YfnYQ+0dhVfi93xBy7BXQe8y0kJEupN15YUAY7Kcqacd6u86mMaRH8I+vxlrbPRuWWHCN
j4xdfwFlgEGIls7xGysQavfdSCcH3BRuwhZliOl3mgmNLtD3pYPI1OLhdm9RJO0/8ZxAT0InqqIV
VsG7TZAelgHIKDrSNoEtNUt/pubJwVk7Aev6gZywi3Hfc9c5koVQ0dJbIrjglqOJDSvcWbUiho/h
bCGT/b9IL2t97B4YKPiNzQpJGZtP4Rn9fUmYAC+8JeQLPuhZ/6uPawS62YIGcupGdQYY81jEbhAl
eqRLvlL/KtORWT12m4KDGVYT74yentD4vYjPfRl5x4r4z4U/inTMcwWvSqz1yaJULjvCLiU+dn3P
tHutMCFdHP7PnA/98hZO0JhoomJiAIMb/E3xjt/hHiw+pcC3WxEhxvAnMaJPwja5cHiFbBly/tys
J5qplkqicbVERWVl9naAG2w5jlO+yLcuxIGjhLckMF/oMM6CkpcAaXPeB0JDTq47zIlv+63uyIA/
RWLH44TrQhVRZ0a0nYEez0pEbUt+qPlV6mB+WhEUSVwTebzTgwRvgNM1AOTrnIzYaiqcZ8GJ3r/1
6rtn61Y6CSGMzFfDgWSuO0c3YImLf88ahP933611JvoGoSLYsqbXgQq0rWwXq3fvoUqMqLwOF5sQ
8Oduy4iKtBUBNYLARNFvoTekLYUnk/1GVRPXErnrT/x4GQMsolQ5OIIeQrAqXrYJ4t7q+Pey/9pc
/J1TdRkfOgjBb2liyc8cyRO84slhsxbhTuv+DXqk/vCboO8CF67d99ciUVydrrQ/2cj+mBNawxsJ
hE8Ht4lnCYh4/bQgZBUIBJrIMl4iWg9phgbFt/MdAj3ckveFY5OdRstt5OHPsvWn83sZW++DMd1Z
b1u175+iWZ9HNjCEB+UgrG7U7mehbxVjMwKuiwQbp5gdwBVC+lD3Q5B4OdJOKrvuLcxcdXSZVKfn
1bNUsyixZFxUzpWqoEd/7Ga6P3miP1T4DBfQH4xShsp3Hz6HqZyuQ6C3Bq61HuF7r9M7fLwYsjRd
IYOQGbQ4gDfkrDttBAGd8Wx0YfItHC0y93Sz7YOX7224JMQiirufCmnppzEVPSM7MecfZRPy/gDL
EOo5T6vlXu7mD5WIPm8nPhIZV9eVKt1bX7Y5UnDuLwyKLJQxZ5mRL+1tUUnfmWwN0nwEfTlY+p48
VJQXsxYE4rGyF+EYBXk7ptw10vn2EB7MQB18yDeOCss+kgYkN7DDjh+lggJBUrhmixh/2vus8gBe
4OwEBvIy89kn+0JUuQMS7P06kZRQGs576wSgZWaaJG/VyTyCfJfjxw8FSZqmqI6H4aMe9++NPr3U
2SBpxOtuFQhd5aX0vlqXALittFqD6dpwpq7Nkr3b8OlAJOVemt2lKZqb3x8utuUzaQcyuXJCh6pI
Z3WP1ypZixtLtWeXyU8DNN9RuvLM+QlJj0k+LiVwyXG4oqpPboIxzjSu/ZaRt7igYchzYFtJgSPM
9OA4HnLGcdAUDvFTRjhyiuDNWpcs5WWW41cIKNjoDvMNldwKwFaUHGi3IXg+HvMqHmkZAQJMpCMu
FO/5//l7qF+pW0eWOm8sebF7l7tH1hG3HJelFqKSj/vK6BDTIj7pPc1+/aim1iijkP8T8wk6XKUZ
pmhh/CYD70cDBISxFQI9ztVKSQY3dXTbCAZigfvBlC84ORmMkJFUo4CptGrRgeZ5WsS6njpRNmYA
TtdDsaEf5eCSwxVDajaXSIxG6x4G91ezSFBxeu5XUByb44Yrpxiq8vcFNqF6K2+3uwnbSwpS8815
XANmWWXJryqzl16ueQjB7Yvr/ihKQ+yKUcd4hCLQiTbRIDYo45Hneg9AgMqgpbirFvHr/vw1908f
2jgtDLo+iPG3mRQc6wWgCAysu+0pTLPPwAuWi4PULYJ1H1kdo8HIbi5oDJuxX6Y9kLGujmKXhomv
fnpoQm/rXfAEn0WuEIyCDxMRkx5YkZLFmwQ4yTfZjxvdHYCvJDVgk4mwHactndslXOkKHIZFU3Ab
xnSrY2/glJUaOaY+pcpx6YnP44IlbViOcvWOs0FeIOO5tfSONQEydtc/fwZRr+ILizTF+q62dEVn
3A92wktUzY40qqPhhZQqKdYomw0mzFr2vXqbpxRtR0aXMgVQQR7gZctfk+RnO0LGH4F+ivugsZur
2sz3qACfSDhm8OonSoepT9JYx3wzY0W0mVPTipfvU5WvOeljVd+es6HI92I4Cx4lZdP0hW8ElgUJ
ZXX+lNjjqnv3HhCTcVGBAyRirzdPgNy/ypC8cd545JPiH/QoWbm2r/dCcs+oWFfcEBA2NlNZecpR
6eDQ52BzeqSPRAMhNRjt67gqOtIe4eowDMTSdNkK1Saj7oeSYmBZObfvBM4wjQitzh5GhY5DlyKw
dNWCpPxExDPk5qQpwADInPNR/gzX4giprMO3SZxuNuHLf9rXShHyV9t9TqYbwse1EeMAoB3qyHKh
rG/LuLmoxj8Am1oM6kRoERdXZvOksWWDIS1RaON8YL9A2hxQOsCB4VnC1Lt8Zvg5+ikT1LfH2Jp6
V7c1FzTyIkkDHBf5Bb3LXSsYsXJsqQzhDGbTFVmiNgRTg8fbXdhDiVmJdgt/OM30gW4ihKtreW8x
K2QVTHb32ha7d/+23jXvUS+7Bg5WmUCTQbzX68ugSsSihBFHe+7mg+rmDV5q9gVEGqZ8ZE1ImCD3
1zpKF3yeedywjz1yU3xsO2CDV7hZE/vwD/bymmCX4p+lNX79YBXntwK5y1sfzMAD4WFAbRIqxT9x
FQRUsgtoqqEfmWmTl5jG6lVIXi5x9+x7LIcbEvDQUm/SMf7QIIAhxs7NCRYPpzgE1N5TAnuPSyqn
82OuMla2ifx8HvIrte4rm+zrpnGqnl4UF5U8QcNzsX9e5kw+pto5O9ZkN0Gm2SwlKlPdOFgMHN6k
3e6RbKNHnq8e/KzHor+hiJbmuJo7R6f2wPdZJvbDnQuVaVN+OcfcF3E137VzoImYCQYKVdstSmow
9GBkTnha24V39mdsdt3vfAZ+W8zJKWC7gJMXBaliSSh5Gz8OGEuwiT0Km+mY8ZdHZpjJjYMilKLf
TIgHXJAzgD+KdUgn87L9RU+cS03M7DewAJoA/rmV8quQj347K5/eQ2LzLab7YFUMwm5qVnvkuKOK
KdgSYMxhZssLMioCAtRh9Hyn4eXge04e+Aa0AZ7fGiiBsiE+7NJ2VYL4eHkx4PxKs5vuu0Z8Gj8G
txQ06WU4D+Zs6wjWLkUEWEwv0fV28ZnLHG2mxR1k1H2SQCjywnt2gHWSxDPZTUEs7swH4jlTX251
NbZuM6cpr7cgQ0wNCGJrZfiHYODt4BNdo9FzPuCMf63VX8t4CmsAk/szEFhLnBP/bWopRhkOnqsl
YecaHkYdIWblS9kBD2PLuHBmsbN/lrfbJfh4K2t+MkRvEtgc4Xlcadb4LABOAGPSapAtYJ1qt/Um
HNBGlC9oTddHfSyz4lUfm65uUt453xSEicEkJKuo9wsGVR75C4ftCJ+6Rzduff2kf+ykDRCTlnUT
e4zUWMbJME+QvGYYWgezrRnn7Jz19Kzt0gLLt2KQhmkhJ0uLgXOkZhRedi8AqCkKQNhwcE5/Yzu/
NnK3yHhBsvNRILPAzqQmYZDlEF9rVp4CpYwHoYwmEzlOOTaCg3k4OUC4rQ868/+awiiPVRHMQO3t
vfsEtYkVticIwCwcXLKZ1b7NvZOpoXc9dKCkNRqOEMw9FoRoTeHJ/7kWmR66IIA9TSMkFg2Xlh63
VIrdvU2v/gBghKjI8sx1+r7ppDT473Dh72hacKyv5Tq7wk8Gr/DOsPEoiQrJK31kZyyo+qZ6XHq6
6ff8QBQ6I+BsNWmm2zGv6ZxgQk9wzNqzrSJy/Bpi5jrzZnZKcJCDPv9KslEZTRw0C638qFm3PuDt
wOlyvwbx5dwc7ikGPk0s7fKJsBYP7iUPhrR+H8Or4Cu0OQKY0hDBfaYT6Om7USHjQPJibdGkT9uO
kvXqA2fNzmEG8vasHp1fGl+q7qqRIrr/xmQkPqPllP/n7hjRM1HiDhB5nsZH86FC+gFTGxVRqM6Z
Cu6oQQQoVGrX6sq8LJE9N7Yrt6vcYjGtIblhmsDB4441fOUwqxMvTNdcwmgJcZ6sCEhNaBHekxjd
uC13G50PoSr0sxlPQrI4Mtw0WnPLyx7Ov3yr3eyzOjZGxbWRM4burXQGgrm5wakvbhD/LtcsPUtD
jBxvqBHzQnImh5oJhsNpeOdpPmWMSpKSEHWsZzIcZ6LRnqmDkZ79VSqZ6U3rA1EupkKaCSN5WJNu
wRuzs4NjXPXV/10Uf9IZyZP1bZbmClmYav74ArjWDLqXLSHAuaeDNuAf5ekXoeIYJQsM3grjn3uO
5hAweF2rY5kBVFZf/+Twqw4TYrlZnl8eMRx93CljhFSWdu31m1hvTmGoKHtrnnaY9fjWMsvcyNl7
1IghA0s9orDwQJbfGWMEBo2wbPnp/7pQZF0mNndn8RAMLKki+RIIvtj5HMrq9wGbZSBXqcSv6kYW
sKE6zNKZs68O7ZAKXSqzV52hAqv/WthKZ15kztjrE0xE9OgAY6k3FYlAS2pDU1Wthfkmdy5CmgYi
3oUVP96xcgpz/JlKTJU/llKO3kRCR3X5R2SBnEcHKNbv5F8lvojZcRYp+rci6+ceeCiWacYOWlCv
SuaMZrh+L8i5+8zviFLAo0fumzHjUxWwYED3sX8j4a8zbIXXvEa86RBIZmhBsb/UDnv5O2/yAyNQ
y2boZSC/atSLyVitEEJeJGdRq80hfm5EFq1PfKOukGnQO30AOkPJJx54MvTKr+roDzdRCYjuXqaM
3EfhYeLgJKCOc1NdiV9k2agKpo7CtGE40FauFvZBCjIcAJR/nCQ35jNw6AMJaVakIjZFNx9GP3jV
OLPisFLzWIptMXNNRW1DMpmVjUxpygAiDfkA3OxHcC0/1OF/sEHhoLJ6uVtaFSILcMHm6eKSuiuv
VBw8Cwn5ZR/Ikqzbrt9se5GPAoxmdmZASzjVgY3y+7flwmdFUp+BxNCsPtbn8T7FfFQSz+AvJpmA
Nzh4f3ilp3kOqtplP6qVXgMRJeQ5p52JqyQT3NV+KwiQpRQ3ut/TaIjd+4puQHwdK931ONZ9AWhp
O1irsAs/Ay1V1h4HlxTnHlkf7OCHGLmuNW6iIS/Hwt32INUs37lNDR2hBuNGWbIwa/x9U+XJj1U4
eMddtSx1k5A2tdJugyZwV31n+rvtCMNMv+wnzLIY6pzYvX9J6L1RUuCBWqrL1+++0K7indyP4jBx
R0qmpe8+/iRMlWxZfiskWcRj1tX/4p/DmFyIGGx8czWjM+KasF8SFjcNn0o++yQfc7aaj8klOIHG
F8AGzIBmwiBE5/7mGrdoxWeqNNOQ3f1Tg3Aq4l7sLwDd7hijE8B7/wznLqAbjgBL73+pU5tsAKH9
s4pZdS+mjM6OvWrWmfS7t4qv0rAjjOgAk5kRnSWHOBlMSoJfE49/tjHHkeCCmaDQE2L1DCltPxci
XQHjwqfBUsfYMjL1PZhM9M7w4F50nxchpoytip2yX2WtsuGBzMCwaLuq8wg+thcTYCRHXF7GHWtI
Y85U44tjI7/hbU+p+mR1/2vfjp29Otb9kgT0NZx1kGiO1TfMzuJBs6RH+H1baKLBPx3OZE73n9Qc
RwES9bmvEBkzXZ5MZiDt4kPz2DPu2X6dRtpMoZKDZhOXdRlxGFSKK+QjESaH1zCAg6V7Cy0tI7M/
nj6L0rBm4XfxTHcM07mUf2/j3+pWBIiOFF+63JypqB0TXdUa6ilTTOkmt84+fznLZyBc0emBTeS/
XIWZ32ugSDTzn436KXWoMqeSV9p5QB0+SqZwY0Geuss/qqE3os/xhJtx6Efp1+zvhj76rdrmwHUS
eOEaZkiYK5w0o/CJCetBD5YQD3RXuqzIuZmUO8gtOhGJu3YoRgMvGPgqXx1AYILvnXbx1E3K4m87
aCcVl0qlRkWzbymARIOjQGZhEihQvPjSnWWvIQxetLJmAnnc4bjUukFYcgz92P9wk15dpcpYk8K3
RqJsVxHYl9QJgErLPZsV8s3mHmrfg3hZ02+N/X1V3Av584vEL0rJvywqdVTQepDaDadtb7yOSuPo
LyBAq2tS8utXlh5UMib8v7xdxLdD8nEk/k8yNYKAR5j+1vp/jG5NVyYLSCAxlW9M3fOwitvz0j1R
CaBQHWlE2TTZWcmgOF0c43GH7MpjC9wJJPq74FiM1ebLc95tiIkMvWngePyiRFGV7LMMBlCMyhUF
7+6ofefjKPyr5TjWoyLWKtUhCFVCUW/AilGAusFBZ9xiLqpz/W+CiFvXbo8MvU86CLpP/t2cPC43
VTiucDemCjWo2qxFHHtk3eXriyyOS3uRD/MnrPOcd+q/PFwN0C5YBO1y1xrVcUoFwixzEsPzOXvQ
rqekGwqbrBVKGYGNSyIvT9W/D5WS6kARWm4CEo2cSIrShmCmvoUczZdaYpNOfDAw6DddQrjiPTHv
3TSn0efR497b14gH0SHSNewFUepo1VquRQM4hYpqmid6c1IOEViSQoylhcJLFWdU/a14alAz/LzW
+XfUwt44FhCJllJNBpNNe/fCsT5gQw2bilnF0X/gzaRZxAG16l31UsgfhJld/+nW4eqn6zWC45Zb
oVR/Q0zak5MBZBn/JvLRTcTSBFi8SZvXElpiCZllQ2wSfACUlur7uBD127kQeWSI4vzG+8OMqXEF
8kzdl0DkwilJ3HljOlXdXC/2SlJ+q/pAjfRDiMOnixLWb+cyetmEtaNv+gPvt152glkY7g9WCmqd
Nzt4hbjLmKFpc0yHPCknasLbFQ4G/waA2bRrEG4HqHT65ZnUIWpLm8iFa6PiJZmwbGOt1oqV/W2s
fX8p19eEBmZI44nCOkNL59X76M5rB/GbhTbuGKOvdrYtmM36d4bNZyEITLPSvNwF9BQgb5SQBSDA
jjPNDatd6k0GcxlU9MClmNT9NtZB9VYe6UseGbg8q0hsp3JHPZOM/K0T44PgRxG4SpxvMvY32Ex1
AZobZJZc/tH8xGz4USp32Hasf1hLIKUU2bYc8UhWYwV6MQXSp2qp6OoVakOUGAvr4pa6k1ybN//t
vKpa5rjIzcchNyhmkBDkMjGOzCUxO6iJXRls8YN58SSui0BAZw/azQ59z1zAoua5fAo8TpmG1qgS
eidyHF3orZrOWIs707Mbw50miJq5ZCtrlxiXl1eYwriFwtvEA97KOiLo/TlMpFAIZAiS0JpEQG1l
szVCv6KhdIrm/9TVNk0W72oxUgMUD5GYm01/N05FGWB1yjt/+8vy+4/1X9L9gsa/TglKFsOahINM
ZdB1vhdzjbsUPxD6TFMX8WgjfGYWsLEYueO/HHux2pus+/eN3GO91Zz5Is3nFeWkScW5eriu5Wxz
HGi5L+GS11Y+6JSeX6PNgnl4QfxU0nBzK8cEGpXp9qJXDFDFt3wSmbNaJiVJy3noFDYvpjRDMYe7
coHUnKv6u0Zc8day2RwUkS4zcWLov2WFtMLK+jRTR+oC8vs2iQqMvtm+Lp/xllxj9v/SraWiLJzt
p5Z4U0Mt9f71hPuK4ghFsdUZbTgN9uyyK4nXSvk5tlB+IQfWL3I0CLcVhAlL9K+H1AN+QnjkEUnO
VMLhTYlkqk1dvBKnKLcQiGD4vG/0F1ZgqCwdlQzVYlxg7aPBhjJRiRfMVvrRTSASpSGsiTf2D1+y
PzwaKkcjprZo1cCSAnVabVmd6t1gGAh2QfD4CE9j7lz5h/pJj+lG91FN2RiZsaU4y79YifAaU/Qj
jINfIwbxXVCXjUCzQ2s0gGXuvD7s/vJ0PKyKKIxulMuqkiEL9jSJsvihjqFAEIW7oEFM3JkQmJGL
9Zx8emSrkHQmTuGCzYUJKyrQIT//Hlh2jGDerNHmCYVjRVHc3kqGJBQURWlLge/vn/v3IO2TDrlU
s63VGjsGqiMG+5dqFNrA1sEiw4xDzZQRpZhdEg5oEnDvOuo1YiSnHlj0AYvhvsmxJ+hQ+cEiT0Cr
xFQWML9SKa6x9bdNMWsbGtCSVu0lwu8Y4Hxt0jWCDpgI8xu7iy0Va4X+HZQKCx1rikoH1sFyFDVo
f2cN/EBpYylrEQXO8fP0uVNBsGiegWpD0W/QY+KEXpM0Fs4JpqJjoV16/r+9js2odfGpSiBWPZxx
RCaX9ldCx76lbyOhyXQqaxaqOPWJC/+WAOtkoSdTdSiATUUsump9Sxjh3L17X/rTroytltr+6M+s
mkaMlJVtj3jECOlKwFZ9mAHbw9iIFet3uCp1bClB7VE7lAhNhhDkjQju1GX+exh0R04r7IbehsR0
BiiSCqGjGtLMj73V+BlJlYJjN8Aln1Nv09aZXTXd4Srx+LeMOiXMCXNLyG615VQdAgdIYXMC1WRw
oEdAbhzXXuO9F9pKUepn7csEAJ9HqG+9bO75GwmxriGlHkZ4z/qDe2KOpC7Jq9GE75hZvfMucHwj
HwEGlAxB9Ax0KKtaFt3KyE/I13a4XwWBltAnP4eJfKTa4IqcOoxjdyAQobWSs6mILZqRkgGxQWIn
YLiuQFpB1T+zSWaAVhFhp49jsd8/N0zpfArQO2rKPVAvs69CxkNrUlAykZciCgeYZ3j6srUzAokO
lguExqeZJuTvlmUItxNjD+fNWQmjIJ0d+XfOTRAjZKLJiKVeDFjvglHoHtHPTRllvWFmYMuwJVy7
eITAqtEsRsIjDcQ4vio2YzfCz1HKMPoNghGG9+hGrFzwjows1ans+De/IlHBc6B45OoiuesIO0cI
F6jUnBQhzHsCBGo7EVFTDyKbscXqE46dKzWAOi8VsaMT2VmxNU2UbWQ22oxmEqSRetEz2aQIGa0X
eFiN01fFBAT7XYfMoH52xnAfLLVtzf+FLRjaIFFRVCTlawJF0eB17ObG0XgZLJswKTiDaCHPeuYK
1hnNgH7mkFUr8JF+1rDCCIRRNLdlQattHrCBaR+TlIlEgA/eVQQyl+ndz5Xd/J4b3rvFhuBJfeJ6
l55ac9M7eYz2iTTmmZWoHnNDp6h1neLIKcTvOcPzScww8xdCOp+ytOg0hj3Zr3KsTUZ+n5HHW7bM
KUE1L2OO+WW/t5H1MAOKcGFhl24LyO3XisHoyPX3Zq3SPtXqZUa5VpkTGOF8M1sQAf/rPs1RHC74
4F9a0+B4Ybkfom1eBbtZqaTDXkNAPy79PYrTptZmf5M2088uH+pz8LTN72ZRIvmDnwWCINDdcMB6
mHZoI79UFo2djg/h5uom1QQQdPpeFExUzK3kbGWgINKN82gEUij3Li4TQkiPvAUnYqnSOMheuznI
gnoFkxe1HsBa+jv+iC9xwfTepaLTHorsAvAQT+BZmohreUE7pFjXwRqLoFEPsfmujLPQnB0CnH9r
liJDzI2F4WIgeMlh1HamXSnuggMCBGTWzTncIwaWyLHuRnTcLsevvaxK7Pr9b9+Z2VoRBwFUr8zx
dNAm+wFT1pAlrUV/k5HwNdpB1H3urmRDbPeXfuhPcrroY0jZJtbzUr71NoaA17Vev8rNCRPIy48N
r5/V8TnXRBsWSaFQaHqlV4WrOPL4AX8Nn9v6T67npuuF8zgKr4QtZTBRwnASb/XVfaoiC2nhF8Ca
U/0Ogo+LrXChEAXez+MmwJH3WfBHJ2LhqBeToJUrW08JWf/ZXQvEP8ypEHUnGMUgok3tv/RPdBtM
p+2dRfMmVSe24jQhRMBJYRBv7/rOvEjx7Itj3NSoYe5NRNWJbagPtbrLHKihJGML0SB7wJF9HRSo
AvQCQsHKL6v00yo0v9NruM1DbMQuDa5e2zZkGIh1Rlj38IRqYa3zEYVoW6EezAczou7EL0C8R+2C
1gQ7Edl3TKGrniLq6b3q3gP0t4c2Fm8mUx5kPhnyIQ7qnySh0YFv+93/bnepdhpMjbIuJp2M5aYe
1KNuRdOYYODKzoHmXXhVes6zCfBKRrEloGc8BKx3Z1aC0avWnwpFlEEl2QPEGTFPqCRF3aW1Tks5
9jFK267GjENpkx2RWHfnU0j3EaNR7gNu1J/GLND+x1aBWnkZbMG+UutYp4jm/HsbYcR2hjGSUpKI
yeyM9/mkgE974FZ2potH6rvmmKNsZHHy8L1A7LujLr3w8oDnmM8Xqx99e3lac4L1Y/rfEvVqyPST
0F0PYVoY2BwajH8Usl+wa46jSeRewhKZ/wJNYPtVCsiegopkC4IVqhb7YzjKy3iNg3xFTo7lmD7h
6w0dH4Js6CrK65jsXU5XIMGoQBJs6lbvyWKCXSgG3rpr/LdY6NRgTdLFZkgAUwX3Z/+kj3V2iTRt
O6+uWCBoHzxG8mzb9W5F3uSl+aFCQkA5J9DpFIpNMO5YvvDgkTsqIV1ex8gQSGy2/DLewhp6kj90
VM6pCypxc78xxmJPPNCQ78O2qbRAJSwQOd+YmhlGsZ43ytwYRDNk73nNy+/oO9CR992LvqkQU+m5
csfhOWXE6YVHAz+lSc148VN2PyuEmnyNNt5EA6iOy2cWKK6d7Ry0mQ3RySqvB1eycEEbsJoE49Y2
RmnpqEh0wEDi6SlH2gmVXqCw1V3xBVMYqPRw17EWuEjcCCaWWz0jHD3UDHK8dJa/mPErCrPpy148
x03v6L7zykdw2GafrkQT6g1x5pN9wR6T76nLH4w+DN5Tkve7dyEp1PKymdNws2VqcBiEAVePNi8V
pxg0C64W4c7mmX5fbnXbqODsQzKg4r0BZ9/vURO9Fd2WL5lPcyf3lgghOE7a1E+r3Mqn5qvo2jfj
81cRt5ytnJrOQOynopkA/TjBdDIO8youepKh6TMsJKvFESZdIh31NUhEXLXM9M1B0JzisXq1Y5Fq
Ct2HLIwv+3l2e8BrBpJEG1mqEb+yXtEEbHeCOht1OEXCEQI8Dr3VCC0MQ8sN5CD66uVTlYAO6y+8
8FUBo0H7SDoJIKhOQxFTjAFkDvh6Rx9KnWtOc+WQSa6zR9oLXZvflf3sxB4lncDoeVqyFi4UA4XD
3MBWRaK4iwSMWt94Dz6UFUrw2EuUXudOXIGiwIxS9oqhAYEPZQ49HYAVI+3ulCZ2E1C5NwJRMSZo
yHKuwgXQ0OcqmHQrxt+unqSS9abraeF8wL/HNfvwgrqIeL460oNSzeAMhA3uKef8gKFGIqcoCNc9
xxk4LlqRUyg5l0/Rvk6fiqaSTn/4ZjDrV+p2cVSmfKc8nTIVQ/WUX3wyxP4MECMDREBQIVkSmEU6
cApdZuXKGwUoHy6ARngo0aVMjO2lS4xr9GX+qu5UsTg0GvtA6k3s3wNgmfIaDmrvjT+EwOJnwbwC
tKZTl2Y53jTBlDJtJzPzKBVa72nKLmbpQP1ZY4BiydhxuY/FyG2r4eYdA8VFi4m9Y8GOoEKLpHG3
Y0sXGPqYHOBRYIiA1rHT5+9YB2fy9LHkd/Las91lQYAZ5i15gzbunsSHzxUntpNQe99MLbZc/hOa
9tg3FVM3tl3jFBcWS9HnXHxzNu09eoMiSrbII6cmIZqGKLol8ltj2a6sUD18ImgNNRs7ZKXYzWVO
Y36RkXxUV60jLHdkATIcfdmVhGiMUMeMo9uMxnRAd/J6JYzDITLoUhL04XRDSoCtfXViMD1dyY4/
ONTP26/qpWbRFi/8mB2Ir3UFnUT/aD8vJCNIJFPUKJWNug6IH92HLBTxhnbhTzgHiauWZEj3dU6m
D5Z8U0vuSXIv7uT8llSfefJ/JpFDCq4neVxDdw9qgj73yYqA3P6+n1Dt6+I4dL8rHlaDsOm01cuw
eDoRmQYzYPpYeAvCLwvY+6RSvt+SS6XjHxxoDVGOom+u3o1txKljYVBE/QRqLQQYicRJH/l9GK+B
mkbLhyXj46PDRXUo91K37gHENG/TSFy1HE7vMdhZWU1zP1VlK5SYj3zrCht7ksCB4BeTCsZqa+Ss
45cFDXH6Rf0LkVsJpjm+8lil4u8nPV46OXfRjGm04He7oekjXIdFk/saISU8lsJO+B8AkByivz7Z
hpgBrYfjcQPJ5HnBqdSsnE10xpK+57QZ7XEN3YWQ8gzkthuGCBY47aH+Wjx7LlJPVAm8MdxE5Gr4
7y90OcGnEoYMjzcZ22Hrh5WiSzg2Q4A5+j6ktFZEM0yWxRX0H2A+MAw60TbCUwjf4pk9X37b/7ky
CW0Wbc+LI4nXVK5YIXB6D7vAg4xz0FH4MSDirSFbqN/GyEwO8y5iSiLpcwk66UByI82Zsgh7nH7K
xJ/QqFPVz1IRj8KOysUDaz6msgkLPALtXtaG5oKO3yXaR9zgYFrIVLT81fTf2/4ZbiJDftzAl6b7
G4oHcGWDJM+57Dy3DGfO63O9u7+ry1Y8i7szLoW8Wz7ln2FfDTyWiXBX8yKaoCVJCm9tZlhwyPpW
oGaUqMQxjMLwj2a6rROJEUTZlkEq4MPCJ185+j5u93Uj1f5TlXdoml4yMhL5QgBFLSx5mVJRiool
tOThyJz500dC6QaxudqHAtrsE0aP/XMgT4ZLtNV224eC4GlYEf/EzT+FPBxV+sdIl/pTKOkY8tso
1Oa+JCCQ0lBL8Q7SXsUIbd8UumlFACmzcOjA9fcfm66NeHo/XaM1ofWJ7DqaGAxRzFR53pU4KfJM
tLnI5DeiOGG2LpGURODsxWonJMXo9MAfIFFdgUCt/BEOjZiWS768MaYTGllh91zl0hsUdsYTas+U
n0ZZx/ldLKFoPEvVH5hr8lN5McMNbKxyrOrEKdonUnygvdvH3clPXy4p8XKcK2j+2gTYic1HZMeC
oF0xGVdF5QOLLqg6mg8UuF3NQz1K7+u70HQPsnDWUvbKtx654Vv6/hiv02uorlsIJCkBPULZzu18
pfd0whuEbgThocXzSG/QdEGvWU+96UkGxiBC1lJVYR63dkrs3x3uC5PIj/1tK/8+FUeK+Dg1TDAI
75pT7XcPWxa+GFI/2MTJP+i35BU6cXdhTNBpaN5t6Kq+/m0oHivwr2biC9qbgMqn/F7GGAsJYjKX
bKFl6oBqiwzLasHmKyRGOE5hpry6dzQg0IC71iNZ2dLcOmMortY/OUcBzA0Nd9eSfbK1lnco5ta2
ZTCRYHby/bRjhZOO2jLTR80NkYBNPKjPgRudM/ZQqvYce2rHuqSDr4RqgJHvnP66nCxqsbFSw9FO
l7rNZ/wSlV93yVTt480NQkfi2bQ2aAg7JHUXn6mDIaDcaQ9ZcET+cv/fTl+PiKavzXQVW7Bdz86c
9UN5Gy/l3opa6Wo1zcsRP1viB9wX7hXhmQeI9RlH+/1etwyOS8NcTRtCtmozyA5bwAUi+3jStyWM
bzCOIkSVYPoEpBvW32Jpc2qFSmz48pbR8fE7Pl5nLLCe9MWSiEyljlFPcLyzqtNK4Bcpp6UDNTNH
rc+TKpaqRsuvciQz3YX2zZZnBQKsgztujiF3Q8UidyRCr6snl2BVDKtnVLiPjtye5Fq5ZZp9yGae
7/w7FngdXf90FJffGwe+Y9cv99OvM13CcVXZgl7+mOYLlPCVkLaBjTAoD4Ir0W4fvdUtHD1Lqhiz
8jOOPyU0nh6Xuyq7QTdcG/fyICUyXsmvFlGJnKnOgmkSK7pHDwA6UIl6YcyoX+PuoYJo+WJDBXBl
RjsNuboz1M9pNsK/qU5D0nP2Ad3+rcZ8ZRQaurDyxKDjkYMbv33Ngr6goXgq2344EcjCLVbiqgpq
nWlWj+mlK6isKMc1+/ATamOamCkX30Hm4QKsRqK3UCSyzRzbl08YXkeI3hRV4c9TfdCxrqbyIQpJ
TQ4tFRPoLgGGeZMVzuz0DIVTWXObD3L+VVuxvoDmlH4LChZMGPcZ6/xUKWHtK5itLkBf6Zp6GYPq
ng1Z3kYUa84oyWIzd/rBSr+l/uNRFR3EggSjfY5fKlzUl1BN/8KiltQw1hlZkZJfWHNxr3MPhIqX
hkUIqeKR5664QPfOI+Ne/TEs1+vPJpc9SuV/MndxGXGJWg5PgakiMGLTLVXlHy1jaVI61PqT08Ap
uKxmHwWjXivpaDnQu+RGru/24EEawLlCQlIKBuqip/fUj/Y+ojS7U7G8iReOEEG6i3NNTT5Btunl
rYSaoe7OR1ixucn1De7/MRjP7hsDfwawCGJOjN8hDgqtDLw5D7YAkVnKIQbFHOsfO0PU+kR09YCE
Q6wTSrcdH3jPiH1jhK5VZaLClfV/gptGAg6VniXMdrgUF7cQwB6PlIn8UOAxZs8ij/L3Br0xHxl4
S7ZW4s3nqq/0ieDd2R+Wg8+yz8uryBWKqvsMhepiSZaZLTvq/JX1YlbyektDYhCAJNM3X3GCXVSS
3iYMA/5ywIztWWKeTfSnh767ikLngAalLyfntugnbz6rj767cCe09Pbwvvao5nHgKKmGcjZwM2er
xFE70Z8Cn1c7hydarMMmABkQt8VOS+eYr53ToohOOPWZrSPFAtW1nxVO9q8WwGkKUZdPge9t7BDZ
/JEAe1slmPPdr3vgY0meHk/qtDEM4iixn6cIUtwCC5gsTxxEA9l9pp9psSZQqXLyQrKLS6FFQyUB
7sNHo3C00wHbjtX1+5db9xUIfREQs+TTplFZZuPr7GuhgM/Y7lKfJ66YOGa3Hf5hdf5VY8ifocEH
k9/zJeSlO5fufK2XQovcfWcenoSOV5KDD6N230ZBxsEh/werrsdOOkECeowqNSZzwlLrbREoksVG
ib5hWdrrhQokPuPzoXSnZleQKyRZKKO7wUa3bZxLMCnI18hsdyi0ViPBOStUkz9WoFhg1rqTNRaE
0vNPDJQTuMPYWP9g4LBx8jf0PbhExUXrp42cXdrv0FRJ+CpF4JMnGYZuQxH0oFwmhtWObDZco+tB
TcygJ1yeMVLbrldWCW92/aROrMq0wNC7hvoWsFFVB5KjHLBqiM3LdHq6NKb6u//ut/EPZ8Q3rNTr
PFYCUheTcNmtbEN1dzQCR9ps5LaAn2OjDq6nQ5jWPA+GxmJPB20DwscOd5H5xP5MJLXooIgBDdm9
EoCXl1rNhuML/l87IkE5S82YNV2oCidSgFFEOD+NWjnDtKb6sI+L3NczIM5aNztZ8M/Q/44GRq35
JcVpH4heMNe1UGzknOML/NcX/qX3PTk+3+rhrlE9cgKhEW1tre3s0+/9AIzJSSXTwdE+OvBzHRJg
HgeaP3wB3HskrzrKqK3pVJaRGjcf4/sQwGv9XrNW3Y5nwiDbRQTXDwtsx+dW/bEzToDU2lzwBG+S
z2JvluFlbPQTBs/AWyi7W9GS85n89r08FwUHfbYbCQM1tbheyWXGFSMIrQj15N68lIhHqLgsgHEo
z0gmzUZyiVYcZrKMeSmF5ld3xSic2zvRSLFIBKODEEfP6fkeNOMzP894x3j/X3adq2uKcrjTDiUu
4exEwaalEJaBbtECDaPLnVOGB1w3v6mb+vpsyylI0i2d8GyGm69y43emNtk0yT95IjR4XUbpUFhi
QAagWD3ST0A4qCOnkiL4aWSqdzf4/Q5jRNuF33htyXeTBNDRYsteF/GyHm9M615XreKhBTv+hqcy
J31pLaznZivsgdAswz+NFFI2eNX1+XepRqD+RtZHNKjtlyfXPtghoKcOCevYaHU1XqT916lIF4+d
I9fXvDSd2L+TWF6+gKj2qZXXC71fiB2g9xwYcoqWBpbah7qanG3v5VrIGhggD2Sxy9KvvOYMKNz4
dH0OPgD2N8dgyUwhkAfCbts1LY5sFLEinHQtXhIvVRzz42DphuxkNLuQj0sxI2IYCDq6J3wvou32
0HQNqI8VLxJujQBKCUCS+akoqqBmY+EpMBjBsH+qwxRmXuvhGRUSqdDJzbs656cmzPCeXR7h+HGT
U8pi342MKPq9Bw4MThGYA+HHhtNjoDx08lZLYXl/FH+wJT/RmxhicZUs7/SYSPYfq/SO+CSq0II9
dHUbwyyDTM5E222b6rtKKjC+QCNuZdh0IqTjlCSDVzV1DaRtqCU0BozipIx4V3FoCXSNPicfv026
PHa6kRmySVTxuEb1byvX3uUZB3M5b65dxz8ZcUDUTyau+fatU9pWFhc6lT1KMv9s3OBNnsfEu0zn
ZHig9FUrCB1SxAGWVbNPMnqidEv7aBLNsrZW1VpKaWiTIBzcy21J2jvSHXyTiRywNDRqaXOUtJu2
LYC3fPbhPcL3GneIbYwQVBoVJU8LEcbs0VBmpFhsZjdP3mpb/gAhMJq4NraaHvH+Gano7QYDX8G2
49YvpHPg1puDG2DZF667QQyhSoksSdqh9fiIQQ70THEO7sjb4SjNHfFjEyCNUDAZaTNcSbrHnJuF
pmYVE/t4lS4JCyo5+8/YRkMsGrPTdYzDdi0td7HUDVAPeRrTtuWZPgOG/7sf1kN6cai30dtfYeHm
avCU9QGeFoUCrACjNR+ZJMeA0j4icFyQ0+yxosUIHAKH+hRLomB+jKziTne3aNujpYndF8Af07Cz
wKeSJPo6ti2iK/V5lgZcoXMCgCQtBv273xr79YvewX2lzgkNV63sdW2PFlVf7lNKL9f9wAxiMhM0
aywwshiBye/4Kd4TxazvbzybxxvbNB7qE4F7tmvSIffhFXeU4zq9eRj6zOwUbuDFGkd0ZWkBV18T
W0u9OHkRaiSLL9GkwQQePsSfakUsoOrqXVZ8rpff7CDUO2Hiy3P9TNDNcF5aLpuTf6GHzQQotEJ2
6J7I5iSC8itg96emVgTZvR/cApGcNiBqyYD6/j8x+EiIEmHvX1UUw+l3CvcChXHiNEqHIQ/NT4zO
2WmCf2Kce6VuFOlXQJBspbu87olIZDIPv3MUkWcG9pxj/0u8nedp1B8y7BmczoTXbYULQ0dhV+YG
yXFuxWNPR3R7r0VFTSmgF79esRXWviOo40hib9/8OxR4vmvSnI4GT2uXhzYMHmwrRe9uOdTYCWfJ
aao2zYLlIwabwwbccgHXiGLDxxOqMzaQLtbgCJK8wxu1/JQnrbZECAkCOvdkE0XS8KX7U993v6vL
iV0xFisFcqb0rlQDmwm6I9p73qha0Hn15Ie8gXkM73aCL/tS4YfqDdLmsE18OtkZRT5LE1jwXUEM
LPt2le3WPDgIsObrJJ6sDLEs+i5MgXnIyXC2PYHA1wyAWneu+q4aPf3LxHKRNqi1/dRSle/0wwCl
+KT3nf5JTYfMrjPXvOMWgpc2tG4DVLIC/qq76Wpu33juT14BzjGYan7UPQ6MpGYu96lwMDDk0Lfo
g7Itkf/J7HtNOSRNM/S1ItCbqOiTpxqsD7zuBN8wRoAC6Y/peIpxKOusDzqWRD+QtNUS8O3DBlBg
CeaS6orGo/BUdnP+EksLlk1xyAABt5cMSjNA9iPvUYivYIAbv+zl3seICZfcSwlrPm6LBee11ZBT
+Y6lWGIw7hvuwuIgsUwXDRYiESzm/Ke8sH+tpaPJEHPvnjV4oMsPccak5nHJ4dfIq92eWU0BYlCA
qnymox3Qs9S3uMByeemdGJGg/Ch5rsT/ya6WwYwhZeX9HvJVoHr0QatBowxggj/VryLh4hSrJY8x
yhnsuCyk0HMIKIwS6lyXE+wpG1ggNcbVAsaP3jhMlH5tuvCOd5nNunn7NMLC2ZxBmIe8cq7S6wFr
ItSaWOgztE1rRLx9dLikADxkgufoZQoaCoJ9IQLMxIrVvorbGkhD7qlay2yE/V84arsTad1ZuGXN
QpZP3FgyHjQKEc3hFwZx29eYnnJOwKHYmhxs9kzhN0daWdt5ekkTP1+WEoJlq1GcJHZ/L/OEQUqt
TQbD+idvX45tBsvkQblmxxvQt4Tlya6IwSbrLr14FJ20lb+MYC1UY3EXAwpQQOFLI2KnmNGHIzwK
yMstjDmvAyhf4FtBDH2gSWpRXosqYQOM3aJWT5Z0VXJDPDTSMKwGwIKtASicvbmAIJqpkVAV7CQs
D4Y2Hv9tpehEi5RIbt2fqPpuks969W3XAKipUOxCdE56gFJ4x0xlvJa4zSUfzFgzIHCHoiL5genR
V16bC3ez0Uu1VjdFAUHWFXE9wiiDvJ5LPxJRtzXSWihNF9/EWab1r/WgE+KKijyHUGw/zZQhDeM/
+42ZHxp68q8NI0Wox7QZFFfS1YyfPd2tGgv0SWS3v+0vslRj1GoFhgZCxO50NaoPa/KFZLdMxqkx
0Xtb+0EQgg0YYkP8VqgDN3fO4heW40w2uFpNjgRwzawlZaj63N0YSHd4OZSpQPQLBQ6oIeDrcFRu
D3K18jZz4Bn5ab+virATuyv6kNyEBtVfmAK3/8z7t9MtCw6UzS7JD73+qCd3MoeIRFjYErZOcG3w
lsESWJI1yYkZcyr+usan3eJ0Dc4aScta6CFO7bwmY9TGZMIjGdab2Pni1iMK1uOqu+a+cJZWskm1
KocO33DXHFeEPvUJFuQHbXSr7wtlF/1UdjsZmK2HmT2a7LAYro9gwnyAKghkrw7411/61HfCTDdV
RqazkpwZrl/AFrukc/phVOA+LT+i5oTBUvkoHC/L4RuZ6w73ASDSo0dHjkcRb+5EqY3MamPCVX22
Wi0620bNFMVIcPFZrlSWiqU0drgs3IrzlSmj3optHYQxuM/x5alktcDufe7QrepfQQa5jUht+VRE
fBxMDtIHNJUbbhIEejSOAo1J65wVEd5CGW88BW35DTjzlBsC1G6DA4Ab2on7cst0v/fMhW2dS42m
SlA+lSO5j3NmTJwz8WRXJP+mrfxpN0Z0q2CM4fenjQm3Fz9s/cKc9vjgn+/wAwvDtUCw+WnvJPJM
IWStS7bDfFMTYr8+Y5C5GQ9pjU65zBDzwjIzPGabPW6c8hUI1jNEj/+USStytTejQ6E+F+pWtg76
Z/DM6mkOhvU4ctfz4mudU8dUlpABfE7abO3s6Qkk0P7JkOkIPouA9mR8WVhfKPoueVr55/nFl81w
GecbIN234SORO6FhnPAYX/2gEDzjIsGwu09LMCPfaxwtdAT80TecrSQJhL2YPpAuL7BXo7zeR/cU
jEIeqiALGtJ6Fu4o6iEio5W74kf19eqJDiw30PVhPiXoBmx9ErU8kFcDugn2vpr9iu7pKEXbK5PB
CERdao6S15ACBIPgLgpBr5wlqgjIFTeot+4M25a2xEl+wjaUuLreXpCBmgSqcC4WTnqQsDdBNatU
O/Lqugrk4kkyR82chGroAovtBwo5+B9ZGW7b1RtNV/P7JG4P92GRrUoX3HwDBkPk2HuzmvjKfxlv
YhaBCk6FNT2GPdOY+epZfZJMyZ6WClCJNcberoY5ZXx+kcZhCviF/WPOoPV1/W8txe1wPAdIufIK
2S2/FLoIJFVJ3ipHfmAq2L3rbsl0bb3b4ZBdCeSOOOhPjb0NNvynY0gQVuuEfwHiQ+5ab1RMu0ma
22P/vM61+oT/bl87VE+zZOhjHSlQ/7kvP5cODLA/ooaj/Wm/bwKJRi0DAKHXK0u6w+jhcgG728Kp
vNbBYQfEpNl1V5vOjuJGqYbQS0HUrZVwCIOmIczLwi4upLzJETZCrrmEKL6xVdzX0iza3o1m1i5A
9rPeuIf8OTgFe24DUO9XjssSzp1K1JouQo2bh07XwQPM4rZAC91GY7ma6L4wLsY/0raPkNUvSqBx
kxiiT+4v3TtWV8uEr6asTcC0ZceFjuvBL2ZT8OhqwNVCvk+YsQt3b2R1p3qli2N5twScdzanjz/c
/WH1PH5E2zK72B6ymzKopQRSlwWLZ0agIXgLGIeu2DWxndHhcn3TFD87oZjxs9AWXHQ7WGIVYJ/7
N/cQqTXwLmHIAlXt0Yb1GwyPuNwbU3hTswjR6wYCG1Zda093Mb29VSAqqh7EbcOrHLPoNWBfIAZQ
B7VFnscrvEuNNDz9I78tq4tUgd5DqlUYymhc9vnZyL8Jd3lM5ePfgpgjW3ocQmZhHccQssPIWdxz
cUcLdTE0n9aOccNhqV2yAHS0A/ZzmW7InhSliyf8dwmQbdtJm5pHc0j0nrpw1k0R4PePSPIOK+c1
c1IefOChaBIBZE0knNfqwz2/Hninuvh595y+1O7szKdfc2sqL80tzdlnJg8eHTIN8TCk/P+mZN2A
0w+709lSei45B3SGbo3OeHJ2G9WOSW+m9OzlDDrBCaYCgsyYFP+HdSopC1qWHshix9+NACuSdNU/
fkI2ppeBvpi5m8CAGNAphbzbYVPLHsTsmUJ/C5PjqBOE9Qk39RScIXQv8yhS/m9bJWFvqoLX+VU/
PWmXqP4uNVYWN670Snw4vGRo0cAtnqT1Q1eO+DpLyvJp7LtA0ZeQYKeswcyIu/5E/NwvI+dPQA61
DuGX/nuPGcOLVbHFQT4PBYoGZ2xAmVbTrTyd9Xys4E1TAE51541yceQZ/C7CezG+1GdRRXnGZDvC
HJ9mXviCMzEW2J4VmtJ7Yzmf23A7lrXlMU2oScXFwObraqn1Ns5P1/9LJklqH/rROGmEGTxvGaVo
8PpKmN/u7zzlTzMSNjpE5BlGJob1GficdDZzFN+TP87g1KYjA8b30CQeXH0a2PR9EX4FkfN8knGC
vAI0qGCQHPCuFKMOCykF7W/5wOy717d1amplc4b3Hdqy7QTa4xcxNLtRNREYJG1IdKphmAXKNhHd
V5KOPlOEQExYt5V2S9xOMosMFKBk0Z4btmbhDVL3T2fzQvss05FFVB4/4SLQdlf9voy8Gu5szE3V
PJ9fkAFuc+qZF4qKrA880DiT23WcKwQocCqeNk5/wK7UmlLzXtqyucH83TK2IaKfB/L93cGP9p7j
HpbMyUo61OBBHXuIyF/OwzdrIHmBTQBbhQI2SwiRCIYIL94Glt5pKc5z790VyufFNoD8e6badRJ3
hkkQTwcfkPsbtynygnwV9mFHzObiwFHvmF0YafWwXGRIwIVyNf/mO/PQwGPDwDWzlxecWzl05yOs
VOkEu3iLGabZ53cN1nyJu6ZHBJZuQHxqyiNHtI9v3fETZZGyvxvBWl9yXLBMTma7Ws+R2aIEFrQd
unURTLkrwXhfRonpeY9wFfY62btSZum/ojmOH7ATjJ0fm6OynZDTjT5XG7YgJ1OvyO5XoTHQ/sww
wyyPTAp7o8/awdoeHMKCPzS8R6k4J1xUxL2W6cgdpozOHrcBo3UI1dQ20K/dRIF+Qelhwsm5wSf+
8g0T7fxDRSpYLAb3juADoYmkOIo37JIeYKxfUoUyaBFcPcnDxoDr83FOTuN3Ol+ZB4pWdt/eWqY3
qqRwKxVMD+Iz60AT6QW8EjvKW+Oc+HyLSbMZaVTa7oGDEoSzy14K/9GRSg+nseKTFmSyceHfHhdd
T/fsezZq2HK91S/yjwkD28/FsmFhH8MS+1amz/1xTTJwZih57ykt/RsnzlfXvzom33DfjloklC4M
5/dWUd1LDzajfrLsLkqqTFLmWJ+NL9+KybQLMt7k9+Wq9tlSa/n/0DeBikYVOlh9U7r5Nxq+srcp
6qM295tLFXBYND5XK/CSJseYX9sZS0IuTSAD3/QGcOCBInuzFrl5KCpF+pFv2V93yCDktENSnzIw
fI/aLn35KngiZJks/tQjfYZ/ajXI9nxZdY/7jFKMY/InUxA35InJyWKev/Ak7k/Q+0ychqKMjRNE
wGw+13mCQCoFB7O8TJznrxsTH3rKGNOVvTX9BdQBMWYrAdgUAFZ8y0Czt2Z+my7CO+VjoJ/PntGT
PA7/53PnGZFD+mmM/+N70Vx0lm8oB8Ik9DZar9TgnPig5fTuHhU//a3g8QCu18+jm5gO2RueixiH
nF8lY/C2gm6KvmAg/PC9wgLZ3mBsovOI+WYkzdAUTGe+45u5HUjvWCRDHErPfpIwaE29zhuQUrEj
tfegqTh39h3FRli/CAESYtppS/Y1Bs3XpXYltM5l94M/2g9+cLr0LYy6dR10KCtFLHTg51ushINm
ba7f7vZ6Aqi6SK5iEZ+eot8zfWqQyne3/+HYA+uCbvwdVDtROOPn9n5HJNj0qJpthia8dHWGWrZl
arPI0MP2cRBnSKOaAJd+6mNQ/xwB/KrVDsLLOZGTsCmg+7ZC1EPEUBJDE43do5AS8PKjmnFVj/e9
TId1mzoRZPdJFfSxGVPlri0FEM7vICAx/t5i4vBvHjD0pFw224k1JV0mQOhMpXlkotztMzzbWxIe
D6itFWR2GUM266/eHSn3dIqg3kuDqnocvanlJeX41u3pZy6oqKeVyH8GZ3slmzAGL+qu7S5smyWq
xGkHJsjait3vAZRzaCqgIHROOPCkWtjodAKHBLB/3pDKcXcBlEhuhWsHZRWIknmvDjS8FEhBWpiV
OVp45NS9uW2NbR+Tmu5bxxMG9PPZ0c1s9xx7Cw7p/OJvfJ/Z7cqPcRmURdp1V6vIPVEYnelAbipD
KI9YthtGSYTr6UItYy+gSViDRLLG/WQ/qA8HDGaI6+J4DIqw5hMHUM1V30o/Ao8nGzj0IeT8vcQV
8k/5Oe8HPx3mOYkA5J4vBqsi8FJUKeNQONYELI/A8kWknn/BgrptPMOBMejH+WeDN+Mj4KqCf3c1
fovSOXNO9mLZF+xofbitgQd+57M8M2v6d1xeE4Ac0fG34UdcUA6mxJb60+5dFl+IqiQQQBDbZe19
aDhiCjhy8RyUII0/b1Aws2mRo+xQEne1SrcMtXcAGR1q9o/g7cpYyKsWbimeJ2hxqgyJEoZXSM43
7VF+DvR8iToPZOYx51zP4bHbazg0/K2eSc9zkPDGyFfrkotuqRmohReyStXOgfmXDFhDSwIbVw/X
D4kcbkNBF8zcKiG1Kuc9pct7X5kHvLgkBEQ32aUDAh79SXE4e19LJKUf9uhQNuJc35ZJP2iGPJkC
8PU0VQE5uGUUPUYZv9YYe8a7qumyCTQwsNhvhnoJDgsBFucUUIir5WlobfOuI4lO57PjLVPcyoZa
82qwonQNZYGPzYdl+ABj3yigEwuoZjPzh29liJLkqFW6sXLtXTT1NMrx+ZpUD1Bn3H4X55EFTj46
M8WKoToGkHg85BThtd/L2IbdSc2kRSLIfRKw+puYlj59P4cxcmf7Vj1Yg5ai6U62tt6xDherDoma
ecySxNasWAkHmVbqZe3xjQZuZpVMCmMOD9z8FgD5sFBkZEdo069jgTNuH0vBJNScHIwsg38lGPWA
blM2veJbVguzybaU/nFkQeHC5odP3i58l77+dptF/LptZQdGMUxJl30/PuDYfyUHnAtGcSAmJlQw
XuNLI3a2RazzvOOpRRAmsxo8gRWZvjk5fSaB8kTrRvGOitgsEAsp7c7Jq9fF7gaxkJ/A468NSZ5H
lUheiMxU/o/upVqcnKyDkYMgf5UIeLtoEEJWv+3+eZ6RlcXPH17pm3g/eUG5GeLFZT39bs6+YiRs
kakUalIdJKdxebphErWgww8zqSUTjtd0E5k/lcP/7ZnoIhtVsfVu0srdkjguIeVvZYc57A6vLzOj
Ihy5K+cmu2/chz211oMHUOwkhRf0z0JzWQ91x8tE6wunUMYjh7QO9h4uF1t/blusA0Ei4BXCz62s
/hWuNhAaNZzEydaLcgJG1J3r1jouzQYF/dl+WYnWfleENFDdtyI2j5GJXAG+UAEC0t40s+x12Ubu
nzWomW6hwAX9WQhuJb0wvOTH34nOA2uNfU2ey79UU53HkKDN3FrAz0laiU8HzWFQLK/YfAj6T0kv
50DUuKK+YL2ngDoM2cwVTGfghpUj9GtVfGxn3Votn60J6qGZhHmHo7LwmgUFJjE6Yl6t5cVg4Zv3
K6i8pxIkCrNFrbK7LawT2S1y5d2+N2E+gnkE2lejPDswn5R9Is2VsfJ34OpQrwI96QnMj0SktJOX
Gr/DyIzWZJi5gLSP7pyZ3EwX7HEO5G4GmK4zvtf5ZqJgfgv19+pvQwlaDu3vwoxm5JQ9QRy6/OA+
nbaSKqlv8RVEEwLBZDQBMr6nFp7z9DdyJpyFWlN2x9/nvYLpqnF5x1qaDnTApEckbVOnTO06lDxq
JCBbtRKMTsD8CoezbNk4+cPRKjlG3I3IS+uWfgWvYR87Y+0QtTPXioU9VYgvT6e841HVpkdSq3mC
sUySKcaregkID1UoNE5ECgBz6clwqo18YNZt/TIEDoSgnYubSsujEVykQEe8BKkiMahqmFFAmDaj
P/VohDBEm1VDwoTl6iI1B5aqgyDdfvkEAmEw5uqP1GbTJVbRjj+orXVX4Q+rQhRWPgkcC4G8VVKf
E7KXO4TFtsr6fFn6IOfAESKCtl2XtuiaefpI4EbPST+iAxG5PI+Q1nTZdtKD/NG8DTbgxjKJPI9Q
74GjdR0ToWBavGVGTPmNTMY0FIyz0xi4S1gXNGwNLIN98COvFTWQ0/uq2DRAhhrnzOAolmrVRX3I
hLIxI4g+OLWdxhSxYQ0wPLjbZol80/z5GTd7L4+Mk0VvtVoa2qI+aQfk+h0fQAnESwh7TnNcijES
RPhkpyO10uLc3/MAo47muqM1EO7anhi7AtcWIFZUwdDfPazy3Z5wDxWWEzZQbyrJhzsBIqsXf4dZ
1a4ErlpU9edt+o7TRH+950gAH4IWPc3tQI3m0tW1uY9ZxNA7RzPrchpOWDF7jcfzbwKdRV7z0B90
7ZXV9CqhFL4332aNZs5X7rqs95aYl8Uvh3x9egyl4o82p2XXnPVpItT74+DqVZjeUTuBRpYFqO6b
8sUTul1j/gwjSxONmkYpVLDw/eFgeslUhPXCll1D8dugwev2O0RqpkmW2i6xQF3aG2+/R+h8iiyM
5IJ52BdpKxRXazPOZ9RtU1RPj1RVQo1eKZ1wBW8DpOsPcuKFY34sCcpPvC8Kc1QqXNywhH+xm7fE
Q68Vk44KMai/gzrqwWOt9V3ltp0PBKBjc8PNOrq0f5tOtTyYHWk9Z7d9jK+qM4/JM0XvXkh11g0V
f+Vs4arBKwnyvf+tiL6Fl2Q3Os563mBmSO7LxVDxQN2u9kJCzQg5i31J0AGqJ+qlGycdtqi5tBLQ
4N6gv/nJg24hSJ8zLie89fKBEI/eXC5oWBmI9cqIz/8hyuPnH4JuS8V7pdH3W7YsdHT4AoD/VAJV
yf2+E3WSCBW96J73tqfOEDCxvGU0TMkq1twKPUIOE3xaC25m+pD4kk8j71G/NpFJ0bGJXKARAmCV
Zfi7CjvCrtk1xu9/IjjwP2mMTqFxZch+aPPCb1BeX1ox4i8/Cb5QnWoFfY6gBbvYaI3SXFF5tjbD
wn0ExL2/ksVXSCtGbJbN7vwBL4F7MyQgs/1pkWCnHhwnJju7CESPrEhjfBDfti8G/8eHuikvIcaK
RePOT5tlnXXIXHYN+DvsKMKYcH45+lmLx/ZzLIKJApdr1Q5HrFSWWhjDugRH3/UFPAPt7m7I0Tuz
qwLUl2SmILfkhaDmtYrT9dtx7Ki1VLhJ9OV18XxhP/4u+twFv7LO4iFKbh+5PnO3vM9a00gkNWGE
ca4US9mCwh2gfEknvJoT2AXmM1qUWsi7HCArKZVCcoituLyR6XZbdMRSwkRMwXBTpqQyg0IaENvM
R95QgFYL4bqPq2jBpo2pzvqD003dxzZUOiZ/1PtLdSjrzyJ78hwGUMywg+CxpW/aeIH/CMk8ZR3J
UaNyUU2obDPR0zaD0p198dEwEWjblV6+8hsvV5WsaN0+ZlQRwo4qh3ikrS4NrFzchJCOe+20nXvs
5D1Pj6mpnzJMwWqwovncEN8ltIGtjP6n5r4wmnY0lKHWw0BQ3GY3/oxpPlZLMSnvFglwCft/9IwV
4GP4B+lqYrSfTT0ZEoPBt9Tm6pSZGm2UfQolKie8Bh8erCDG80GtOmvwiz+9qLhayL6dXtUSCjcd
Qst5MmPz2yrDLhsbpm/FWQK5Tqw2etDWjk4FP2RzXSnU5FSlgLfxkQH95AuvqUu0BT8AQQyt5NRB
3C/vzHm+sAs3Z1WDMpdTudAu2c0uAvvNJKPZnEDkoQ9qQborw4DrvwQ56H+e/z4Bl6tBBQxJARFz
Sebm3sIeQBjg3fKw93NM39A4rVzHu8zdAK+9TBj6tWAvfreC7VHir2kaWnzkQMJnZqYVejGzaAzY
K2HNrPy310fB5EpXQbuoFHvb5855HyxMTcnSPmhflBg0WTZHM1PChWni7mqhaM8poitLX1mFC152
QzQes46AVuclnWVzInj8GVX58YEMgJ5IEvZZ6KFTgeSOVhUeaIADHs/z7Hy6zJs53zpjdDlgYdmZ
nJozwSSbNCXiq70tkoNp1BNtSN1W65OtAttMw61FanRlRzT1Eslt9VSSh5/4DWW2hosc1OuGD0eG
zHGtEI8qtm+/Xbi7sAcA7NeNYXpGR9MlUBi7YrPSQiPZJL2O6BgntOSu6mcvkE+CMRVwtO0DOR1Q
BeyOxAWtPGONHv6mb4tYAFZoLMn+EPdm2ob7sQ+NkKhD1OpOuHIs5oGh+CbhIGC2zXfgysI0UX43
g0Z0K9qbYPO3vQvUIgB1liDtVvmSZes9Uyw4IJ6AoCTt3KZgJ+xohjNGGOxN5lZ01tCPR4GvS87Z
0VfA+ZabhXiIK2Uhxm1KlGvqxBSj8XQ7gmzXk5GMsOJCAj+HXlePXpsksbiyLMLwymoluXiuDM2+
3zTBtYtEEPTDrRoGl8+4X8UiOJeBYZgin5vs14IrVaFCLMek7qc8pTsSEp4YBYldx5tIeMKVl/wk
io4geLO1WDOHjLJ3xDmNMosnrfRFEsaUILEdRmaanN922ek49xVCUHtDGTEaX6Dg6+njwTEpO3c5
k8XT9JVlzujn4lMPP0vYmpsLDowb8PQ8R5qc9S/IfiWowz8STO/FegjCnScisEw8jPL0s4klTsia
+eK/iLYbkwsK4CGsDk1ZBXjwsbTkxG3NstMX0A9j+mtpMq2Y7CTnGSp8oItkjJWuRIoykoSeBwP2
2jwjsqOlWmeZ5y93n9fDFkNCzM6r/XdjSYIg6BcUFldsSA69jSeShK5KgkZaLq16ESgzfrW0sQi4
YYXx3KbjvxlKP7cGh2B6iWu8be4R8cU9vIvKlqUVYKzCIgrFdRBmo9ZPyf1Zu0yelEJGOYySucMR
yG3H9YNRUbOVDM5CPNvx2i32LcqZNAabvTJfrr4V/AZ2SLofffxuyguH9SImPiNWV2G/2CMQQOb5
ncX9EEJFDK92rYQhStNnU3WaRwl/aR4pU+dc/mgyG5jmP0a7ZuE2WLayURf3zqEf2bz1xLMHuc1/
+KEJ1tOrQAAtjqxs+nGds7eIFTY53+nSvyIytDvDLqdhFfhCysMhRrR4Fr9dnGr8BwZakRcP+yqQ
O+giQQk/+h1606B5Cgv8fi/mT8OqoRFJlCO25cWzAKGlKV5GoQOxvRRbn3m+P2b/8wx4GTkZ3a7H
qah5r3wQzw4gjhRO+sa/tlG0yVIoEWnvDYokG7kWOpYYINH9aO5DkgVOcB/HUodF9DfXuQXlypt8
FpzO2p8rp1kODU7YbNP/kAAl+AYU/yJ7XGUa5LHebKA/GX6A5P81idKFT3L7jTniIQ4I64VM2OL6
NFVA4Pov0wlKA5juoKiT2lyxKZblbKFXPv4+hSm67dVIdrsVbHQzFJY3agTx+pe4C5bqS3qu3mxE
1AJLVdPoaXFAbnlnQEm/YsVWJmV0DN1O6FQCbBoUgzwYaW3tKqVBNjFu91rnzewRy404KwXkeW2Z
vy9hgvEgmb+WrcBVn5jtZsIu0M6DAl4MXepnFpC2qQAU4qNko4nkawYViv8cCWcIyBfSVbVn4wP3
CoJCXfr3udw8LH5GFw6oAbCa9KnbHlEtS0L5qNsS+iyERDx+nUJGohRR4ertQEfx33i4YtB4JEd7
IelDSeIZ2zaEt6B0IyK8IZFwdCV1psfLIkjDE7et0MOxkbF8m9AfB5UR8vPoI9kVk0hs2M1VlLDl
fAaFrz+34IiL3Z+hlApMwESYeF1EYYMLasC2FaB7f+QVi9mkGOzLuPwxAa3hDi7CBU8Ce5zakO6B
LlUPpiulNi7scomRBO6zVIgz5GrMlb1SFcULAz807YJdm46q3TTh6snoX12b8mFAR9WLOT/lOTcs
OFESV8uVrk3FDMAM1B8AyjzsvSnT10vm63klv54q7GAunpT4+4uIGMmhj2BV+RcUjSJgKKoN/w65
jT/vNZF7IqOEh1Dbi4I1XxW8d+F4ZZ3Xavbabw39iQWPxybxX8RU4GOabowXqt5vJ67QYUx2DGXs
OXQlHWOdTTuDSHype8/LcwEUjhdoQyAu3V7AFVf9kJGp9xuWZN1l8AxESoRKG4dpjtS4fdkxvJYO
uJkCbGS1jcWC59ioNXFPuBax5vM5FaDF3shbN+S2b4LZympwMnJIKLBiAJv6x130a2yTuLxazmGE
KY88H54oxwhNU/Qh7wgsP5Vgn9iacOlN3B7NTmUldJOtYepKEaTT7vApzUGB4UPMNpH1wErBX/0i
JFhv5fX4nWvyqFvMaK9zqB+I6a87wn658Q82txfl9NKWI/2q+XccRAsl4AltWjE7x7xMfSMd669o
rC/AWaVYISskBmW2t1O7OxE6qvzLSUOZSgJCavf+Bb9PIuv5TmBKtcjRsfrLpMkpmbTKe+VVsUsQ
3R8WvK2xZyJw/H9OP5Ou2QEoPx5Xh6C+TmMPYMgFSbr2mmQ+Evv5iZNZoDaEEXV5rxfgE7nJmvH6
2S72T5ZWSaKx7hXxrr71IOIikcE+IF4U3wbQUvbUdDXlXK6/cL96d/nYU7P8X+1jjybCaiBnqXCX
ttmcjyS367W94jdHBoFnpJXz9Z+m+17cOPAY7FySR0lYjaVHl1m9JClXaOhjgDzpmpKlRz8loRXF
Eu4ikqxRJ9Dvu98Py2WvL7uYfntZicdRVuvMTlPJBZgQcKfGeEBdoQOqo2tYKrnn6q7K6XqhBE+/
RfN/cGU05cgYRtcl9SY3GBhHD91A6ZiIHo4/C0V8mGK4zUMJTB9pJf4GCdgLKirgFr8lfxQWLsvI
jtIR1uHSw8/Ko1JXXnK3uUh97MXUPOmEnffgdB3EqvMx3IsicL+WmQO2C3U71YlhorT0ujc2VJth
ShOjPm8ZgIJj5jc3JiuBjEK3DwFUxCClVIq1sGO6OqBc9bMXsFnNB97xGQta2HfPTZEYtG4SHqOX
WAuf+H0z+7u9dOV3k3gXdKNDH7pMY0IGaqH4A2ltcZCz9+8ub6t5fh51xuIMTuvnkl8D4YXR8lBF
c5xWXmsIiuAN+RnBwxjfEcN5N+zxtykMRHe3t0DwR+yqHjKhIa3qHCvrd+LOzASzTmL3fP1iaPT5
VlinoMBWQthMZhUXLjmjT7PXIfbPlvZO/pIsQY38wPlkY4EgqJtfsOSFnINHZ2b8eSx55TfejPrZ
qF3Bac0UKtC6kmnYv1AkKxZiOMfLoJhpm1ybdnFRI9BUdhZI6ZIZMFSqUlGoakm/lWNCOGehhxsO
TuUl3oiXacWLhRJjo0qoLDIWG703vlLCoGxrldnwIQp8122tpo/daKYfpTDrTPrgFTxZPaYVldvZ
+rKBJT1aArL3aZkkW4xpRpsFpSFjikWYnYIxLQ2kmCNslc+a1hsKkgOA/Kn3MUrTB5l65CkS441u
epmUZWsZtFp/UPNUUKR0Hh3ohksSMjN7PyTjA7Xw9pgQxwk8UeHv8bHSxUZylY3b+vsB8dvXk/PM
mrPKy6jE8a+nM2aMLTxASDY20qRfh7r1GKqEAj8igytlzmMXniS6tmM/zVhdw2B31E6ipxjKBik3
nS3ldQUlJtv1tF1aQp+Zgrm1gr3F7hGbZGQA56SlOegFOHmQSFQpmeoACxHxSCqidfgXULCwvsRo
7NQ75Yr2EVCZr+2TY2nzfqHTqTBiOmpK/RuA4z/dzAeyBp/qybWWJ2ZFbZVviVYWm9clw9iyOPl9
KoFcCmX3MO80DWj3cD6vB+uCbHBwRDPsFg8NmnHxd9UKR0UKVDw+DigDP79VxVN+9lbAy9DN63S2
MEiF+duKw1pScrcXSd8M24YVzzTXei3ZgWwacc2waGisFuakFomQTimXkGXcfErMQ5P7489kihhv
v8ho4Se771HMBWA7IaPZnyia2TyT95lALC4I+/vr0Z0EeSFRlzUrUdeP7tJPztJPNg54GsLOYoyE
KFQ7B9lpOej//gNsP+nz4A3onm4sQDxA2GPpUOu5UIiro0fwpgORZQixti5SJ075v1+tDEvgRFFt
YQzjKi+yH9V+mn8I1BDBl6NfzL9aYT0jssUT6STqNivOJgufU6bWl276J0DP6tGTyP5+adxnPvkM
rDvyriD6F/cYTFA3/1/vWSuP4IHQt5/J7mYuZoTENo+1iRFfKz4oA/aw9eOoZbRiMLvQiHJsnrRM
A2QjEhGgjnuZbi1kTv8mYkVv12I8EbSbJ5m60bGe68kbRvBFwFiAgdmT3se5EZ2qAp4sUGvNfVb/
OBPRJnV89WSa0EA4XFP7BdWibxKHYa1jF/biQIiSBrpBMGSTzAmn2qfxyIv1U3KwUQQbPj9NeRwb
lhPZaa8K6sTRh6NHHHJDAj2/WcscLxao/qy791ToZ9TrdfHJK4N+b+AlZB8NyYT2I0NDVTA08jrM
vm1Xtgtaw1J6LVDhJRZ17+9RbJEGeAo1HFLQE6eTHb8Egxmt3jcolytKy1yA23tF25FyOfjGvIyE
u/fWdfl77KB4KfN9qO44caYbpmaqgp3KoA0cAoRr1H1jpDK5rNAdO+K1QSQRBf3qBIj7T7N3YPjv
QeIy77PlrjKxFTJw4C7iDAQDcnQWJhvsJxM2wfTUmoEjee9lH3yrxHVmJ3Xpoz8Gg6DPUmtIzX8Q
p5ZdUJtspHxA4ao6RWBLJAPoQBWzs/MEcL8B7wc51Y/1gUIbbxJyy/wRkPNDo74/K2jYLP98MFPG
w0tuehDfVMLR106bCYwqfNiaQqFCkUaCXintkJPHMKv2h/faaIc/2kSiMdkiC98sRwEwAlObWviq
tSGfQsqmKpe3GTZUhVSRzLlqKMqGbBjfceBeE1RxAvJTVEeGN1QoNwLLbuE7N0IiQim3QHelC5f6
TAKO5PNPhqbFQsO5rUAD40PjQLPWxHghHO9P6DTb/cH5YZdY55cvYdMXcwMclrnW1mACeIUgE3BK
+WnHUHn7ENMilR2ei8DEV/iBX1eAB8Oep3ubgjpilAmIDcucwYzojuFcxLlBSPQb3pJkp/0yzZx8
oNuh4HLYMDYAVyAaog2F96LgCttehWqPMVuoiLNH4AbQXn4gJ0d3VAA/8PBnifdiGmnKReXZBbKV
YEkohLwg83hQkDGMF6XyjCvjce+/hFUl0jPV/s0KI5DFFVqZ/xgk5U0pxny6VhQtUsCvLZZ/uVnq
hywBD7LembDLgyjtrDQU2+kWqJlW5yNH+hD80kPvW9/iUSBGZJL/mX8Qfp82W/rehW268K2lQM7o
Z8sjfRVvCjswvEN1RrjCsBDB4esi9/9nHlooooAzRQ62twyiQz3avcRhtgh1Ea5AOwKSQ5jJtzEP
evlGXAAjf+nBn+HRp8VZZqshkXZ8oKb8Gz3zugk2cN0zLMBkkMBT8M35VSMKP8ynZRmTg4tRKguo
i30D0KWJ7hxCWiQG99X63wgp/GQGrMGDtINggWblY+lJAHNOtia2IO0I3jgh19ZbLiOo14FsLsGL
d9yhzbVrUdraSsncAmHYc+WxxbyE/pPVkwmJsHJq/0199ogFu2aBqIAl4JFGeZQIO1CTtQdC6ya3
SBquJoT7T+EBXPQqvF9oPksm5MAUXOyeXO0wWybElf7e/7yuygQXV2e63TvJ+N1IWdAfsI+R6hH1
Jtjp5qPOqM+DpdjXu64NPWhOAXKq+mqATKrgkrn2u/HlYJoTOEGhajGl1MW8gUUZpNnN9wDvXrYd
pfVVaZpW6PiU10QNdZ5D0YIE142WwypC/7Hq/BYFLN5m0+8ax1m3TK0Ihxz7YE8/28uTgSe0h58S
gaOS555nOUAgBzc+qyd8qUfnYGYX1l2Cqp5a0fcdtWB6/DrgfpMlAuqIGVr5GRo1aQnbOcOxPswK
+Wma+dA9qM81HoZ74rpvcBmKq9/j/129aHI/J2PeM35NTASGUNICaZzb+tPgYv8lVw7VarcCAZOC
goMI2hDGI/vosZuunLI5Y9YIWCZKxtT/FjY9SJPUbAoZRJRdnM7MywGBVqMjCKH00py8HwB2+9VV
IArFj1ZPZyxjL0SsqeD/XN0tWfzjdOYcnr8eZUT52wOeQzpL4Gyync+xEQdypc7jAhzQZ6LPkheg
8CSQEiUIdy2w/e4qGzlH2MWXMizkVqh1ZMX++IVe56yvSrP9aIgOK1JrsMdwSozZ5EtJfPYorpxW
GlhkG4CpzLfn0YCFZgnqgPERYE9M0geiKmMCxVt0eTFnuN9h80DdmlM3lVoUEnG4l8bSutFUgpsY
Ehho7CyB+98EckcHgfX7MG0Bf0T0vPb+GDJMquCiq+2gSTzmKSSCtWKs+GGc3EGwcWkPpZez71dW
f1UAH1vL1Yg5Xi4UG5e2K9NcgZFy77PNnMEh9bwM9e7vyrdFPfkGOwfEaUSLzoRaY66QEvc9LYu6
+CbUQIAnc740eYePSumcB29KT68leZ3LX43iF9At5XCd43XBltvPHf1UQDHs31lZFxq88vW+md/t
qfwiD8cTfwBIPgPi7x3B7DefI6zH1EZomnioxUJSTH/RkZmG5Gnc1W3eAgn6QJdwra38zUvGptrf
WfTz+qxZMKcHfdCvxmdPmzQms9IxX5pVa0wnVJ2OJhOkCNdGoHbG+UkWbpk1xejDknb5HUENrxK9
yfk/HwoVqRUY5Psm4ghRF/JHK3ALqb8LbJaHi0FXxJZIKW2/g3NCO+CRIF2MqxgkveCmU4IrjjQ9
2+UYysBbtPmfaoEr1jHce7VfCFsPGqLtnq7bwBZ5DTbarXXENvxQiLegvoT1yMGrK/Ul8UxcvzJS
NyGhyEkFx5Cz6bPCT2El98nvpS6WHRxbOapODroxb8A9j0xQWPzkPlfBr3+ylfalFLZs8nWLsbJg
9rsPMGBCESntzQaOGFVXjoFJR7+3M5qyki2KTz1dkhndtPm8eZZQhRIsour90B+Q7eFeIPPYJNxD
KJMBTz9+DvO5yHym0DRQ6+eqn6OUZ9Xq/XRxTNiKbUoreRZnE6+Jv0HR+tAudNHp62231od9XUMg
DKgkcum2DeCCDxXd5R+jx28RkgZuGN29daPAcmUfRKoKCzeiP1bJvBXAFE/YWH0mnMmDLtC/eMsj
jfyw4JH4aJPgTo38S9foVjEkVXoMgo8ZDApZmiUr9APsIqViRftuqtETvkInohBI4LMAeBIaALFX
krG6Wbe5ziQ7JX2iZKbFIDp6D561tc8f3dtr6T5YDptXDW9xQqVvvij8K8hfHy9ZBEcdQMzzFHiq
n+M8brBpm/tK1mrbmOMv6pjeUUkd6YxwSGfgiPWbegRdpu4S8MYsMQGT1H2FQ1wAKW05FMHSYDMm
YzYPkrmo8Zh1GBT+vTPjc6yZ4FKXb1zU0CuywiJpZoHrrqjEQj58l5yaXv/dBAVJn1xO7ihokJcD
fmsIs6zalzNo+BhXq47txKhoRJ0VFKkWWsaX4N10+RGqvRHO1G+c6bz7sHuDlZyN2jCxEDcCyZ4+
YGik0FXMXyW9bbrNW/xIpAY6/ufQ5IXj+1CHTbmr34DtGRjj/6ZXgt4Nq5xRqDPn8xEBmcA6L/cJ
uWt99Vumx98RSoB8RJibuWerpCPLR+k0Ppk7aB3FdGqKGLviU0hMrBFUxKb2D0fCk30fwPAbXT6c
W2Lwn1WUQ1MJfXP+34mpPi22Mdjx9bnh7gQvcJIvO5iKkSZZJ19JDvWPC+Z8Ty2sosRNwNTe5DZY
segxOqUcrAG5bTEReFZ3tiM8sRyGk5hvRS9Nnh+OHsTz9lEbbTPp7FoSQlQ3PUiD7C80y4oMbABA
87v9lIVfcl2WE9waGlveb0BE0mhwzuxiHNRK4rqIv+Tr2yS8l+FhjMOOUtKsrWMVXnL38o4feqd6
jXrEJldUnJQZuO/GX+/u8E1tr6D9HumagvpPCPLoyjL1bN96kepsVCci4DEjkgJ/62dO3M86fZpR
kB5cuUDwKDx9Y3OxY7kZuyQNByw2nMgUgxjBX9ymb2GyIEkYqKxp7wBVAaiTttviqV064kd+SkTy
rZdG9I2h77p/3UVf7wj6dyAIHIKTcFC1tA2qBL9kP7YiuGoIG4hHSFjI0TT/6EAQp2ewodoGk18x
TEQ2cjkzXdtB5sLbrBe1j26puvOxSfhqbpUSEnuV/CIcs3rFpTv0EyhMjg9BifJdqqV8l6yYnb0q
vYS/RBtah6+X6lCJJAkDpwlaCaeQg/PBO7bz3uUtAMFsL+QwcAlMdx+VFu293rqbTsVId6zAojQK
IwXino3747rk+BzEByUJOO5MMFngNUEh8H9i5i9zM0675t2FhiAISMO91TK9lPmhwPJlqqJuuOpG
5cg9MMxpyuTC7JwEBHWc6Koa/WcOsBSqEAFOCJdqZW1MM5suxpXHifDMdEoK2O40M1Pe7NyRB3kE
OkfbbyZO0nVyFkUpS/KoBTL08aNuu882F/DTdqMNz2KAX6k2Wa+HiGBB5c4Zu9/tgddmlA+XA/8r
9kbYMuqmocM4ncAeDOR5Sr6jhqXvweotHzzIsCRdCSuQLtu7fK00AKH5eEYUNlDhkZVjERTj3OiU
PF+m/wn1DLZG+JdhXRzRwlyfTbJ9DNzSXqIPPbdIuMBu939Cd5h4lIqmzZxB6lk2XH6GJh8EzuOR
tG4McDCLc0EqDHmNQNoRPzDM/dGNs2hWfBoc9wdu24I4e1ouY3AKH3kqT2teJFWxQwPWjnP5K4vZ
Fc/h3/YLncCWZHkQjyD9vzJ9i0044qQKb3YuOxNu6gk8byRAO4WXXjRuMYXESxZM4p2pZHzihMD3
6W+6aUmF/LeekVJF2jimcQ0SErhF0RQHnH6nbd9MtUvxGNW0uGBpHx+GrgjE9gKrRBtjsQS0bH2/
CXdFLyQGXfF7p1c2mB163PvfJJrCOOpaHWXb5FOCx2jbr+rkFQzKF7gUpOhz0tunKydDYR2iGj4G
vTk1XeQgU2ZJz2FjJXR2wvkjSXX1Wau9EcrmWIll9t83gcBd0HcacqG0r0c2mrMONq8fP4K+keX1
EAHc4LIHSE3oOKUX5LlbuN5+L5niIMioG7j5eaePiGzIw9yYq4glUjqgoUkvRTOatbuv21nX3ASj
5Wz6SMO81+ySWRK5WlPTJzgbHV0tpZI9lGZXlINR0/kM7KSrHp5PMKk3lD5zOVWDk3oclETZvJqb
DazknaXTd/1CviQ3V+hWGosO8XntK8mhD34+gfYUTARefIJ7SGEFvDpymRPVXjCxpqNBaQXCu5N+
bVzo+RncYsNp4jDual0VvlyEyKaP6B9H50EhJ3duzOZwB4Qdux0nM2NTsvuHlNF0VnGbg6HjVbwr
U3GydlXDl833/dC5Ezi0HLfbhe/o1nHAWkjHNwUZqCaP5odbpW7jMvj+MNqUuWxGBxGRF1rM54eT
0u+ceRWfBh4SHbhapLXvSN/yunfxd8GQLwaB2asdLP7Ddswr7/B3DA3l6FMyudgwmUPoj0FxVOAI
QESO0Z7Xgt+E5AZAAEEIoIsTGuQJ7jNKIm9CEkshNZKEgdSz+mvSFO3uBYdkyHig65lIIwvEWZ03
lURh7cdWSn11D+ym7hF380H5pXOORdRNZhgDh1W1xfx9gpaoTH3wKQC+FlNy3dZ0J8Uml5gJcbZL
yIO58OE8Lk7Q0jw+mbpfSIVQAn19ufScHlV4nKOSwx1P7FaV1wCx2H3zhBVF1vXjE/OjlTYO6sSs
kmFylD44XKixGJy6hJWRw9qrjbz9TUDQsznTNDyCQlhk5WNzrdRRy9a4AObOvrnRcLhblawjMqVK
WDPlh/Yq3n+HrZZZLx06vLLY0lvuEtav1v15NISUiHq1iy0uj/CWEGFUZVr1LnbCuc1YMPrSQ/DO
A7jfewetW+00En1fPddH8Xs0qkUOg0RWoRij+GuLUlgM6VfYu7jgGHrPKNcuKEkrn0EJ8gGjOwbU
pygq3hR56ppnD+FkX2sKGLODw3tOd86tbbB0MG6Y3L+duuC3skCtRMHkwtwXUFaiUAU9pYzxra+j
uaLUeZG0EvIEao+7s5rEjFCAUF4THea6i9GNHQhTxdzjoijlHjS1Sca7hnq6gkakX3EHi6z+/uLq
o+9QnYm9lj5s26okYNq1UGz8Kp8F0BtaL7ADIE4fogaQe4k6cFGZL3HSkNcSSuKBYYK0tF3N253N
JY0GnkGAGqAm3vbCjVcjrNd+kOIt46fI7+FtZ87sDq0EqkJWlg7Mkf7Sqtf3uxCZZyEvyejW9OSu
5UhzmBu5874COyoJ13bsQ4qdsEJwpJtnTVrn7WkbZU5zARDvWqYDnqE12Dzsn6sX3FQV60w8S5iF
11ZgrmFQl+qMNBQ/8GpkvrGPpcEeqlzvuhW4MwgIDhSzsCVjmBRaV/fYilEgVzYcAGEVGcY5k5VA
jsd14EDdJ5/L8AawB/pLEB1miCRijUCpfK315QllUnjMB4nmNOCh0GdsPWw71wElkqC5eQCvACBg
OwAXqirfQ5BwyzyBiWV6geeRDHBF7FbuiF+k4qd6BZgfjLet21LzYToCBTpLCbYZpzAGtfqDgqJY
fMwqouh/6/OPCHbW1SExBxQHvtCeyjpTxJ9eEHEaaX4/l9qvfcs8hpADrE1K/36aeMgD8zo+prQE
5T8v+6l3J2hSWSM5GB7LfLhgyNu5vMI1EsySYqND1VXqcGtIJb/b8n61+4KDpDl2cFtHZog8TMOL
N8syvGgzpCESqb1MFi8d+EAlftF9RZBvDY02me+0NP5ImqdsJB0t/NQmE4HSOeo8jxPNAPydNoIG
oSmvGraHc862/mRCDrH+kTuT9DbhkbsOPP4SP8uwPGd+3Ltgov55YXtlqlc4tMpVIw1B6ns5L7sx
78ExbvQM4teMTgr1UzNOiec65kYH3e5BoBxZqlR21AxRHJnBQ3U5hZaWU6Uamet+8I0ICH4JIu1F
jF5lD5ALKvdM16twI1svmh0vmzZ7qU/Avyd3b5L7Itz76cjs4tBEvh2colnbDuiAKy4IjXIUegWT
JYVmxML9OFZWGVyKkd5DqQKrDjvWGO0NeEyMdV/BM+D3Qo4cg5Qr6MuJ9gwkeshxHTXCwrO3+xsi
SQvRtJBrooruwEKm2kf8l6OMD5NhnY1P6bFYMZwR3Zi0txXuQ+v6wtbBNOBn9jFinE2TfJbjbmWe
KRPzwcIwEbi2OxyLLiDfvYobUwF5EOnl9P8dR3lFpvMOq/SKlrjdbUDdtf9p3MhsEyirsslqUx5I
B66ryLIBwxbriG5cEeJJC8A/OvPRSMaO60PJ9usj2srmnYlhrC3zAPw7FJeLkN8xgRpmeZyi9HKD
swjaGspZWzkQHwjIB0931LPKlEJMafBbFmJoNFuWsEdOVbqZNLXG9jqaj0+DWfHSI4K2hS/7nnM2
HRjmLYbHcwUqgD3Z6fYRRpe3S+H2AvKcZT3lJZs7gQSdoh1wa0WU2bjEJvn1UJelis1FSaiq/SGp
eEPwq9+u4tC5DYgF9U6uHtcES8NW3jIJVeJcpItjDJTwrG8bezxZ327enB1Z5m3SRXBAalOLMQPw
A4SMDHIk2ukXZ2ZLbQH+60A/i6WSAo0hT3PSYKW1HPNDQC3OIt2w1KmlfqVnz/7SClWVwf2f0bvi
6JOBfK6bsB6RYXc4Phwx5KCfuC+n/exU1wLhv73VjPKgIP3cuICN/Y2+zGo8tFMMqw00Afi6UG14
aVeE8xivSjuQ+Nu+PI5sco1DF+ECqUNl803JtyhAyOnx+66vpugrBC2om4TxXe+yd6CwtZmRzLkt
uQRNJzwE/HgIATT13CCjLPAwvSi5rdg3AmqBHoLfl6dvSH3yVXqQug0FlCUMZrT5z/RS3PWalofS
hTewCrPXena9jFv530fKu8AyqpjZQ9Sd+b4Te9FE/goWNl3evpF7UAFLe2nTO4khlgFiGhj4s4zV
K7qfGp7XaugXbcJyvY4yLaMq4obNOKTHHwmUWw9CB1QEZ18ylmlCl3J/DeFQajfnJmkE/o+xm3s1
jwkZRlEHA9uKvvtA4+oH3Dk4f97Km8CzVt9pMgSWcMCpZIaI173FOnzaaCYpX9kWj+Qtd8viGCGZ
fnElRcr5jbrtjQGAOPp/u660Vx4ONMbMV4nQZ3heMqmYX72UMvMmy56nFWnihj90UVH1rQ2KJqsW
f0eKEPltoEthxb97JYloBa2ImbMHpEthQaRebm9WdQWePf5nJafe3FZeaVLJ4FrqjuIPRg4Ht0kz
p0no9Ff8+RIus8/4kzwWTfeezfBN0ZSb52vqZv4KJoU46M2zLvp6kzQjknMKEH3uL+o3eb4zTvf2
efCybjm5ONav5jKUlnGKrx2+EIZcI0CfE80boaB1b1Kha6DwcYQXjKzazqkzeRqSkdAv9JUashPB
X0SCTmnA+MlW0hQY3EmUv5YmDDDPHMxIIpupdgU8+4EIEmGCNs10DM02CJd+syde73w+bCMpriLO
/7jkOLybsYKuE6ZTTILCuBD6BGGvZ4RAmgBQQmCz4Nz5OJgx4bwfEDShuxCVKVP3SZb7vcAA7UFj
vjTa20Gcl03DeIU2pwapmg+1XqztV9wow7Xn3i3cvyM/A23UxT+NszlSzEV+IFUFaamS2aKOkzel
g95htTlluzzI3x4NqXKCx3EQtdnSX6MG5zlNsYj2SyxkbeEqVPu+mDt+cXn5cclJ4ZcSZ82jVuCB
qFNudKRAxXc9A1zYTP2yMiclTzVh7056t2uMI2p6ZdPHCRAMgd7569W34nHdvr9ZtwpGMn97IyyX
AXIFHajSXwl/OuIkVyE5LmP15QQxOv8vWVS67oNHL0PeLCadqq80x3V/UbhtICozjsRx4h9q6uYH
DeQs9PJDdn73EgEhECegBdxee2lfjxoydUTFD9D1Ey+ycGMlo5+nIiFZ5yF8RiuNKLH2j1tXxzPL
411tzvGA1wYQFotpGUUM6EFF7L+Or5ER9Jl70z1g013D2N03l/+o6Axfz7XRqJZjTBQDJKERiYi5
Hg2Nih7mBSzrTsjeBeWcFYoPtzwtIPCOLq/YsuNJ/RsxXcgBcLRM0781PVFBjlTGg1d4PqNvMq7s
UhkGxsY6rMnOwvnCKYSCtsKG8e94to9B/VNvqVj7YZGq+ewDKcPSLsTGRDNs+RmDHh5yx0phCHpu
eVFoZMwlJ2LPqZ/4TNgkD1mHQSKQvERLNDVQJgLhsoeO4YaVgF4vr0/0ugy/Wna9FPfyZxtixcew
qoCDHfHOT4oNPJw1p72TRw5Wjzgsv1AEPWP5ckZcMmYHLoxkO/z5uPDJzxJfpPWSr1wT5rCQGX7f
gFm3mxj/sygqAFqOxG7dGvnonzRkFdoOjTLAM+toCi5uCfVDkAMAoN84hs+HT9jwE7r9fL8mYPJM
/dkyup+/F5vLPj5zrxGvaEiRy/CT/EnHl002XZIzlxEQUN4ffLG9Zv3JjLvv0lgzIkhZuaIGh7O1
BbOGbs/QDp2ULbQffX0paKkm3fxOdDHQMxWZZ1NyrhhBFCa0hHDEFytwgG1tG1mt5WC4Hpld+z+W
grKc+H9jLTwmXeXv+EAu56igO/G7XS2zO3HwYN7a6+CWfkeIzXzbGOb8hX2KnSFJxIPGXsx+jqKE
6lWtpetkSvItLMOhwlUTQJKTI5Y2hI5FsH+YAiK8CGg4Crn7xJCJg6kSYD6s+JqtJ7UxppBFMV70
8a+k5VOtTXxeOBAzMYNWvcKeMbfQu5ageDnxGlvU27bKW/q+bS/kPQOgdbuugClbNSWstmUuq/ib
hIVMA5JrxCUrHb3fYRI72TkS2SowMN59zDve3xLQ8qp6kdPsvQqPiBCtXkcmw45EiIPASWTjiYWl
CIrAb4zxal1QNAjB1P+JEDehh7yQcwEP5dKnhneU34rVhqouXFWBNtM6gXXPk8Mv9UiY+T8vQNGk
x0e/B/nrlMYo+m3Lyc5zyTKTQdfjaEZqNEgcyABWLB+o4zqMVVEffRSSS/yP/dI8Env4DGATRbRO
/i+vPseiwNaod92k7WuhpVxNflE+5tLbmpkhB2UNuFEb9/Fo+fmypLDBvOeyGgoary1KLD8qHOf/
giSz1y5VExHLATxfeTViIU6DfDsAk51YvyoHyKdKLHESVh/4btwTvf0YaTNYuObCCny/oqGfZVe3
yLFRI+QX1wcCvvk/u/PFf/HX7ECeWperx51B5M/8C5D/XDXYpgbnyz47FRMHwEKnuFj7+/pXu8sB
so5RCRfGOXXqjPwnq/QXOChjRmOc05SmqAlNksc6glN/IU+ynx37xAhWZOpeRCeLWJ/AhZAMovZX
AZgCwZTuo1NjvudUH6PABw0YMGDMbTlrtD9ZAfOgoBXzpmwL58W2DweKABoDS54jKQgFnl2JC9Oa
qmZ8qHZK/+aJOKpHb2A7Pb1p/yJoMcmoBOtJS/hOyJU07/hAXbJYyBtuSKqYTo2KZqsyYc1ol3I/
kxJaKWTApANB1CkWmS5WWtsSvwnq8nlIDmKnoYa5duL3mJzju4jq5m0hpKM+0o24+/AkQA0L5jdx
53R3JbbjmRChIQOZHL/mNvL522CfFiablLkpLAX7IhSWijBAZkfQFhRv1lkijuw2xVXq25pRyGck
wUTWNUs2gsN1e9rOVxE64cZwXtDZQjguMHpwgxRzj0IJljwhDzEZumtg5KjtZRE8jAaXMcCf4ms8
P43pMaazB+kGuKO1pc+sGoRus4ZvCTZmBAIdI/lEmLwZQIL+hr3IQ9JdjRmWbvaMfTnUN2QNjKWk
7rBluF6zXuY+ZjCXMlLl9DYDPgwJgJRL1DUpxD2gZr80oXmgHEYJ6XygCZo+UPGX8RKKE1xxxml3
Iz7f5fdNN8aKr4JQm1SlBvgzxQC0aHtKDTUP/W+c9N/C/wjFmZ3cY4NQtahmXTL2gWGGD5ia2Lb9
uoIemIlveUMFWl01qnxXdR8stEqX8/DYZSNzbRZWQmYNdYm6h7TVyyeemrNiU7WkqcW1BUCfida2
+dLtN7ISLTptWqtmpuJlCSFuVZ2fXLyTWXMDWIK7ikMqpjTM917FCEEhjPzCdBQkIFX9LtPANyyt
+tgIQl1FXfWWZ9zbeOwZsQDCZI8Z0bBtd8dvStrxLncS7Ast2Ll+2vXl1bt2/dPbOE47zFXE71hJ
2FXZV2tcHEub5C3hGM5l/D5u1hESLCqkv3dsHTAjk5t/oRzKNGURcMZiJWceYqDctuGRLDJ2FpOp
Gf9d2gIKCwc2Km48Lsbyjyh/+It7WQr+LFYSTkn/+FvIcAOzj4berKnoWkcWcVlME29EVSZB9+4Q
jnDcllEz/21Z2O8742yCw1/UsTtK9ppf+K6zDgRPbqZRHXTSHf5BqftYb/K2S/qTLpiluLGi6Aul
1w2UX4/ke/U0kUuvXIaOHKfc7NTLFne5Fjk+6G5rA1/Bp41TRGqlUnDeoSXm1/B/z1SCJfO6j+Um
agW2fi/Vi+rX02Z/v4GZX7l2CYV/v6cRE0ubzeewaXd8KhbK9cRSVkB1NqXRETwB68KEKvLfno7n
4qnDJySFgCT9cY2B689pWbr/OZSiqChWF5ZfIEQ5WUsxqpVOKUUCc45pDRgUECSRzic/qoubH1vw
Fp5aH//aYqHMDuy4kzt42tDCmitP7GL1sNmOjDpYYO5YcAL0rEtQRz0Mqf42zVjEZxPGT4xRR8xD
cxs9XoNkc9erHfIT1GnBGSkjNSJd9PIlVwh/xN8I025EmpBdeKFzlVcW5j1tZCjU7NOdZuihOlpf
KTRCzmmmD2W01vJNBMTVX2zA3TSw1BSA72HL7HejV+JN6BnupjBP29hkqHztxoX8prwNRj92hgRc
KMXIcNEB3NWRa7ZEHm4Ky8mjbvf5BmRo6uMXA7w9t7kVXmu8OGXaGjt3u6Uta12+inkAA6j8b6TL
4S19P4aT1u1ZBSozHAXhj5az08UjhDgMQch9u5FBIkSWosMgI0sDPLcZFRZcLeB/mdwSyYKAMD53
HPwgBjxpxlEWyZaIWo4fZQ0IEr15jGhRtwn/pSub6jyoEdArjpLMul+k41X/YekxrYDML83fiZP1
C8p/5IUGExsWj03OoFkBzLjadvb63FGf0yzL3obqy8cTCXYlbf3+A3oiVM0+pzKQZeooG7ryttc2
3HGIEsUmJnkiouLIdGpMyaDn2qCvUsx3RvwTdn8/mZEjssgUjZ2qKBWNdFDF1l7mErt2UEDE5HCu
vzx879vtBvrhtVVE0KY9XZgPNPqaOvkN7wP2FtBAvYNWuZvb+UpgIxul+/4sD7aL1SOzBdD5M+lK
76iNY1b1n/+gPQvpqg1GKuJG5nU8N3Nv+cb8zu6dOIeqicyTruOJEX9yKDadpHF2+VYCEEPOt/3F
jOb1xrohDCVwjflxr2e/LpjeThMneL13qHUcrt21R+H6ibKmrfGmwiA8fqNUf1fykbfTAnrZ9Q7v
P1JY8vCFIxVZj564mts5CDi0CmneKloCcwQqEdjtTRi5Wvbx9fdkvdK+4TnVjCRl1FPdEZdy1oG2
iaj01pSS9K7f4grSx10eJeO/5B3FPbMlPoWqDlqOT7KaBxxRNv9sYCZT6Vg4uW18A8Qu7Mitc/ub
VOn8zwaV95WoQAuUeU90fcbHFx4iakAEiYf6kZ2IiO/J4UW8HpBUoaOOAmDiTj7xgdTmbz0R9Zqm
LgALlJRPDHZDIMMHohv67FzEd0y3vfCPz1QkZY//y93+CDdNJZU9inWpPMLjhbdY9+wlz7as3ac2
ZiiEIyiU6ZuIiqiQQsJmKVY6a5RbEsAWpvkQffSBrJ/xamqZHarFWTzGTDJY8wqTLgV43JilQHqc
X3XhV3Ae1fZrpt7Z9liUz6KOI4EsQ7LtbcwjrarlXHfyajAaFXlycuT3Ffu3YLtWzV7FAWQ7pYIe
8Soi3joGjxpR37ZqweuVOoa4bqdSUivuL5qmDwITkGPUkjEGVi08JywcfD83pnrRuyXEz3EFHibD
AWyx/Dq64gxdv+kNwblcVi7MW2WmcYZbBXFpnhICaQxrUjw3zd4Wbdx1TQ8h7WJX/uZySxxHAKy+
HEvZtr7B8Kse9+UBDjfsnKfjN+MSpQRcG2dl+eqttfhAUheP/ykunqED7Sr/RhkZMKDBMVEdnumn
sS7A24/45LPCuL5cI+R4hD2MwSzGIHLWjSOXhZ7sbauMspF6XKNrQZDRers4j7i4kTNUolEsRI/k
y1Pz+J4oBI6d6X/wA/7b/js1egCDSYyxGrTPsFrGg0Nu6tLu+jqloFPgjQUAce9jmI3tOFVMVaWO
gTA2GRqe6VzeMlXagGTkZeWMEEZqOjI7Y4xBQ+vaJ9l/UktlCUFWtxkX87VgoWdozQtgbCUucwGc
5A3I2g59Fbvm8xSh0G1iGqfchDqyvb4FSC+qCeUZFLMpwqOr8CIlWHillg3eC6Ajg0eGJnXErG/b
daRy9gOa7oXDxlAa9do01LaYDVPQYPa/IxjWw39zbALpDO5knba6wcYZNzMYvHpTJim8McrsRUnp
Zf/IlW3cPnCg0/c/n8Tl7hpKjS7iEEP7D+1BpYWj4x3hmQpnlVzmbmMMm+33EaYw1mVhbLYiNA4X
/UiokNF74ML/o/SJtH4O78lF1wB7jyzm5gKG42qufPwOG1zLsFKJduqr7q8ZUNYBtAIfkchKyQpv
BnIaGIFXVLe5LZPKZHExLoKTKNxSjIo65eGGcYPmdu/FM6yB9RgG2ZrrRbm8agSl8/grHQM+WRPo
F1PBVmpDxB+VpoydEDUFG00U/yfIsp9LaBbA/6lFj+EvPNFFrOkgGlqhBhmRJo5ARlyvr1Hdm+Gc
UsVwJNwltXmP7WUe4oXxM0HrCLf31lUQVM2s5Pzer4Z3M5552QG1BKHMIwv9TK3C+fAEMe9QiDiW
49Dz8QgqtL8HWk+CTJOG8UVkjPU5BqywQvUiTA54FJXy/7Una1nzalaoRAa0GAYbrEe6as7n7HKD
meRktS7TiaTbw/PpLXlD51SYUGRvH3M2Rw0NlCnJrPquAte7pnY+GtcblAL04ac9tj8sZ6bSvnVv
tEy6W5tmc2kwPa1D4DtnSr5nZ2c98jqZ9YzUIKrMXz4LedKgNbFVic9E7kMxomjefm/xM5YTbA2d
Y4nV9GFKvE18TJzU+i0yDRFxtROFERL7wWYoPtG4FbpFnYyjaoZpAD2rsmXPJyn16Kqftz/4m1Yi
p107HXmZgz01UuxjssK0SFqjTKpl+c9+tcu3SXxCAgSbxDiHSDPlLdv4EYrChGrsNtHCUO772tK0
U5d4IW7yhuSncqFlzF0XM//Zaq2J2ed+0Mnm/ZD/OsR3YZlsbPiC6Q4uSpsbBx/oIggvQGRUL/1x
RguBoXQdAVo4V4TwRNxpGda7zyW3d9qBax3Fm27a3pi9dCyOZ++3n5//Ya4r/Y8Kx3Q4I9BK83+c
1EOpTR9XsFqcijV7+lcYQmntv4gL66WYvDbG9AryQzagXi0FpGXrOReXmkOPBW7TQKffeKWN4+/k
qvAsTAawEliTrIgcUm949nRh4SLDUxVbWUQ+Jh5aOluzcUJ/IF+hNx57JkCS2krrw5cfG6KDd+Q4
0EiCWiWCwGOCWSfbKsDpUqcr2CtAdZ9mE6rRhpEyrQwnLWtJDfPJWHQ6gq5cA1NiXELOOFdpw5vv
MOg9WZA5O1bUABU3wkH8ZfOXmWhhPaTd0dfVFdJ+WTjrnMBm2+JLznNukmr8L0CZJgXQjE2ioasP
0UL52Tvo3Kaf1zeMt2IjcVV8+GRkCPLg1HiWjn6cgIsllQqqvIatafP8sCpFPO4j1LzvWm4MzdIf
KQUHOD9QWjQlssM82yp4OfnIEff+E5jclCZkp7TLVpStBwK7rzp+/fYS/wYX7OQ4z3XahHXboQc8
CC2HZwkfcR9l19yPCvhaHbdQBAJfL4yciq/8z4Kt2Es4sZPvzvDajoJP9Ac7ll03vYksxiU5oYfS
0n9+7Ifjcjr/7xqAxKMdz8EcWc33q8ESR+wfgDs2GCyAbFbBgu8lCA5Z0WOhqRqDzMUKFWmXBNLJ
lzNjqso8QAF56dab8B8f49c8vsi7dsBuK0Yz7w4rsyWfn+h4C050ndH10NNnHKt/MqIKsYJC0RmI
tSEjht0/mwYi65/ucRwx+88aX7fFJMeNvuwsgbvl0+ttWU8KxETzSxo5BuehTFHzpbvB23GpWvIJ
7JLLaBKaEcaODWvTnL5qgZW8gUHmw89ItgR0cAPRnDCFm25/Lb0pieYslnbp7IBUMNHzWD/PZxlb
SRkv0SbwXSGs6xk97vL+BqEWeS2WXGIRAjN//x/Ds2YokJnZtY63DoNgQgKrEpyKdhCR+ywFhuES
86IsNqXBawHsJgqVRsuSMfq/4s4xlh4sAGeFUkU7D3fj99QHQA4V8pm2cV6HBajlVWQuR8VTCKqM
exdxUb5Yih+IGbVzkfsCd8f+mDSgTke6Ghus0ONo1EdBWRCruRYjYdpOQppe4iyuDLOW6faL+3zQ
l/RowNOU31X0IMNl3FXqKFH1RA8vPIQljCfvW1//BCvCu6AAdZeKKxzZK4FxdHNH9YWGmgNo7vCl
cA6m/iLec2y/9caeOdGl3gw+KjoflJWloCr/2t64450rdyOSNPwayC+GM8h4wQYIfL5OCTL/NTXl
wHbUGoVA8JELmS7BnEnIVf+bjXeQlnQCuImyR9gc1hoiL89bgZFcQOUC9dmGLLVZNvFnC3wNYSUB
04N3GTKqhJVy8H8qgxg88YG7KBYS2aKgO/mpocXTP42o0mJmVKGPJcLTWqTcGGJm0Cr9+4tqG8GL
YcI8bbaIzuodEIZ+ffXGF9ju5HKYg0Fd15I17bqZbQm8X0IW+azoHQw4DKWSQFDv7uMgIcZmboi3
SSjELRwQENmmaxtZbs5hlAz0rEkFU8p/tRJMGymuM5O6P1ReiehUUQX1m0mLNsa8/Bh8+Vao9OA0
wRd2W7QjwZJ7OIJ8XhtjEuzw6cB11SGZdyYwyE9WuGnYgULAvf+jdPAh/4tbl8eUv2h8qXPSXWci
EDeVXKp1wYSruIThzVf+AfX8Ck6Qnj0UJYVMX2eBzbFtz+UI+8heHB044ae/YkAYjpT8d5BuGumW
eG+6S5azgmLRVUNDm0HHsT1f0OXxNfydHDqvUr6xgBwdaWhaJvvXe6nv64iuZRcM8uywNinG0tWL
AcNkd6qTSB4Zs08zrFs1lgi7ijWQEt2IMDpdSHXmAWWw8WbkTduzGEA12MltP+rwCUlVQ2MxKt7x
quFh9C9qIcaEF7D2l1YbqZOtZ7m97DOVFVj4DEJBQ+9ZGw8jxqrXXvlYyEGxb6fFjS2y+co3HoIU
hO0z6OR4lHOzs7XhLKZhzYTvhT/5dpP/VaLqahPlto8W0qKLQcsnEVM8FF8P4guObm4bd2HjsF+t
ohKuftEefQ8V6N1/YqKsvr7FgEQjkwAubK6PuOzVBX5LgCGUHLWIoqAMnNmTgYTp+ju3MNT39AFI
89GtHZnO7q6BvQtCRjf5rWP+uvC/rFuyRNzfL2gURphbg1yLStSq5Nb9+oVRGP0XewAx7C0h5WdX
fB46irRpZf41umSvcwDI51/L1jYJeN+I0bWQ2rWbFOXT7vjVcsP2sdzGnyv0SWMi897rnfdGaBuH
5Q2AJ9Y875DcEG51nQk/3OodXSDyjXn0v5ZGQly8WIEMqxvKVLWevuif9cMKzh6iZ0+DkKlL8Il8
TgmVM8MnitfywBfZU7h/ApWJ2nyLrpsfOTKokkF7w1HZI44kdeHKTY9cfcyLLXTszfaQlKklZkE6
CFOXEIGAU2zNCKLD7HYu9Da8o5u+GowPfAZSuNuu0ExNSVG2ydWrcZb08iW2b6psuvoa3Kek9Mpj
EnHnk7Fv8ZIV5WeOMPlcOzRaqcM0MNVmGX4vWbqLfZalkNtLfKjA/d1ZYBKnH5vXV3hHusH5mwlA
KZy9WArK+FGr3N4s35B+WBs0kLe/AKV3J5p8wMdv2nrW4PrtvRTcmRnFonRDqgY11oQVycnb4cqj
G3Q/FoGwUYOkaOeyDUHwhpk0JXSln893Kj/FXZf96pRA+M34byZUt0mzdks0smpJQQ/q0QgzHO+2
vUhWMOOvGInVVrZsjS448ykjk3Tj5xQ428KdaB8Iz5ViQQ0X627vodYxaVjvmz+OF/UkYnLcZCtZ
gP/EH2DVPs3vigWn9aGxORhuj2YbOi42mQgtcx0Q7p3kv/RCeayR5cQZ0z+G+bt6YDJHEySdcnOc
uJhDV9KGQcUlpHqoLsU3sb7dCcaadVMwt4C0Fb5Pj8+1/mv3yIrYucySRt5X5t5Tq4XolwMkg278
4zHkMBP/zjgsdbWhgz/2E+bPIurc98n9kfMd/f7zhBZonP/6BTVuvxeVUivZetbyotytoJNVwjBE
y8cLIoT5bpq2LXzTOMezwObZw2EVOs2uW26LFaclmHb4O1ITQ6swphJoCCZb/AtPTyLd6yg7D0Bv
WnwPEVcHlK8cARFLJWJwwrBQG0p99G92ZJHo48wJxX48Q8E4/IpD2VLlXfyTBR5dm8N5tgp2ya+J
rPHbl2K/qAnrkJzplE0OU1oLhsd3zXeWIyXcSage8iTN1yc2zakVfsGpWeDDlk/JHniFHvQFnY/0
QZwhrYWZuP1fEhwEReld1uaVfaEVW+ujYP6eJadTWXzWv2AnCTWP7dbzr8K30kaFrmYtgbojQuqf
Js96559xGyu8cH6QcpXOkquFInCbxmv9maaUK16dSGLD2tL0vxCIObAx/aI7yBwxJ/Jmz1/nXP5o
+n1xnDsXeAW8fXxDB9O2nsEboIcj8hUfFHQFEk5pHWGR9hcHrj7B38HbvbqRiAiYG8sXmtdBHQ/I
SSzdEE8dTmrnQQLS1OEG2ap16y775QTsuYLvt8MzCA8k/+HIVlqh74xewYlCVaEyKuUW3IxfHfsL
BYpzBh2ag82bG6urYOPMSve3aNTxgwqFHy/kppPWbPf907qfys6Bem3bWqxL2EVFFsG26FJUqleK
7ynLWm8l8VKU9ZjE0mMI6xrzH17ey13cqvfYoh0l7T2Yb3G5K45nXWfVh9YhuWqdVeM46LusnTn9
YK9W9SrQMlIRmq7+YgvQ3nfjHzfhSBGLpLuO4Lnve7b/M8GlZFcGSIbM9CzAnRN2N35dbHnMcgl6
1kJpoQB1D+BzmbxHUNdE70PvHJCA12dYtenW0zWMfMJT5MAD3aDbvkUZFKHAhb5K0xUw9HocvWgG
XQ4Hl4/5eJ1orJZM5QYZOSeMxzCQnieJi8rxGvatbplX43PZSmkPT1MA4iD6z449b2rUvDOSjI/r
CpnE7szQfWy8v+bZTdU8gRfHBAw2gEze98OkdbeJHA8GD0Oq2zOLovycA2r/DS5/+eyA5vUZKhzS
sZVvLNM27MmI2oXeXmrAEMjESIlKfX1doyyBRjVCDzs3ZHYeMMQ7Mt/FpQHfG7D/Vvl9wySWwszK
VM2Nkrb7zSBDmYc4+eP17Qe30pd1y3iv2SqE+6SnhwEj/p/ylRGISucAKEB8YSBB3KFSIdSJB9F+
wyOa/jo3fzEjCntW40/VcB4/il2dbbZEYuzpF54z9beh2Z0ulyUuUbv3Rc7KUpF33hbd16LiPn2f
Po1dbn6aDB6UOieUmZUms5DnM7wdUjZzzCcGtTj950GDc/gix8L0D5/tk0hp+yQxmA4iY5cY40jY
7I7I6btdERT1yM08WctlJtECmFpQUums2gLEAQfskcLkozJi1uf+GrCBDn3CWEr7imh1dXAGorKr
XTRXx9Bf2pUb5A9vhAiHNbA1ul0GPrdo+a+/WH6Z+o/MOlVrwYzpmG/b6yO1MGXiNeiMiX/jQxbN
AR7Rza+ZxeoKrMgaD9waVRNHyyUS78p0o8/+sItucWl933nmaJx5PZ2sBH/N5eWOk+y7hDx8zJ9K
r1Wdx0nGvE0+rkzjja3pwRKYK5PgyjKCM0DrlieJO+Y/fzstQM76IHi09ng5latdopj6csysBBZZ
4/8YIZUHBRg8mFxSzGP5WvOPrG0veKAyWBnyJN5HE9grgCJaWN6vYgTFoahfb2UQ49cwoi28QZdt
5OOq5sDh0TNzD9mMeJjENIXZmD6/yiCRcusQJWHUDVw0iUmkCMFGSX0RvTbTu85lmPnKCs0Wh0YO
bCU0lbg6b6iv9QodsnLXivFGoHNIjLKgxagjlvcnTW+BU3anQx9KJ9g8WZVYfmPzhqHWPXdzXrP1
FCaEiToeYydButP0ADDg3A18uOze2KXa08qvFA33MYEk+wiARGE4uhqr8lgUNLOPZvMaghpGbYTk
VKMdyH/OEIejkR+ZPcSzormpnhJTB5gnEw7b9lLN8ZGwLINPFF03f9J617LhlLvBnQVRXg6PNjHp
ltwPfoBFjpPI1E6iSPe21SMMYp57L4WBegTs8wVnt10Z8lt+8tu+NM8+PcA+55v7g3KD/pe5x5OE
0+foWGzRgGQeel235nPGQY1Bbx4yNpwbOjRaumF3ICl5SGzo7V1YBnJsoE4TZuNSEKnBYjDm7qUS
4MImqzXs4UApECYdVB0Ww+RnZcGNooEH1Dm4PUjvXcSegP8vRf6xjm8PRoxPLmpKcGmK76cE7qRe
pL/yDfpF9SdklDQlwhsJIGh7csRiZGjbwDiAhfhg+Wc/8F1J2YpgRAhe84+8etGwMHsHLjBcIXZY
vwAVMZzDK6Phfnskh4HBOaLdPsANeAevfioaXTkTjFCjtYCIgSKhXOKWrVmWKI3zqNdnR3aOfPyu
n3tBHBu5BYqiC/k38GwVfmIIjh5oDzEwsKV4sSHqoAVKOiYZkZ1bP2k3yr/JfhsUUGphIXpLbBxd
5Z5U8WC+/hzLGcLy8cHk9mrnGOfosJ85kbrVbYPzTmVJB8DfWWocukI29RitOqT9ezp0ufo7J+XK
ngWHswgAv1po4QEqBitUx8j9GRiyEsK6JUX+ZHoYbAjKmtgJXH0L56HcaUAAdHzusN4RxO8OJh6I
7BMjq2HL1SkERBTvdjKo+ICx2ZnuvE9m/fdFoyyLB6DhNmSGtfuxBGAzcAgOSPoSbLjM/tvBrSOT
N215/D0yqiofeYKYxvghv6eI+/kv9z1a4idpUoHhtHwYBbEKaKdekPjqiWghoZFxAAQX9ezNJ6Nt
K4ryKqNi8Lq5HnJoWz9/nA3icDRCn4HD0vo5ussD5Nx9ZHadot0vql8NJWa9ebG3Sd+JwzmUDAsE
PU6qcCFGQsJzY8g8/DprG3bkoIqe5YhQWsbR8wkbXxo3bD8sL+Li69ls1FvP3jxdwY/6abKCZpzb
hSOlFBwlAWvxYeXguBsX4b77b+Mw9upF19/FIBc2EnG03i1VSVdOlsE5dV/NC5/KY2iNedvtc+Co
NR7jti/rs5jyCNdRVuamLCPyZnWdMwr+BuAzQRup+xAK3uJoHBs2/UyEbOvlkmWXxrOX4Ch0icSg
oThW419jvlyu4sTr5yuOtpCR1rYJlNkVsTj6cI7Cl79BLU0hW5q4OSnt/TkqBekzfOa94PlG0ZuS
fD+OvWs0cCgkmxxh0VnDht2BmpveKXsbaAftWj7N5lVQP7yE46Yxmkoec5nny0KZ/hRqJDApM8LB
/RlUcVHMALQRi0nll325BgLuqohlnOgyHSIb/XEEQbQUVj/WTfgY9nlsxpJPtp3gcnhr5a2fBfbP
TiVpHCW9Oo4lfRRHzHEBPU46J9d/KQR2vM1V8IkTFQP4XOUj42BMLVmxwv91WwQU0q2kJY4xHs4f
c8VOnXS0DBpKx80sm52Tj78bhuq1FJbTuFD4b0TTVSpBWi3iiyFTQn2RVXvbLJeoVudbiUpfh+8J
UJIHZnXgY8jVYbDuoXdip9OAct9yZATl2vgYIzFgeA89C/5St1dQ0uazZ8GleVm04Wf0VyD4Cb4M
tXz4aDrpnmRD9bmJFwF/51loshitld82LE9lGdVq0H+w5QIpLpV34+TY14VlXC5lKZZPE02IAaz2
GGw4bGyFvhPnfXY6NHGI0uNdqkanHXXLj2XGOnEGLKF6DwHaTTRBPUKsERoDUsZlB8++D4U7UL9T
MQr+HEyJCd8UrUgdEqmr/LNrNYqKtJUwQHXcfRaXXbTFBSSznrNFUjuqU/bNaoXXV49xqsTSjZLp
1b5DAAjO7DNRe2IXhBP+WaVVOJ/gyhbHXPypu1V+8NHNxs/N+pAVBmmikEvmF4zvN5pGyKBSTKf0
EGnikgy8cx+9Ket+EAkieGt9RhH8Da0pIWu5Q1f5QL1AiUFBatQAaPztbTxvq9v9vXQ5MGwcwyxC
lWFVekHPeN3kzkBEy+frw9bKLx6yRWXe0h6RfOL4ukwbGxlPbo3NNwcjiVsIZuy53yFnqD3gqH6h
hP1fIbDxEASJkwWj7CJnQEtv2mpvplLkUxskSRvlTTdrPHqM61M+SMWIwl9Hf/5U7UXtl8VwkyaR
acEwrOzj746NgbzjI1GlU1efR1DD39ZVfPhwo5TMykMq0I53H//GIrA8UwWUVjAM3rdjJq1WDWu1
xBWzhLVRwBGtRyMH0u44oHkzCtUt92eEHt6NOzlsKw9dkGK9maRdPdQclO84I6pCMmbr5jZIPyin
o2ph/cYQutm1WzRbztfblmFUUXlK2uqxUakzM46u8MG2jFVQPbvfwyZ82ZSLi/zZ3Cu0pZYT1U8v
KpYYIx//TOIB34X47Xm44e4V4sW8/SpmHopBj9gtZFWrUE3qNT20xRx+8HJpDsP6F3lg1C8h4WW9
Nt+XrfKeHP6ZaZAoRe3Rr4pV2nFUG4Eirp4nxPszlK+s35Dz/ViIE2eIzWQkrp7bptijJqCjTC5Z
AAqMIBT5amqp7Jg30vyimFQPD73HJBvGWp6fpur35Wl18IMOaCBkJRD//H1ns7tFMRf+8iZ8QnRO
aP20cdkZH64dB8EaEXQw0DkvJYbNRqaFQTbbgXisveK5hg5jBh4PIIzBKX5m1v0qXWYP2feo3muS
L3o2jbUE39Fek/qOhcD5fKWrU1apDbArT4JJDpWkECZz25XvoklSGRi0atgflJ2aXQfBdOndDOP9
OV+w7L1eBwGmQPsjYO9eSukqv4MFdIE9jN9wU9nIu+cim7mIjZnxxecM6qHVzjcSF9PR7470XOtU
56Pc57e759i/7mwRcF2HEjw/5n7efaJR1IGP0Gh2T378/nnHbizWF4Ke13GSQAdFPaCeFUACBzhc
IFwR/ADvGYjjPmXvygMqelCnONlsCfzODtXOiwY6YQ5TUfdDYU9a2LN+7bIeXGvW+cqFvj0D5YCi
xl0W4PbRSO3ndUOrgVel9+OgC4ZuHh5bjyT7F2sQSzLr94XuZqcvJGrmB8wojRb7sEuUpToypTZg
EPCsppfoD/PkXZL0YZvgd89DoHfRYj8EfHx/UBZUa1cGoZhzbU7kqHFfFpzCKnkIxjJyNf0Ct+NW
AIcpA4GIPphBvDOqEAipf96ZTzfmrgdp+mXp7sdrbBRRJ18XrgfAH21NmDZxR0zAjxe663kEX23X
YCRmh4pzbcUz5JIjmhfzM5XJeQdQxNQ5hBqz7IjJyNFNPSMCuNviBTFylK/bpdClp9TpbBxsslba
KAxXb/Lw+bJTUlwFBqYJtMZtYe+6vvxmJvxMVzl44Ddqxh8W2AS/gagGjXdhx8m+8bHEbLA1PkAe
ykUSbhYrILqlUrZMgVN30G9i9M783aLGC8aYNLE4E4ArUyMY+j3QKDeYkbSgs2mDpQ0jxugaKPyE
yKpxh9z+SRJSSvQF+lL5PhHqLspeXKkUA62F4cGX2TyztMuaBg4wmyb8hoGjnr77ckmyiDDjLqe4
NSnKJ9d1iCxJkZ8j4Ussh+GCKJK8oP8k2/hGivN5A1Y6rWEjrtJbpzGrU1+UdyD43ngQmbFdY6PE
Oi2p34/0Kl7ScLJUcW/uZ8OEVFZKP8lfQBbQp+7OtX/3K10Ze5j8wRGZPoFyQuS6AFLutFn2iyv4
BfVGkTLU+KihRkREFnfQrHUmLorZaFjDyC7yzpFpdF4+8amAbgDbRO2VVWl8xbd8FzL+1fEEvxWL
aSdidT5PpYLqNxQJ1FoSJjrhjvuxnhxstUDoDY/3vRMgql39ZVfLnEPJy1Je0NaBeJtwzmXNPtzF
S+cplUM5/HbQaBnzRCY5k/Z9IeSzBlWU4OF9helem+tlt2V1/QynLGNebp2JOa1B+dJC3wWcA3h/
68DoX95cNoDDZFh09q9auzWzli7IEYYpdhX1Lt5xwpvpUjyGqr9+4L1IkIPdUQmEu7TpgNFQtp4X
u2ydmhLyLyrxumeP0S8bK3QQxcejoHQxMNcw2BWLgRPYUGaqHzUmULM2ivh94vVAH0S8kCdSaDs3
+YYKAaexTEqi7IjoB63yUcu2vpbq2DJoMKQpOZr8i5YBBZRKPulwmLoXi8hVaSWkge/5I3K8lZOr
umLQVhRCrr++IghxNQJ8N5GoVD4U4CKwY5xx8TFL2WKqRTPgAVyY582348ASmN27SQj/kQZrWK0a
kQCouBQU2T6vZ55WORk8jKAdMKi0/gjqDVKXIASFZ1TtScEXg2jAYVuaaIxTHM/07xvHM0rDa0eI
DDAzftyPugURt887QLP2pD7dgb9x8g5ZOzx/JctnvowG9j87iF3LkeOgaQjaWmB4pyaq1Htp/oB4
PWExkLRu5pupe1QBeUgFMHCIrCbj3a+7vyuDAZH8E8EcXdyRdRdqJr3YmxzXaqEO2lPYo/FfzB0c
j9Ue4FHJyw5GVd92F0VgP/b58/r6ZdADyFgU5Dbh48wELibpnYEcN5SRcA6r4GuELrMSHuExRoKM
9f5eouUdzmwUnyP7QtCj1v/X9BotwEz9G4UYezwZg84hOQlkUPTC1AKBA/3bifZ2waEXAQDMznTw
mrTY0oTFFPlsAGTsPgHB9TTAuMO8VMaP7SHBP7yl6lMhMHpaBbXf2XAtOMV/jssJ0s40tDx2gwTf
sPbccXrzZ4bLUaXXoi2V+HYfC4TomRlsyRfhrVZ8OtC71ggkpYGUNn+icAUrI61KMwpqlQ3JsXuw
22pk5R8Z+mny973YbyFSy9wZN6zlETraFQOyPCozEHa1ZTuqQSzjAV3RGTgfl4YKrBDoiE7Uqwn2
srocc4jnqro7/g/7ddSfS1MMUL47Eb5ZGcnCOgK69EJUycZoHMUTy7scF1r5fCWGH2ktMrNjWIDA
0nFmG472krPicvDv4YshMLj9vmX3XiCNnN6Xv28hFall8peT+7TXT4SohWmlpq+7o/x7SWFK1hRZ
tTb0KacCMi69Wu5fCBO2PVN7hDJemSb0MxKjK4NrOTXZn4w8B4BA1+Qy+sp3bDLiU/2LxQJwHS/j
QdUqobTbDajt4zmiA0aluFJa8H3/g/O5Y30T+stVuNOzuok/lSIerNOoqKX7y7Pp3Bvxue89IYU8
Ppj6Ywd3xN93emRv/6lE7toumB8u05/ibwzL4EAyUGJOMbnxjL5Ws8qGDiCH3U41LQC2n7ac+g0K
rgae9O/CsK33S0YeIUp7WCum6zaW6WjHzV6J31jdveuFqBLkZWdKAGfp6bTb5swGrIUiWpA5sAyy
W+UkGvAi6fzJrRlm2HU7cd3jsqpeTlKOER6CH+aW++6QSlCy9A4mvlShIqpGyLBijQAekpAzHjNj
boVMeBU7NkBla8UIvRVlVMyd2zfzLZoA4qJ1FA6E8ovKSb196KrsfMFVLNZHZTA6hfWqMe/29Lvj
RLr0tbYQ73eOVmk2FlBUiUNlsvgrMb+h/SCc6Y8zt9DAOeTkwdPdbToUhA+vQq3hkQtGV7aG8S/1
mTub1r+s3QRwu1EZF86kvxm2cAfoEj1gR3EQRa4XlVS8YXE7M1VfvQqqZ6mjg0HbHARX7oxECYn9
hu6avAsSO88S0MRbE+NHZlQ5+TpI8DJ2We4rpZJZKqzrG09wZ5GXcwBHjioCf2zif/ApSiS8Nt0H
9ww4aIsXo6k3RO4DDVGcQsowO3faHhezCy7Pm2orzko6KZ3LG1BSgagINYt27dvb5KWQUHXzavKj
rULgALherVkg96KzDsNez+aT/YrUwtbGMQwclNhYXH7Ts8qTXwDdleWRw1HnPOxIi2YrxUplfs3c
xNK1M6zOZb7lP625fbTGE0sxExBd+DdYxp6Bv70Pifk7X8Ju4WjB4cu1qvDB6TDEA2bS+0GNfZ4I
+8/X0lFNPc1U9fzsdmTZxhPg2V3YwM/hjcEbaHS+oEFi/KLWoKqT92WGKdSsa9/gaX9y4KHuYkxl
LXRd8y6H/5xS/8gt51Y75KTUoZMaivhQgQGBqsKZhrwbbJAGwGd2izGIB/uhpBtsA2y6IQOBfLOW
ounddfBm7iPHXhmRFBbJvu+E5RtxRsavs8kLrezvwL1hfVfMuyv4AQqbe2AuaD3zL3tcvvq+9Wun
XHCNB/4ggeW+ZyqevCZlXbrN3wap+yaQroDNGVZ/dQ+EuwJnLn9IAApREc05DkD9Dxw72gC0zDL5
eZkIlu92+U38QCKnZrtwJMrgSBy9+UxlE1Pl5Rp9reiKmgI4g/Qltm0HtGRtFISTbktfbpmXmpNu
w33+YZwEtAVlkDtmHGAA2IPHP5dOWO3mBIbUgVvzk2oNDJEM+AcqmCwZelm+BFgcai9noxRE+yF9
gZMrgG7XqdpdUpe/t7EyxWWmNu6gjIX6cN7+zBu732gqT0yH1BEyuBywohPiR+Le+gyvBjJa4EH4
qCyVY8gCf0incRLR4B9MrJP8vSd010xVAWXmb0zlsgZw6ITU0Xf5PJkh6WwjqF/aOR9NZg5Wy0tb
ZIwSfo+kvuQy2qYBesfIIZagYiskyPJNiTjR7ch4PGJJ+Nloxajt9OtxtUJ6J05Xf2ct7GX6zLiq
ypAvbcDOMgjwtb6Z9mZAKEYgOo1Rwq+i4Llf8P7xCoo9yIUtqTIi2zCpnsJP5ffGQvbF1wpHEsyt
rxc5a0XTLxBg2pygmszVVa8xCA11hSOVPJcvcZOucPC3Nll4YHw9VfR3jzuF0eePhgmmU7LeH1YA
dqr8CRyQDJjsrLsyNsCsIRd9V9JRNJQQc1XFf4SOpBBWY61Y9pxH0ryUUsCTVKllNlFi5wDOo3pw
DUOv5rBLZM9+Fhs5j5vSms+XXv9OkQKVSr4M+74DTn1Act8ZZwR74Xu2zYu8FXBI5T4SsEwq5wbe
nHzDiSy57w6SUGMEq239x16XsyNIvBmBI8/2dgoa16V1vP6XEDaqRvS0hSEsYH1IQYWw+4n6/JlH
A2Nz6MTFfWur99w6fx8m6WNQ5czq/UJQWaQaxJsJGh4ybDmZnXEDQgpTXDlGQKFMZoDBi3YpTtWA
SpWJigknkt5aliP0gBgtxpbamZIQBxrjLax+XgFgo/M5vEYq5ZrAxCLTS4bN3C+kC/d643Y215QH
AaNuKuK79MrZ4Bn6X4FSoiFIy0/vHZ0ac5UBFQlPAW9055Oxh13ZBu7mnYVULZwnDGgvYZe+ga9n
REEoaIp+yumIecaiNLcNdkj/DIGoTtx0NCL0nYfSB8jKPcrlCUKUk0VxTfiPIFs8dKN5oIwT5VD8
9zm8WL5T5mGdJ1UIWjXWBN0VtDzj47tCYoRHEVi/OPRVuNiVnodZbkgjwQMttHVzIFmXPCmLyAKg
PUlWUeMzhwWxeqMZ0YKPf7zrY6oeAqS0yS2TFHhX8sq9xpYjohIR+/suLazTxljHMPVtdiLbv/W+
9IZLatF4a1NRuoG5bLMhL61Q8p6TBQouxLWtM3jpNbgbZc0B4uLo71mCBSRand6UhiD21v7tjlWr
PSjnoCbuJBujU7gkrPIC77Jr0MYEm8C211T5D2vGlHaSA+U/k3GkH8Y6aG7LjTiqvDfhq9QLA4Js
rrH9w18L7kvInt04O5BuG3PjYH+TbAbyqXeEGRiQ/BYYiPCnB7NyNM6C2HhsTeFyGn1JpGuG1qEw
FEHRvLCMyR/JmxgrQxh5bQ2JjD/wlRCuFOV8R1IbkQaZHQY88CZvKxEIDarXnX98mVBn5W49pHfh
427pQlGoGGTkYlXQUhJrkRU5GCyWYebYrKd6wuWrOhyW8S9QuTMgVvqFiUyhrmoGR2FoFrOPs58S
Wf2VTlKLb9CkjqagT4wih70X7kmkVF8CsX6kiBw7AsHh2emGKRkxzpNdu5qSH/gcE/cv0R7mRnDF
NNEqg3qhxj82xAeOuN8vpBBQpQJVhg8vLKRF9pXaEMYGFLrW2J6a7XGuV0Wj5qUzRROPxr637SBD
R+hWYNO3NeBoB+4FqzfxVmpl+jHnRIvYu6mvG+s9kx1gKx7U7nqYXT2FRvqPm2o3Muq0Sn+lJbA4
jGh6FwQBuVMt+xMAI7PRYYvgzKB1Cfocdj0G/KcJtV6NFc04yJ8GSEs0/SJRnjm+R5qZT4KmvO7u
Sl02xUcxhbXBCirYhuJpguuRjHdpxisgtdCShTCs8uDszDWPasled0vlh1BdD3S/CN72Ku6NzPo8
lZuVB3h61ikE4og5QOy2AXa7X7LRW5eNyE8dT2ipSfPyK0jpMeOps/uvwEFp/vBOIY/qQ4M/5nXC
WZZcre/wkU5FfQo1/50L7ooty0tpEZMFCXxaLEoMVWRRFNqt6ll5yAlh9vji2Yf5XvEs9WIQfVjG
+Nki0x2rk6BBxBVLLgn9KLo1Gu81mXnYvWYt7D+3UZnGdNpS86L7dGxCdND5EBeLY0AyEPWNUchq
Qw/A5wH0dWsF6iajNzHtHmfN6b6zFI8EgH3IuzEyJrS34Ql3bIv6qIA3yIwlfDY26/92PT7dhnTc
tD7ewzEQv5EcE8VAJIyBjfkNyAlRPFrbijlvu8H8rYPKLtAwRjd9LtOfs0Nw1MdcEwipjRDbnCA8
bBAtLR2TLhHCAu9y6h5ULqoYSpedy3TCuID+Xymh2w37QIHRtDwbw+Ao35xueGPaMEgWJzVOb8vB
z7NS9oV5G6xPrB8PeFWcdYTCZyMdQ6c3UbynuwFI3BNtrZ3Rrfw6ZZNkk7N8l8W7xFSo3b/W0YxX
HYka+xVgpNAgO8QG99TL33G4PQ6kaEs90U0YQ5Hv4sngv06yH0PdOFrNShHBeTdUYuZJIAMfeDVO
12SBFS+4gjhfquhKyp0yIMuNZCPFZUkyu+jXxgQ3W5nMXkvvAZTEYGyUzA8qKMjwMNGhXRWUbucv
TLDNYrv+y0lzNrh1MF63x2Z1rw5Ou5MHK/H9/6Gb3MIboL+E3cFGNsM++JGqpuC8L2gaIqMQqs0Y
ndMsVKGbdh2gGgM22kzXHCoEZx7jo7ZW4z8xLXfdtjGkzaQVOXPfCcrgfR/KFgF2CZQjE97knlyk
h/FmyubNymBrYiREu9u8ULdTFL40JE76CX8IKs5iPn+93ZeNyqIUPcpido7LIUQ97zDM0ZKFTEMK
Q1Jg9t6oBX3vWjnjrlY61u+23jXTptcvUKyg7/62DakV3gPzKbKHdccprM9JICfzlFIZ4/pQD6MH
MDotGyrGUkj1fbpNYEmJpDEs2QVopSEJAR20m6vGpE46FU/rvJO9PeF1Jw+wvSjSttQZ8fk/tTIB
keslCmLuCZK0hwfEoEnRtNUWehpW4C5wUMOiI5EVs8fnpRQ68HEAUOORfEnngFwuvt+B09nVviP/
FdyLvdiRXgH30DrGVho3JGkZ+8VsDzp+VddG/4bUKdAWiXWBlo5zPMwT5MF9sJfeQFjjWRZedjY4
KjVUF2gJ2meQ/iSybQ4NUQnbdy0aKKNrr7FvOmHOv4vk6GeFep6sdMXMMnUkiIUf3/hlOENOzMFw
LJMJ0a9FDAz2PA6OEq/TS4aEjnryu1YhmZhQ7RYpLAdrrY4R3D8UUS+7OpoSpmTlBGtDm8DEpcZ8
JQDDn5V7BlIzXWH1x/hTKRJruO/bk8dYnB5xgzitOWO69SR9Cvtx4r19tHwEk2omGavV8kp7qwS1
MD0stiHUCumQ2HfYZzNcwsH0XwMeVnfmiPCP3Nn6nyx2qgWynh1a0HuI1VRcwc+TJfl0bLnXKgPv
2jQ69dLUzVCyaxTeywDhGHLJ4dg2QvFj24E3qSjKmnnK6CPoIzl7ku1pdUdyF2uav5BuE63koR11
gg86o1H4CuTvSwwWi1H60LKAGAN/MmWQgIXB2et3a7V/Gh3rW9yspTaGTlykvCPrbA4ndjsLlqos
cFbo4WLoLETrTNAQHAaS3HT/vafcJyjpQnWhXpSkkoHb+F2PdUWAX7fD1rCw5N49RQZvUSgUqFAc
klS5J+JDBS9MENk/iWio8yMdiHigS1FdDevfEP7unkVFN056C5y/AD2yzY5BgqfFfk09qzFvGpOV
8GyxNPl18Ucfee/L39/FkzZV33qvMpcaK85uw2iqSyfiHg5zwfQXTzNeZ+L+dfJZBoAQ76XTrLGL
iz8X5SL6HlzFl9zbbzeatVmU58tgFqTDKm5sJC9PwCnqMkoIS+0vhgh1d3rmVgZZIoNv8Y+ThrUg
VdJVIarWma7kDT0bS/ybMMudR7IRWjVjlri48OCX+J2PZiSbY9itl+ZrkAgdx/Z/t6KJRZqcXung
5zEf8t7SJ+DYhlrdu5MQm8EALsfg3711RPjVnF7dzgbMlZbRyqHiQEdoKFP/JoiLb5DidiXB4jsG
v6cjsUhRWbk3qXW7CywUf0/Pl+bE6nPKIS/WXHw6j/1glO/TPC+xxpPCxFqJ1uVSr3227wLh+aRI
cKcXuxUMyT31VpYYn3TW7+vtmdLaWkl1TIpBRUmbFaccVaEfwRTJB4m0TDuL/5qu/fpXt8haf1Rc
UL/dGvYUgYBTcBM15xFVgnUSqnbRbVtg1EHKdODYGwuyVI/bMH9BrUYrtbesw05s15MrqKPh3Nhc
9Jv1bnwelOcgIi711BeqBF0Q4a+Q4zQAfJuHTpN8rQETfnynxgRo+C0tawzvE/1c7tMCO/ms2sA2
XBAv6M75HriPrWwzq8684OdTBQFw65C3jJql54gwwrBFkEL9VlcKF506qOVYhbl20BIH8zfyCORZ
5UgM/uQ91MJQeC0Yiu9TV6MyyeSK9m59/YYsPaiRr6DMLRjt+ZG+/7bIGqCrWINFCzgPGZ8eDSvb
IgLE/fhJLW06qnKsNPVrsFbEL5r3x5Ejsv7wNcMmSx1q3ayG3Kvx1BwKKcFhG0w44OJkSsPTSB0y
3amV16OmW+my4aX52LIVFI6d+lCbMkfoYhAg6JLwQrYA2mx11EUfiAxPZU2rGaHCq+CqgMH0DY14
Jt7EqSalpQIXOCbRzHbF1QfjisBpvwHazI7rVefGryAGr3ktEZmxjRfPjkKBheaFE+7DhWdT9YwT
F+tbzA3Sjpr75zWwFw3p0He0JhRKWVU+fmzv3I1pFeIivwllysFfiizMk5VN12SRkJcoIl5Ri5c+
L3SoLYvfSAmU9KmtbhTgZWtoIGT/REoVWNDEU4Xj6NgkSKPdItZ5LYuaJWBQuphBgGL77dvf3Ggs
Nk8VjY5kQVHG27x9sTV8mwW3yJdSqW0t1sGdJPOGzzUwjO53JR9PYZMXNxHDfd6Ge/l9DJ3/PB0M
RqujfZtjBCV9KTgkIc0iGXRhdobCKMLwubUczR9wxqYum20zKCkmOo/A0lnlLrQW82W9TrNJ94qQ
owuiq3+ka/eFGBzEuBMDwC7gAzl8Z6PysbYXOYX3R/z8pdv7jy4RZHTLedfB+5a33G1lk2Oowyrv
A4Re2RH1MfJTIis1h58dzrqmPK1maGUkJCTyOZl4uCsrB0OlMHmXEb5WtCmWFA0hs5oakKGXgpHp
zabgzKfbbvxI5ROr0D9wXIEt3dhzInPn/1ilWojapWASHPHRCuyfHIV6krA4JC3aWXaSp01rTg3A
rYzzeXFeZCKcnNfhhTqbwG61Whjvn9TE8aATM1sD5yKk2gxHf+D9z5RtVw00AgHXALpszExPNKMh
RrQ2mK0XApnNxP1ZJv9+chGAq5ajCVp/cgOFix72QgMyjHu4Gvz8TlXzU1i967I0RSa5w1DiWDXV
Z+rTrxORn9GCLtxhvfSJlfyDlTwxbxYqE8nY+wvQIUujVeVCKV00RWbkQGOvw6A7zlb+9eEBwqRN
LZmta/qLCCnGknDvd7Ez3+NPVJWEPCyU41mgmV4iDsq2quk/YYkVL5Nd9qOgkUzB5F2dYZCWVU6u
Etd8s/ltT3Pgk76p8wzeYjEtXG+K+knoR7NDDaq9LvTNob6f3NP5wSBflhkaopgl4HpiJQSebSrC
QwNdyydlouW6OMgUX1g4trz+eYDd8V7s+W0Y3de95/gJKiyYL/sefdVBiuD4yGzhLR54c7tnDeoD
VJcFAU2RKoswMsa/0TLQJDkmJ0MPWDT0fmF1T8bcFgRvQvLFOoFNltCTILDPLL17KZdU9eYG5f0k
kmen+bAEkFk0eYQOue+0l+XqQuwN8+z9LWNznpUoqIHjBzljMZNskrIz8LqWjbVGbE5CSR2503Ir
SvPHpJfXWtEIyRE1P4y4NSp/h9UFQzmiYkA6UQ1S59XUxjtFhmLWpt52VVEYGOemoug9dW7sHV8v
4I5CT1XZGtz5OFnL0wxq6AfX+NHXYRZ4ML1jncX9PaLHtSJwWUgBxqUgysSNEgebWLoXfnaSOLLR
xNJ9a0y4U+l9MFstrrSmMf6u7P1zrvgBm9e/h1Nl46qG2raQJGPl6HEAQeL4Me16B2pc8V5Ttnwr
JhRfnMVfDXa8zav8rurzCTsK6zCnhBWTfMGgzD50FA3p/EJNUYYyJ6AHqJ381WQ4V/CdRmzpyw7Z
tSvP0ys8CCpcVKpOEGEpr6wf11Kbk6DYT/fCjwIVj6jt5vdJGrbPiyTMHF4Cv9wEQd6pL6/Dbxm9
sEZz16A5HpTNoMBklpQuS9T5CQ1QPL05CUjrkE6bmQ2S/5WUEo96fILCtcoHOd0iT/ZVitUuNids
BQy1i6h4jU7iZBc6WCy8p9L8iN/FPU+SJHaW9ZiygePzyO7r7IvGTlHHkygxOvZ8xdvu6yHKZdyC
Qov/hkHq+efyI0iatKgnWBbL9LtCf1bqu8T0nX5AciavL4t+Tvchwl1X3Bzv3b4kQ7FAvT8ZQBat
karadM0+8a+xv2WSIbZtqIQ5r53M01E/Uv8nef98t2OnaxVUGaq/2flL8KVXGI3OvtiKcZsp4Zjw
sjW0Vu/g69tPWOUxf9+6JIBR8HZaqi4nOzUOcUEoKvtWW9kGQ4/XfX6PIJdrTA4zkVVHE8YUsqKY
hOC1NvtY+AJXPwtz9z/jly34U+h+jItyWAPWGy2gqd6zoB3oS/B6nkdgbz6AhO+Ap4A3C1OC6mq+
VsO4Ywoc4/clnvSi4eWokyGRsaHK7mssY1afXiYncD9TLRdepXafOc5pomIAptQFvWRTSWfKjcWd
rPCmKxb7BlK4owKanIxpZ70UAEoIqq/x+a7sRpUvogrCiWkZ1rI0n2kBV5q+lM0FOZmqU10EJkUb
15wSSP7rx8NIxE/axS8QUlbB+kz0wwl2+mYE0+06WhzQWYHtKq0Iz6xqfZOs3UYO2iHI9xUC1dTY
sTOUbBbrRt81goIDem3yRy0bLhNCyLtKNzru/C8OEHSchmfryHl28ca7+YQsTXzAroWKNgBe34SN
JUvbMB1GrA7ET4UaDGT/s5WMGqJCRAEGe94XASvaFOtEVENl19DPlWERXv084PbCF7lq8hjwawTi
sBzW1LRLc5fWHXXhkn2UGJDgaQM21tD0KZJl1CqKTPxnDZ9xHbQqO8sBXDcGE3uQOihErVxUbahC
sXGttbwBGmDmU0IozhyTF4nZ1hsvKqt/xAhwoP0NA9+PiIe0rR40nXHSyOR7Vi90BPeerhUH4Tqo
vLUEFLdHDJEQ7S8lflsPIjoX9zIqItaKevj40E0SmIgqF9Czx5D1OBZAlW5SiAH20VwUC8v/bOkP
Wv6g+6YR2kOmloxYHZP9IbnFdZu2CUAnl5aKWe+Hc0UdOcq4TP4mOcEl9Cr69JORINdvVOCMaW62
JDyTzviSh6cVKl3KMQiZ3rFGU4Z3Fcza72tAmtrcIXLAqOuijbS9O2V7Vxt8umzJ/vM9bOa+3wWi
dO6gFu3XXmBrI4Pt/7KUfOOIAyPSCZZOx4bjwIFuBmcIzuWpTUgKIU/TtWVCG+kQewFyJs9mmCfL
8CgyiiFItnBT0oCHXlQqDuarWY/G/ZnvlKvZ1tgHsSlV+W5Tubwiixw6yiCGRAB7ztlkC4zYRBJs
tY5fk4T10ZDhCNrFa0MM+xKBNO6XYWRtl4nh4BwgIwmIvKj0MOZibB/v4CbK0tOEDyg/HqnmJEtW
rDSeoTuZgIIazS3kxKGje9KDIlEoBvoecHw1wX85FlPTr3Dd9yjgA8Jg5ey6i/7SsAL+Y0J0K2f0
YH1kJUkHSuiH/JplAd/c9DKeZBKjdjNgtJf9/5UC/GQkn64rERMC0LXzOiK4/xmHamK/tDSPo+jW
HAivKZOAIgPNrQcE7X4XYKES6OCs2tX01+CJ1l97LQTpi4hblZMUOzY3jNJiuV4zSQT9nmTMzZ1c
5VZ++/IDFeaJdv9Ofoo1ygJ8vEh6iGoOeIxGWfzPoIyahPpXr6kXe64guXchUMlqQO6pft48d97B
kHh6pepxqOC2O6ZvLAR8AeXyI7frIhBTV40vmrZ/AowwKIm29JKG65DVt+AJgyS3eBJzFF38Hgo8
zL9sJy0HKmVHAPvqKwm1ZWxBGBL/FTBUR4zlE8DMAl+3Si3a5RwiEtkI1hVqiit0ctiyL+9LM+FO
Ncv0B+hZkn96DJf9jwwTQ7pJZ9svdmeNGTZHF2s2v6yhAENwobTG4YPXe7/I4LTSMQpTCDXYQCEH
ud4A+bPsBvma0D+7Xrnal0a6WXISO7/N0IBzjDbY6YqCoeTNd6azB5c9zRyd+mFTlMVqDNFp+T9J
2cvfh9LWQQEJRa/aGIKfZP31g8b7JHRAYbURPjXHFot5Jk8EDgpLQ96x2J6ZyGDisst5/QLSB9Qf
N4r7KTM9oPk6UlV+8W/7d48/5Mvp8SeoKIkAYJ3jI5S4xseRDayTx90zZPMl1eExJ85wRrHlpE99
HASGQULXesUqJ/x8Bb0Fk/mtsGrkFemQeg8+EHzP/9beHrmrgOGDNQdDEKvMMf2cdpwNgZHVusdv
+0SYZ0H5Cwomfp2rbFrgOCNPfTSDx9lISxbHlphlg/zhYmcFCJGa8MG384gtj8913qmtSJvu+cFa
WPa9/BtGJ7VNLs23ATQNfqad7BAaiQu03TxmfMo1BHA8y434sz0W7YQOLendmZ/SnEmztYnZVVL8
ZVOqi7y0zJ6M24xAEE6TCV489Vy/fsNlNJ+enTYJ+KlcIQbtS7w9cO/8YoDaUhELoho0fTKDLDF0
oiX8MOVoHnom/n04k/SM/4SmMdx774efZuDj69/3dmKtyWHNwIQCBentC+8PG++ftU4o/d7iCc3i
Me88iF8yBnNJWRADAx4AJiufgkcDvG0PZCdhcfTQ8AQ2tlWyJaP5feCVBRaoJgCwED08LadQlyua
FmpuI8053q3Qyu/NfFu0kD4NoaHnZ5V1BRioposr9zT/t+myU7QaYiFzcBCn82B1su6GO9ba4K1a
DJSQ5RvuiimAir3QfFtzT0bCBS4wiFKY9w4bN3XZ1sl+BGdjvdlmoB1z3ldPhuXaTnqUshNOB2lh
nF/zgEeiVySjlGUz/8RecSf+uXhdrJcxQylcC8knga/uSJMdN6YcNPDqHTkVTZkRkA2wZA29KJ38
82jr9fW6Q97F1FPzVh9DFHg/Vmw4ozhrnQQE3ke3ntL+1e/4gIAK+jWePCfaqo5sYKBhKnmWbjYS
whnHni8V7LRk2JSCeJx1Mz7OC88FZX3uEheFCd+Lnp+7CcqvnL3Etwfot7IfRM3aDU9OgqkjiKoH
kUmKg0LWDCez4rfPQLv5L4mumBbkXoXwm+EGIFGX4piGAASmgbkyhhZqqMmSboHsdwh21QwOPeIB
hCNGHrJLhjaKTgCKNN1C60nIJu9C+G+AWhlFd97MS/HTa+jeNdINqN3mweORuH9k9SsC9jkXkzi1
cboD4D2dR6xspi6r1zhuRjvdD+kJ8Wb/VjQxZ12dk6AsCqJM/oXKNw7NEBLZEMKDVt2n7hTct4T6
QOWMicdl+qTFRZBd559lanKJw7rekhh8HrEVHUr+c+rKKOx6i6UlQbfNC/vYgy1xeVUpm98i+NpY
UnXJGMZ3WTTIE/vSTR6rxI0Ho7Ef0g3DtblcD5HuvNjIlPeOh6onRRYUGE0ADosQnKBVfCxV3gAp
4PjL/3t8J5tUPxoQbIzpS6lUvE3ktv/X6dqFEVDPppskhUxqF2EuugmovSiB0KxbxNrJOwc1oTY8
LE2B811M7L7Mp88A6hQS18vOlTVNpvQ/fJTn6NiANti9QicVDelJphHpwZ/+LQs2b7O3KEVaGjC4
jrPO6v+1nRUqFd22VAXDxTk3jtpOHLdST2sLDCUiVBIlzA8s4sdRPKoDw2sNgFSIP0YT4kUUZA3t
mhvLmbovcQ/SnHSovSfLcTSBJYFj2K7fllM/hgKwc9Jjz/vmVi+29y6SIeaV+9TUFD3sWumueDkk
uXjmYUX/oLSxmxlAq/69+y2MMBQ+bAhCvShCplTqMvHUI0u6leOhjaceAZkOn9Q9YSq9C+u3m6d1
1IqXZGbLiGprIhlPXe7nnb0s5H4TM2UHgXqTqwgL0dRGcxntCIyzK19xTnDJeBIUG5/9NWKKJXKX
7uHe2havYR70dxoRT/wnRP5MShRqIA3bUGY01S8cbq1hsDszOpd+qLrJMW20dvqtwSWWPeqGFgDC
BgghrFGc2v0n66SGmTug33wN6qtiw/Ox2VR5S9NussPR5cnu1baZfxkRnpPv1bpcTdyEEZIfjKDb
MNEzOlxJHXTzLgYEdgwPomawAIwhGQHGgHNOpyA66t7Z5uRHJ73Fx7WjF4xeTk+VkzwyTK6hk2h/
bMtLGsngaZK3EOPep91LnYSYlRxjut6ZqBlNX95OySt4OEKGaxvdd3KuR2PHwHZgeQXYFp6TB/iL
HEYFpUPJJMuVM13CLOD1HRuGMrc0yFTDv8BbSSzMPJbNn22dixlbJaLjVl1z7QqXV5IPA4skYe0x
hJTt214gnxzhYQGdBR+EKvlylM7uKJthgoh43o9q6HZ8OCgdFXPzsRFbh77ruTl5T9ykIWnYBYmE
gecTenDGVjS8C4CgeefLjDUhh5kkZ+hq3bxfIhEE6DLCpfS8Y8ReOJ7kVWLSLbIOZSEaYSqoKStG
d5KPExPeB1RlSUSdmi9SywksBx1Dn5M1pMbaKAH1b3mGJ/SrRYdPCgKPNXXEmbxChT3i1wB+8Cmy
xJCiPi/P+IH3HCMhGQ38oKtQEHNdWVcSrCoBCdZI0mwqKfe3x2Y5m2wYUVZkRZmTegHCnX9NknGT
UJ08tgL0qwgjkcEC3K+toXdWqaI5PR39HD/xmu9us6ubYq0quYvDp596ZY90p1KegTgbmW0m0lYA
1dyd45nlXYeIVQSIdKb4SL4vz+zn0j14AHRvL7d78WUFoMu5JUybF1roOdgtvCB+cpVLHa3ljuT8
w7XbmJEGk1UekJGyX0F/Lq6mfHkZvRvRYkXKCt6YrdKhSw5GIkWIOuWWwgD9kYcfE1i2GV5crVIK
V/Pek+q+/IbG67tjoa3zq9c8oIpIftigq9uYerGVDdV+w/+BQ51KgYgY+Q8efs1v3iEIRdNxp9gB
8z8cZpY2P9Wk5ZKpRGiairqANH0OZULX4RCiCLgade9Kv2lgH4BR53Ogv+oDcvFr4NhGQdNCE8z+
5ErATHd+T01XfO33Mu77Nj9s861zFQk45WnIMo9Sq7yLm5h46EjFqazsVGYr/+BaMaT3E5GF/4TT
UX4jGyHTP5V1mQP7k0XSyX9GOJC9RYrdIcIfoLRzdSYo8gB+sdxZUVqz6FZm176oB4yqPV1dnO4x
4YffgLLeBWL/d/ceiRSPDtmxrTd8wBuesb0FGwOUlegzrkBfdy45EyFLPZzsDNsMk2012sQr+Pes
TqhHBoaJhgByE+5KTy+q8q+vZAiVqSj5BGfVUfB17DsmjiNQFl3E7KKV2P1Lx5IMUVufl3JVwZWK
GzHW3U+EJ/BAtkYz/UFunMNLnuVjj5xI+qbhxTgK8/ZxdEhWVrxZXzPZJIJl1dADvfpQXIgbsOu3
mGK4tRZsq/1pZG10UzLEAf6cn0V1PyAUnYzyy6SP4zz6d+2L4QtFLi+wecEVHchPrEQINc5wxnaf
2/jUU52pw7AiClzNIpvIt+kR7ms1BuCMoKD6TMcMrB9G1V1TaxbVa8f4UENAiCppDjOZthfv11Zc
t/xSZVAnapWOgy5HmzE5iNRu6EifqojU1ZR9dna1ZIc25o0A9fxASYTX+zuBu5QUvQaIG6ctqW6G
Woz3v+EXMNETTA6ASr8RkSjt3u8se+XTe85AhepPktrGC6kB7zWzJOTA6j1NbKsjDIGy9v/hQBBk
V5hJ/mZsP3Kt2ba8+x99tDDYzTysvAAtLxYRy9/m/7dQOm0MnDb8RMHyPwRlT/rs3GlSy2jlUS3o
rYtPtgeBROg0UwMLb06dL6IyKlfRktijcAr4VY8hNbacgqpJpsLIalstu+gcDEo4fgrUCUyGh6VG
rB4JQXSrqXxOXX3d/AQvcOo0GLpPT6UbTerHIC08Iwlcvv44zu5zDlgjTM2bDzLxVdjQkg++xJ0K
ipl8NgevnTgGJ/7rz92BqLw+pF8GL6DQRoXhIE4vdFH1T7PtgjnoiPNv/WjPXVUA+JpBaxRiR80z
RC4GWT3dNqrBVJMpbndCT9mUld18KZ+ukkr9KjVhDOdHo12QP6HQTQ053ws2sP/cl/MfZVDGgUqE
9hAUMVZfPwfhNp+zD1ckixg3kYh4wWuaUDpi8by+lL8FZorkDlne0NxZcxBNiX9N7K1J+4w6MD53
kADs/Jaufj0FsjNartUMaUE0U3njIxGo9UEBCDOTFHvkm1+J0vL0n+WYdo/InnxexwOqhB2xsZqY
t2f0o9sIkBaz+4IpazJ85bW4BGy6SDr9q2WLnK+By3aSaKgGwI7EIrcTJqM0c0SJgBd4NMOGjCEL
5SkuOJLjVtnzMHK3+HH6n9naxbo5jsjDQH4jBvBO4c1hT2LedDJIrM9Af1xATzGkV4ySDZBy6rh7
1TnHSazQjGX3pI0ybiI4WIeGtHGfxZ92lt9waCgtC50fdwsS9wwmehllkE/TJPcVJsafDJoehyX9
un+aJj0BV3ovQkVCVt9wfqG2M1i2UP4/hqHzLOljGcY+sr9Hg2CRGtcPK91cOWOrQsXSIL7OQ2KM
evknU3P/7xzn/vlv75d2RuYuyoiktBUFUzx5TSKG0toXeFmgRg1QGMZyJ2cA+/VQh8qr42DLCJQd
HENz+rtgU8G9eBAwPBCp+pg1P0GrejQs9AtZh31RBSh8y1OKwIiyzVwxLisEbe0f7OT+zB8uC6PQ
paGSFIa24i0NX4wB2Zlf+/iRt+rVtKTBH2Dq81Yfe+3eoQ1zjsWM8gBAfcX59hYyfO1MKmjzjg+Y
XLUZYVgfoC7zjxW6Nbbzw9oXpN2dulZorOalYpz/ll4AdK/WT5wc7bQ9QUgn2VT33Nr0jCH/l2wZ
WgBJUfuWMFn0KsmIh1Oru9/JKslzz3XD53RyH3oQkQpWHLVD+HrXQUGaSsG3XeNA9//Q7D1kOKtT
eIDAZeJTqghCY7++07Dqti1Uq6v+nqiFlEfk4Eu+qrK8craKG+yWHOxUpwTlkhhPZc5CyBIADre3
hmmUtv7AZPGFm8Pkn9wgX17I5+EZFDB/54GpCppur0+v6utz+/7MYYGg3wqWef/vxhpyjY9AHNg/
f9Dt36qZPhbG7R0utaiBDuYLHph+mIq53IhSAe2B2ChV4UZfW6jUDJFhNqAcYyzY81E/8JUVoRYW
SvOL+o2twwnwm8JTUr+qFHHS57WJpU8F6J09G2XD4CCRrUbEU7v7xB3+Oul1iD3drHxQtDHTASSb
cQ4U9Xgg6sI3EHR7GdSWAC4XWDmEynvj7MxCyZdRpQkmhHGhkaiN5henr4rXZeBqEE+hBgEFyDM8
0oEKa7OITIgOd6s4+QQo+RkU57KxE4/QEyEbaOmxHi4vVYDJyeUOysTYWywyZL7fU3XKbBGWBDaR
q3RtVxwsGsW/FjDpFrcHt9B/NyxVw1Jw7r4y/lMOSD5LiC1yDVOpO0rZbwH2zEnrUKvybrNAd1He
vyyz/6nDzHr19M+QD6DwBLE8UyfSdMo0roDBH2DPsI41wD/6anZm8/ZZDrZAh+3AeOpSfDOUIvrk
iaJtJueWkISk3CCXm51gjrfnuhH1MtU2AYlwA25L1Yt5WN7J0dIr9aioAVz03tBUSRa4QxjZtpRl
Wrk7rT1LqBk29ljERYqaZXq2Bdf0btw4DWFex4j8M3BYGPaI/94bz0NVAtm/rxHw11zaIqeIuHvx
w6bVGY5jEgj2eYZ7OWypeFRH2AbVvlTQDFpchIkjgfIJBmyn///45RWiaKybKB+/21l5HzqfhhfW
5A8XfIw0rofX7LeTid472Uj4qAz+BAN5we4PnPGDozdwvmw4vwRSEzQ1MfxOz5ROIat/sEHeYesa
fyKQ4IkwzW6V4261/1EXUyJczjZETJdjO0eIYBthAeV6caTv4IfV0Ns0Y8debCvSR7byxFGvTKVs
kM2Nz5roMvM7l4/70OZZ3rU2cJ3328zWfflVVFDdRlNaIdpZieWzh3MWCr0mME0qCmDyCPVlDTlp
fE3L56RdE1BLHu8L+MbOu/QEDLsLOd5DG0ry1PSajvpzJsgjuYHBLzZmiIu6MlQS59GqrJPulzd5
RYy/ApKtu7bMymVudzeAonNm29k1so/ij3SDzxuGS7Zum/3OdhJoJQgmO7uu4LDDM6Ze6i0cD8Bc
myBEuLGEZCPzWC3ayRiNn4sEPANh31ZXNPypCLMpA6cOBUx2KPRAaWrDoY6Gpkt3hKdz9VVIRFU3
7EhIoFmBpN/0ENMulfdLrdoAhBb+ngXE8jdndW1TVL6Ls5bwOuO0c2Z5/Pl7qpBz2Z9ZQmFtT7EA
rogOGvkBFhoLZXevHRwe7qVuLRfEUNNZuhxBaSbLGaElHzxIAMpCvzZA5g14WuR9oIEhNqWETvg0
3BVte+hQxvm2wi+FLs9RSrBgPngYuOS6fIRq/oM/YA/xXcborOySgEaOSfgPwcxCmi2WSBRkWnVj
NJStUf4ZYVMqnCrM47NPkVKO5aW15Iv9BiZ2FlFgwgxVqaxJQsPSG6kkTx/6OEEWsvU/hvA68yuV
26ZF8yhQOFRQNyAC7OjRsCQjaU1unruaEu42K1Vf+lCLDK4qCIW283iIeNSW4pOL7cksSOdA7WLr
MCxVXTYtGNCxhNwuZxOra4mnw3wn+ti3g/WUfR+U01CWd7MHxL0wcBdOK0MOaj5DCiPLGNEyZV3L
zcUwB0T2HqyXSJXShyAtipQ6QGxBw0/0b6fKeOR3p65hOLqZ4JOwhoTjU/+7fN2gNE9+9peZuO6I
7tQb5EEVJ6U+rFls+23pMDkV0LUm4NX6Hlz/p1bo1mGqwQFsmp+1ZGmfM8RK2j5qwyilVrOOlGsO
PSoO61+rejA/J8V1Djj+vh4x4sTPLvvxTkzFNJopEUL9t2GjR80ymbAHNcsmu8I1EiiwZJ13mImX
TdMh92r694MAzJaJjbwQATpbpj9cmuLbzatFTVD6OFnUGxPMFPSrSavWvBibq6QkXvOlIyhRbNNm
wV8VGgxKDee7tuwaNjSj4ijWgFLy9ZUwnBYXunUaWcXM8GL3uv2iwANb65xZGg9qjpRp9bUjXfs0
sN5OF6fEtHj5fIXL7xB3TqUJq+JtHE0XI1r8MS/g+CfF0TzMZshbA2cbhhoWwZxcMmp4o3GhnGzs
1RRVXtY1/UKjGoISmzUzNi6zoNsj21+08MTXuL7vmjvOEKqrvoe3kEajcviKF2gOesaeJ1aN/iQs
vmbd0ZFRV/jGF0uCz8rf+qzfv6+bVIClrceAi0GumJzTyDVYdEF6Ed3iorWtZIYEW7rooAIAVBwE
Xc4RD3Ol3m5hvvQG39YROYIQmRipmFY4n8nWlhGF+iPto9wXLfMPFKtXZQMbzJmUAhbDyQmv6UCz
0VnxQAWAtGaaOASpN9YMamiKgDe0UT2Vh3rL8tYWCAH9mx+zdH3R1ElBXUQki1bSFQ35GsVc6dg6
64FGq7chNpVke84xes+mtqhDTXZJkBC7QI3Mhz91PiQ4LflOAekvuYxvaBxmhbGMqtJeOWPFNvnc
qcrym0ngQgKdCMWS7XF25gSYqPs3eSerGrxFwFiW/I8PgS/UcYwo5Fa0tKXDOgAcaZH8nvryGWTF
j3JVgbiQUNn/PN2K2w1rVXIt6DD2t8/CwrPjal/YxFqsp8VV9P07UqjAWIJFlvGrfyeqFtrl1F2J
6O3b6e0HqlliXft0AdtSHo3OjZNwDgyx3H4y42NehuvNnRdRJzDIjE5v6y0NHf3wTR0s+cKu1Glu
RX4b9NtuU02NQmPl4nSEYYtk0EEN+GfvMx9+kpyprvaTmQp2SlDnbmmIS7lq8CX9/I5U42tyTHx4
jjRsSLsh/cv7IgSNy4qAgrfyCaoQj1shXKkOX7HmW+1QHfbeaIYNaVeuhmegFdP9fQxFmmprSTeH
gcmANhTF8Rm+2kT7FhcmFb0t+7rscMSl7Bd/8uRNID+UBEACyQkuyUHcDe0OeUTeMAA7/oNJXTj/
r8fJoKr4Ur0q9+h0H1hCHDKt0FREdwEeFPoemJjKvjUMxjqbRbl/ZiGSJD0PMAA2drkcGZdYjtUg
pB7ZZOp94Zg4EUtl7IWKGwjkZNbW+SQfZPS8r1RCiqhK1MXq6PBZUsSHPYuwlIz0MZ5k272A3sS3
ogiv31aF6ByHjnHovJBUuSNotO4nxJ7dz41UVZYfGYY0zDC/Fl2ri1UYERpzpfv82apL+mlbVgCW
Hz1ECUXK5i33QX354MIyscT6gvEEQfJ/lttKZ8xlXqdxcHe8PnxCDSlW8Dxi8f/CWTIjWd3qbkjx
VSeEgk66HziWB++4t8O1VwTc9pBbU/flpupmQnj762fllPXYfSPoPOk0x6nRIRTl5PSnR4wci4J8
UW5d1OGO2UNYpbM+0cZZzwbT1+rNBnQStJgdLplbVoJbPLHWAbcSyRYDNaJKnnaW09NcdSWZaCFB
aAbF26XNNvh0abD/CJdOwTIIu4Yv04GDZgSLR92zeP30aSZn2L1GtFgT3vA05f4+bx3h35+3XsNz
PwF6tlGlRZx9fxhKpqzWmHgzqBWaYO6HJoKPNjQtVnVShUkaawmxCSp3D4aGkBVY8sqpiQooTTCn
QS6m5qiIvsfpe+7dU38x/rVrgxiy8uYrdkm441GLU7/KMQu08GZBdAr/h40jPlojKfRf0v0DYCGP
mGTT12x3tyfUHFVm0SxIh7hpr8k3rH/hvz/X0rSpvcGNR/CS3bgc2pfcI/PfZS183O6L2wbovMrB
mzXt/sGVVYMbkoQPMAd+rJPHCcMl4N5mrH84/tbOyvn3aWdKfnfeIlSsmYnnf9NF5PygF4z26Xw1
yMD+UYb0wa/UZnLG/5egMTEMBQqkv53Efd65L7MMxKqS26kiiA9Fri6uqcT79VNiOcof6ARZcbfH
971nQ/LutwziPQFSUIVbFLGrGNkqYsowpbDmOY1GNbDX9h3abr80CifE0z2jROD4zmUwZ8Qvbt9r
I32WQBYFjDYtEWF0qobQZU6Nv0007nR72ThjSX5JalTCiHIuCSjU/M2oyzopPhgAuqlktNcj4xnD
0dduKsQifwPLW8NA21eXsXbGf97aEEyZBJxSC4KWvvDO6zZWFGy57uUZ5qFUwHWzzDAEiyrGj2eI
eR4bzX4koJCLPJN/Ve7QsuKll1aPIBrxcRWHTK6vjvlex70bPNRAYPckFiqS53AHHBSxe6BGJy1k
wbPb1Bb0aJpPMPDD+2yrMaPIJ5MmzSDpJ9CUVmVI63PPWF2Dda8Mym2ArmcHD6YHJHLpdIT1+oSb
5dH8K35eQLS00penPpvsgomlPeOX99GPUf0JObCou0YqcX8uZ9hTXks/AYAqwxhKMUXCAR2Cg0q3
9GJ4jl1UmymP8c7ONDUKJ5qWDwhGGG2PLHT4WQ3r4x89csTn5EraGGifjG4H/5AgqM6cVqx8dDKJ
DFIcs4kB6eC4sZhwtTBAsTim3yo6tOjJpaFjg/e7dMldQM3eYQ3AdKyYOyX8lfbnWurpacS8Y6/t
9b6tOxmdlqXAmf2n4QtYPQZBTPWmn0hycF9uP25ZWXgNhkdewIJCH/dlJQJkv6Ogrp3JmRLWOh3w
nSNVEEnCtQ5YzS0rEHkln/Az5f3S3r69snc3oPGjRGFPlhP8p+l2VKKSEEBHsbWxAwHiuQKSn3TR
XNbmt11V7nnRMPP7pqCcYc6AtqWS73m62EVROoZnrDLbreFB9FqcQ4IG2ik/T2rxqoRRtj5VoJNG
q/+CzrIevp8OYfnClBJ4dF05YBnkSivdHJnjNGrH/MGjUnrd51U60j7li2EJsu7SJ650r92i0L/O
wIvrrwH4jHXHFwdHI+sAvSOJYeB4uKgPBzNs8qL+WyrpYtyIkmGERaZUQ/pUwpwbklYVor+hx+An
5WNVYUcjkiXl9jDgvyQnU2B161gHkbztawuA38oeUP7g1iC3YKYinABwVo3530YEoWj4ofn1iKOb
JLf3XU20y9vMc5iN9/HgjtyGk9tZkZ1mlX19umN3oImCIV4zQifp9i5eXO8QbZrb8PAXffaYLc7l
VmWJHAwmyTOuxOLUPhxtPRY7bALAGq6h3cWPXQRt5Kl6Ukvh1h01OpQq6e4KeVxd/kol5u0COSIL
qN3A3POD9RTgIR+3oEXC4/Zv8qbT9z2IaCwBo1KKRCJzPWn4PuzTedZT/lJ+I3eiFFbaNczP0d2d
biCPSZdtXvYuUXiQOggHqHURvgW4F+0q2Vg+2qyRCREMeiJB8kHqzGELE1lDIliC8YOABqF9+O/T
6h23IZzPN+upXrqyVw0rs+m51i6uMPrut9aI7Ply5F+8D1FdN4yYQTNClJmxKbip8hOfnhTGKnDS
BONGx+ofgprvvOtxZt8f6VKOWcHtQW2h0MVHN3/9gVHECzdZr7vODNENP3xO+7VOoltIPAvZn5ZU
7EyH+s/W8T9fI07GRqWpHWKl3NHNwW4vIuSAu4wcBpYkAWlqfvloEk++I6kE/CRN5TvuXd/4r+P6
AWJPxRjaNS0kmsqkxQ2ZHnxUM/n/rtNmta8iSyM3DRkIQwU2tfcqtirpyJA+8Zhtd7jjz4eBGV7u
pVE6e5dU1FykZjaD8lIYmZOeGAzNMmMzGeNY7aYJ6SEQBzJLTgSO9L8Yyo10/Uc8xQVy6kMM4pZh
rf0biDPxIu8cl20gRlGBy/4RBf5WRKXrS+Eb+nWnjXb+c2X9LCvBlIxGUyghxReIdRuiZscCiYAE
TMeOwwmziAK+Z9kiutw/uFmpKCHvkwdoEPsQLzm5lbJaY52BwGbBbefsFPTBNot6rTa/luQvnlH8
Sh1QM2ttjLtQW5dY96bftSm1f8UNXDW+H/ZrDekez6b5MFiT8Q24nZe5T4dmZ6Pr6eSGNfBTz+bo
+eAptXRFBEGO1OyzGfLz+oTDm9KRtII3ZjqkfoZF+Hu05lnkPctqRMzKMr4r/OCu1eXY2s0yR7AJ
fj2J8Ii057BvNX2Erv7baFCi92bp5Kpx5knHSOFTfrqKFb4Bfg/lAhRIkUOBcj3fQ25aYk2i2XjT
4ZOMyLRVYLgqHUcz/x0e2TOEKySPrKYjcyIUsPMPrhK+IGBxr9NsTPMQyCzTaHIIoRNWFTDjpNQy
fN0JqdG8/d76QAnF2Din6yZNfy4nGKl73CSgrcQky57BobJULaX9ciwiZq+hS2FCJCNQy1O2oiL9
645mW2pedNBNz5mTr5OFqZRmsIVARrP4XDzCpWDZM7m5CFfZDo+g/aukRflJc5hwgX4SNHPS3wT4
8VJ1cDUZu/IopWvDxkM/2t0w+MXM6YQ1BjZiGdc5A0wuxFnNYQsFCFZM+s2ydNV+loTJeO2rm3Z2
kLOkOAK7X3XnycOK0MOrAdavYWO4HA4Cvk1UJaUZUYQlmoWQ/Pz2JWXIaN6KiMefYPPmTSPASf9n
8htkc7B/z7LO47YRNF0RZEEN+00atd7SSAk0kXQFNkS04D2zrm9haQvUfc+QM4RImHdEDtEI0LAp
99aHr0EmB21Q4XKoYnHtkmKG0ZikUxgN9FraDjWXRy1Wr+5K8dserHTZjhS4ijJxT4OusOcLHieL
oF9hUT8njT8nR2nHS2hUXyu8Q0YFg1lgeI60gXI/ZDAifkYV1CRnAQ/XYq0um3UNtdtwHgWE56E2
0+j9/jWCR4hlD8VGY5EU0mR2fJbt2M1cpjBcuInjy7SXlAXSXjH697rNTgj49ENP5Ue9OfGHYvDF
T6NorEFakZXVILwAdVXbo2kT9QhbA7d6Bfa4RBNsMA2hpw9H9MnjLkQdqbhE2Z0yINjpETcMAYJJ
9Y/P6B2TdCDilWyHsEoI0w4GmDAaY5kdU3KIvnyH43+NRMSsyqFU/KLt1cG7Kk9sjk8LPjstchIU
UrxuxPaZi6UIeyEmZWiX61t1Kilyp8BUG/+062m+fa3L7i+8X9aIZJeNTaSo2LxhQAQ9/amFXr65
ZxueKtcBkNUhVbUjpwEbOX8xaXA0llwTLRnGGdv1DxyJYTtPomOHFY9R/Um0hAKG6U8VnPbOD9Ai
g53nC7SJ1Gj/7zxjq0cO85OekV4kTeiwdLgLzRaXMXOEbo6uFLGPHds/cWK1HrsY40upeyVs9pMe
hegledLZYbkaGR52x5hmmVGvduqCR2YMueTmXCOx2Q6mFEQfPjPnYJ96uST1ZJgOajMHULfzm51v
JVKy8OjTy95ysgjDPzopPy0EqgqVZ9Cxh8g4HkCARDxet1n6jte4e/cWXJ728ZWFAOgDdCHB9bNG
+W/l6AzflNnXK1uj2hV2Bc8LV/gf7FacTIfdkwkHdafoLe7ZCdP7j7/p4QqqDHZuJyAYTtWf6zHn
TOY1ODBnCU2/bSbgGRaAMUtG5xImXM9xnYfxkKtisbA8WgjCFJjmz6Rc0BdLjf4FjOg1sgWD02xq
MtZ5QwkwyEjL+QwNLpoetIGS6/I3a2wFWq8fCF/XbRCmu9lEZ4PQoHnpuWHBjjKss7GYmqw2EYOk
IeJuEZiAzvAAMo1W/+H6SriEuraLbbd0FJEf5TEhURrOxfm8wUny94/M/hJSuxwC8w4Ww0X6mbce
p4DULRLT9AJHjF8wg9g8Q3ESRYNm4K6cfDwM2oBPtyLIlREqshghQy6Zlj9ym6hOsKtJEx8UznMd
1WxuV6iQWo9VeT6RQ+eDJ6Xnp/XnTTvlJukY/wBqiWdWADa5PvXpGrDSomP8uSYzkll9krNHpnlH
y2Xn3+iAINqKq8CJ/ZUSukQ/Jr9UTL25nAEqqRCLbZAQ3ZXeYaW7950xx/hzMbjMmZ1rUBud5GHC
JFQcNGj3ITH6LZnVFjg3lLY+XgkYUetlBNHp1Th5atGTJMAm9Db/1gHMQ1pbknFK/Zo8mz+mN7+0
j5OPwnm5OEw3ZNLhl8FJ3tm+Lc2le3lu0s8eEGDROTs1QtW1FHStxbfr3vlvmV1Wk0HPXy09/vXh
WGvXvLJAY5H2t2S6PQh7ojr9MA4nlH7WTirKEV6OGKFp9g53c7m+Lpl3mBU8271ua9GR2OS9D8Sa
Co1hOHZ/mGum95870JdoYcpsa+Jr+/RpenXu5awBtDF81v4rU19DBIJ/x1zn9XQUlrGDEjE/ZMHU
YI1nUygJKULThi06PR79mTlg1ObtYhtJbYfcjEtYEV//sokJtzM6Olg+vU4Fbe6YMZ+WOUf/Bi6t
wUSfbMOztTq9OBEbpCnG62v2t7JcSDjNEZqXfNCXSQJftO8dMO5OIQeUSmpblLGiiWDhbIyIh4P/
g8dhOSosyNay1BydYg1ZXljRtddJBRbCfRZK45D2AOLtHAicNwWt3jFFitvZud4ggqmtCvDn9y1U
IUdEK09YxSmsSdU4jrPPJUlItZvLxgDPf0pdq7NQUBitVApc9q7JYpxHk/xWIwBjah9tn1eANgWm
gQRlp7FRL8zivTVolDEBYIURDisd962uUi79xj6mndcLmETGsK6ApqBIcADfJvmKLtscmMwuzLIv
511Jp8y32AptH02+MeWgo82TXXT4L/4TFH6IlYyQR6VKA7XLHoxTKF9HYd5GGKfz4nQjXH/INmB7
3ZLiBIEInmYzbHhLTdVE0rtLTv7aRgAjoogHaqjY+a+0QrZkVRTqculbeYiqaXflKGKFidh2APft
WzA6DS1vRlDyzRXiec45l1uJDDtZeN6MqpKt58VMTavFU5aOh0kl17XTQm+RIp1RM6wUpTHevWKa
aZ/zc1zO+KmsAcCCjnGxbm7nrUkAHHurT2d2D48nrmQD/DRnG18WM1Xs9QLTNoTHhps7KNtQtaxU
7CA68gAeijTKmMcBDAXg26N7XGiW7pmNjmMII24wckCgJoQlet6CA/wKefn1Z4Bur2dNm7xkivNr
zZUoZdoeYLVgEpP5y0ZRWBSrCoI+UJLEXa/IFCcfXKJPGlXwSNk7WUA4TM1GUsxqCCULAU1a98TX
zW7cU6Kls9S2x+T/Hd4RyudimrfnawdRJbMx8/nOuQGO1ZqffGI5lfD+cqRzOEwe+lSpwK/L/FY/
Qr/0l9pZZicyiUUoLXKIgLhgm048Gr0EOySTdp1RH7IA7VGzcnnicHrQIVKTjxW2tmxCZyOxj9oT
9Xbh9qPU2TVGF28J94vZKPyXDI/WejC41B7fkAl0MPSnkw9OkcVI0PAZuW7wqxnXVoGr8PrF0MRI
9r1wJ53k/lk3eDT6/wOo1BsMWAOMCsgji3FzR0TA8FUh41QZDmOtwc1CoV/XOYOhx861cCf5d6oV
PIOULPYQyCt0cAdw+DIJ2BxqpgjYtwXn53ryI1FjVPZOfzVeRLqBd3sickx7wvwnDwC2CoH+oLkU
s5Gqc+FaCkF7uhs6zEdUzWBYoPkNnu6tjQHnpV0VSooT5CaX/9/cpDA4J5aY8+JXZPMgmFRK8Wnv
4PbttYjV6t0+WTAACvRCWfwCiWGjZYngyZjY/rsoSwQtICm4ZvWQBQHiwRzILT1bKo6uiYSSLE4a
rCcBGibpMfHiwYq+dMLYf2szY4q8tiV1evpaSxTP9Z9o3CdW6GhEvL+2Ufpck3oBBC08BxftioIc
DpA8aThHd/Av55Cl0kQnteEXT7gZfp9rVfWLjnpoDUVAwxD1QsujW5lzRKF2OzLUfDSsN2Sfs8TN
EFF11vGKAfPCfXFzGwgehQmcE0rN8FGp/YczyNTGf5mCXtmr4e2A+rlEe9m4LDaQm1ymh2b2b2li
aMRrqTp4tWtAAA7WenSRa5bme6XUSUHteAPCRw1GQ/gGcsyTYud/q631tWpYfIopnDeTUiZ+gg8l
pKOt8YMT/xPEVkW51nIBsZbZAjgDQs8z6xzQVb09TdIZ8gYkytRz6Ds7TvubSdxUH+wC9dVksac6
8HCJvd/lpzDMXh0RB5kaUoZA9FwyPmBXsdLKKBCkyCiBEpJMOFfYnnE7A+j4eRRG7762d1ta3ZGv
TBw5ncHAfT7dbWEmVqPe9x4ehxe6wmRw+MggbXQ0Aai+0SIu1FL5KWWEpg2nn0h3JQkxey1ULgeD
hrYq4he/0NMyz+jcozxsvJUYMu2jN9OU+V8fuoyorcRG4O19zrrPwhkerTRhF/0LZ6wHKByTZa4n
fK8JjJ+F1dq6kcrjIFQOGPuJzPqAuo6a2/L63tFKKgVF6POlz0aID9nsFXcxp5iGevZgBekrFqBx
T0wZiW0IUlH4UBR4Ugc/belKhhSHieQY3ybAvtXzOhOy4w4PnZeVjcXxEy8/+pYehqYU0hPQtTlA
OGlhS3SfcYYQioA5MACG2I9WTUfhnqrDJoBrwcBcJFVGLhjDSyGMIXgtgSaidRONNvcTywD1lkJN
LzYklS1o23+BtyT56MZ9QL0JFJV+W268N7NQc9Zx9ahXklATiP7YWca1OqZ2ZejCYugbZmGxg1Jm
UWPL93Exq1lGSiOlCwQDOeLY53sn7IZlDEe/a1DlSLvjwIcX+7BpKe8T4XM32XcCp6ZSTfi1JQCM
fNTOlNVrAmDyJPNSoJU57619qOKnQy+UoLK1ih0p5oUFBjSIaLz/K0Xiiz0lQa5lvStDHhSoA2lE
GbCZFYbc0h4dueqrolGJTML2XkKEucifL7eedzz9z6OlctjJnOmxYa+4Y+YaSfYm4PLFlRCBXRHj
UuYPq0exIvSSfrEt8UP95SHaWboKXOYND5WQD2dwtvjmrCx0BAipTFGk945wlBr21y/XqA7jp5Br
tgqncQZ0Ayhn6Wnr6O+1kePToWarKQqXuU0GAk9OSLa0/bGiyQZxY2hepM2jwUAvlHUaCcM+OpKP
cEyVWb3VZHl20btctatJqBYK5lpqOnmockukOMyTA+/hIeBhjQYGikNOdmCzMgwhsJMMgLwVW7iv
JaO9KmvFAqydbycOjih+7d6ou3Tu5cyJoPiHEnqaL/N7dtBycGHrJHnpoqIohZaC6ZKF+1Utngtk
hMHXM/cWdFtHmhJYU2FeYX7q3Famm8ktaV3pzlubpCp04txsOTSFpJkcrBEIMkGMjnM3Sf3+hFZ7
moCfiyRT3eb9QtCFRWv6wwSABpmm65QRG1HjpkUiMc/ZzfEmaHkMMboDTvueO6/MO3Tk95sVNmoi
ekJdLvEQEC1oFngbMvhJXsJ0JraN0Z7sPqpyBDTELxTbK6iRA1AFX2VEw+8oubFEqbX3D/H/oKw7
D1vLc6Hb6DJHT6VzoGNwTBlZO0EV854qoUZXWrqzNYvEUHUy9sz5O4pzr0itTfw08bvKqz+l5Ico
tOOWbmuCLYX8JaBAzfiKCwZyZ3HzJUXJ4hiJbvwT33ZSITMSPNJjMt0/h0zaeCNFe8fP3fZsCPIi
H4yIGQDqfAJUGYcOciYFO4eI8NN8NN0uL9rIW1eYyUfWjEiNf0AILIt7ms7Qv78dRtLRiBc2/xGr
ZFq2G7VXQHG8rVGNXGUUeHLg5XbSqdIgH6rKgbsVrSE9getBPLjaYR/rAOV9XpJxZVuySpjr2awC
WTqwuAn42hDyHoQLbJrx9SHs8RIu+yDiTiJXlxwUHdPdnbxMbE24ehY86TmfbDmId9w3ZmARq6nY
ZQAlkIDpUxPIbQxVRaZCHg+KlqWZfudDziTOKHps0fTeIMHZc9/qIouoSWWUG4ThpTLNnsLRynjO
23pJgeCBzQjAw8MPxXHZTHMFA92rdOiYuyy5GrX7ZHmR38BEg/wSlN+SmChDOgonvNHegkfLkURb
o9Az2qpudmKJFMbQAXH3mzgGrfvQ9h6OkPj2JHtLZZhF0HWJW8i364M28tXB/M6TUcM9a/Ukf6IE
SsPUBAAtXMpTfzQ3Xz88dWk3dmTm+/0O4IgJJbZ67UFLSE6qzQ0aLQSJgm2z/rToAJhZVJcTQhT2
JjgMGSIfNYAV3wCAJAVang5YLkhL96egxjx9RVqClf3870mXic+LOMu6aJ94q4oax1WraekSeR88
swf8rM3hBl6AU+O4s4ESt+fnTX+qtO40pOE5nt5AdV6eHeYPH0XLqW3T13PksXtLEIY6Efe0qF+0
agc1JEto+7NqTFCmsN2LGKYoV7v2zepHldIGXbF361nHp0QBkSJCw/+DOCTZsnhxcqBRalJKMP8v
unolCUH6/K1N+CUW27lkvXmp/m/a6J6WG8Zo5BFouuwK6CtG+tK9nAqsohhLIkeHiGHI0crctHUv
oRBzeu22fkOW61aJxEp02qEq6syXSx7/dYWhCRJGFCigZbhn03epw+bW/y3QvILakqHlcOemr+Vh
hM8/5ZUWv+UB0fX14SUcfld5cTbJViHYw4a06fp7UfZEavSbm4hADbjKr7uYDyIZRb4inJgV8lGW
3Mr9AMokcmoIwYrVzYBU2MEZ6QfrklVjUDNSyqGIdNoYqs4Mo8CJGnYtT/4pYi4e696yshAKJ4Yr
Hjh3C6K1RIDIF5sKHLjgYRm1UfMaE6E28VmU1bvsZUTNemgVqsK8fqkE/+V2BjsB6MtVidrvIThi
sjj1HL8OHKGOv3oyLg5RRuHNb9VhEsy40kvMwjQaWsa+5u0aXdBMXEIFpjr4lLV4HvHxF9JQDi2x
A/Erwewt9KvgZZnIKrv6jYRxfK49c7mUz/P8CSyClGpgMdS80waXWQzarfc5cZPR/nByeOMt+82a
f14wS8HR7Fklk6MBeZ8A0pHzJWF8wP8dPYNpwEoqqXYnzn9rfDwQIqxwF++UXeqiXAS19wBn+GE0
VJZbkYSsFpD6a1B/Uim9nENTWceeDgNm7wp1jz5U3PXxYh0fiXh1T/HTApHqXAJnbRAMyx5ZVo4f
glm1vaW9HZO2SxvpXWCF6I3Uc/kh1IBw0zhCn6uuSx9bwfY7VsPk6+uCI68Nl16Cqe+58yOX91Rl
VsS641bXeMVLeMy9S2VqbL9pU8UoDAPdQ6p2vZt6BhLAIsqbTB+XhYKGoSvBTvKQFzprWVktpsal
rglvRI+bvUjE5uCQ1S4//+5apZOcAlklH0AHSctqLe3rk/SCB/e2QvY+McgQOVaWItrtGgeF6KeV
A/tkhAy/JFgRNNpYuDqIDtn7fW08nAC93eGQvXrhA3hS4wUkKJDFOpGZQK1m7btsgUViB9uetbiy
SKD8BG+GBw34MngQfo4G8EVbOK6OLctw2cd7sgA2Q/XcsPDt7OhGt3Cq9yMFozDKIwzyt+P/PyYK
fF6jYzq/xZ4ot+aGNMTaXVb6741Z9xXABojA85+77faMsVRZjfTZYAfcTv80046wNRwQlNNxtXj8
RADi5Oy1oylwMaDpUB3uFVaDbR48TLvYy6nuKxlFgenxQbh6ED2T8uREhOw17wynnhZo2D/HFzbm
O5v5GkGoRbo/d4Y+z1ZIxiA2w/hIwhLVxmlDcPFJ+yKr2QcCaCBcxGQ5AQpiHlXlw6Eo1QxubcYg
G3e3L1T9mWbVY3p6zjoEDgoMp0S/VpyeHBpoKzqb/NYa5uquUanFd6VM9w+GpQcoH6VxDWRhOWNy
ZAIMx81siliLDG0ksjPus0hRtKQf2jL2XuwoC3WcROFGIchYroqidAGiWnMjdsQ25ftbJ+G2QIi6
Ewu57zJUf7L6P7HirCHD6F5kq8UXhKaifNBR9AUbtYMpBbB8Qq5RBB/rNLL74nyzRD0jY8J7bfSo
LGhxFISk8NG6FOsSbDcmOV9OWGsXR0hhQORkDMJbswcwtq6ePk6CUOX81QQJOzi+HLB9pSKTPect
/EFNHs4PEkqXZVoIm3bvfDASvflIZJZdX6wcOxCYx19uHYRDI/i+GfOP9U+j1CDSutRveBNZFebY
jBO6vIhpDuxJAj20FdAsMF/DhSel0mNrYiHsr8pMUuie/1RfVFVJuylSAnrtXslUTdxaXcZ25W8s
nQtcspdvMWgI9KuxZyH5BPvNLuGZ53La560NrPC9djQ80bimY17oehkJx0fQq1i3vLWoMVNFGG8W
eRpZNP0CpF/vW91Zqe4+7v6e5PWatYA3xdD4hVWb7n0j3h2+ZaRp3qzPWrkcOJMiLVgeKNRJpO/9
3wCPhe6d+WA32xvarYkim2/DIhOPARQ4vVRa/M77lM9o+QFtoQ8pr6/WrP6Dv0Tfq6b3+nDUZ0e6
4TuEzvn9jT0Wl5tWSMka3YAlOwq2qgXUe36sB7LhvhA86tGdEKp1MjhSJtA1oxX2r2pEywzC5n8u
umlYUakdOxv3lEoO/kUTXaDqLvxvQdbt8uDKwYZBYuqjxYIyw2Ct1142WyfdQrT9ciaZXqIX4a/j
zoX/NXpNHkik1FsDLQWuwduNgzgL8GB79SPpZPtNIdIriqmugjJsr/PhbRuxLDamdMe6Ltan7anf
xu3daxESUPiPpCf53P6nkAVFTmGLwPKtezMXnF7/PjDQw+nAfqbCtoVEnX5Fq+GZS0e3c8CeOYzO
g8125lXKKKB+TqibAvpbEFf133zrrzEprZRArjKMw2VvpA6NKUcs2m1Pcj0nGVYC+O7suoZg0I0H
sIB7g5z1bU83e4NruV7KxfEJuviOuv4vYnN9m7OrtP57CrnKJiCfHkaR9/SEm890KhMY7+4IYRgt
3f8FgzkVOQDNQJwGmLuy8weuUMlR02s5R+IHOTPElBUKi4m67OqwJEyX4FCBuSVhwEJAixqpIC3o
ep9tHweKhmAXx5gYwY68y2RT+RtA9fwiUe0eUuAM5DTHNrcZfxp+FQGEVOsIGUNdzTg1v69gLK99
riYuqK3ZIryz1uiQ0jovbVWgUDHcu1g23ndMBS5I8O9gKyin2OZ72kpYwFEOvBlIbgYq24MKx+AT
swTDP6pqkQpvKtfYoou+uhJqui7JUnSFf8Xp4ethua2ygVtBa8+/hi9ADpEOkRF+HHJqGBcfq207
L7AEI6Do1jpUMhuMGha4+A3fsZplRIUVhsvMItMninQBaWU0jXENQ+hqIA82ram3nbRzNhlUdjhH
TCoIxHJtD++KeYAJlX/pFtYLLHjll7hYYWVZ9CIj80lhpNfQVuRFmKGh4UTyIkoU4ab+tnVjpdhA
k46EdVgm8dOKXnL7aF0wKeVQyneG8s01CF6QEa3epHLbqqAi3ZkDDpgnZGQZRB4iSNgupOCX3Uxc
uENVW7bsRBj71NjlMxu1guuaOJ77Rfgywrtj+SiktsyHj518FwEGjRvLCCtaGXuMssVK556gp8ov
s/BFq4+rs2WEDi+ePcIb9LvfFR/xYJR/ZycP365k19z/F6pJtXDmkylqyvm57m7aZuLPXJQy52tw
JT//1+A5ySeUdwhfE1scarhl8Rm8qmfNd4YX6dMQy6AOfHhUZO+lE2jiPLdfh4tYNfIBgN8u6dpi
/g8nx38oeSVWL+cBuWUSe5Nx6Oha/GhVPzqPEYe+mxWAKFM4u9NdxmMwg8U7a4ovgi35jl47orMC
XMoZbazvqbqdKSICUEO1JSDbR/olPA14FEXiihcNrB008HIPIkbC1m02BvZ9/16bo0nywQo5MuvZ
4Gv4fg0BaRyGgufNoaPcaaI7P8i0SnSPt/haQLnQHi7/tTgyWSHskBZgZbh3YfEYtuy5rDgNF5Ft
9zWW2zs23wXOtvNb1ulAL1ekrx7BKpZcwIZVD+yxdM7QNCjhp+ECWuleWulW9RPJPLWiNSO82nWN
lSq5D4fEAlRCDpGXyzt3aOuq+a2zqvTJSL2q42mTyEJ0RmJZBD6XkRyNPRCt3126n3B+TXBKMDgh
5gnlXN+/iy84MVyeL2hT6Q0pt0+j2LeX7PSz8ERlYTYe/My4hpMg4cDnLo+8YXXmHwt05VZ7YnyU
GZ31MtUxGfPZUPQs+LzAqA9MOluLMHC6+25tXbp6GEY9w0wiUzbrl+rWQ2E5lJ7AFh8gZhkVyT+c
fLe2DVvXA4Xf+bAzWgHJCqQXbKEhg4JnHQyFofivgCtT/qy6eqWqE1l2gZIVyQGi9OMkdgwrV6jF
rqNyJmKXtrn6VzceQ8Ih5yg0kmH2jqbBtbpGgaFHAwKy2bFK/PBcyY2UKSMzyJaB9DA1ejqOa3JS
3yv70OgkztzoVtOdIJSs/IB2GYsM6N7sQb4UB9JC5V8gwMN6sh/EWrtSHtI2DGi4FG2Y5aLYshfg
m/V6R8n5hnzxdvHXdWLB+aunIBfeOSDDKUCLZlhHZMN0e0+WdastyxZeBtc8CBeU5+NpL1OEuPPQ
s1sw7RC+YU2B7pNIth8eO2g7U0UL5BRXjl6Xfr6XAjnZLS23xj59kFMosSEfwB/s1DtrfaHw3o5/
RSGJr29ODuBc0aa2hPZm8AO4WPtui2ICO4yKJEQKWQG1dAcPFXxUdMSd6j1d762v6BRdx1g6KTnF
vWfHnBjN8VjTifpp9utOBFY56Bt21YM+QuBYCukNoBjOk1pLAxQt9vD5i/hp9KsQq5kg76i2qT7C
e2iSt3fTQYVncniT/3rTC0bBFf+h0klxxammK0JYXYIhjnIDOQWEOSaVpLhQ9j+Ln8b8mboyE/YV
J3z01lZXpBCTvmWEQWpadVAb91wpKv2wkLjD64Rwhj+1Qjjpzqn/mLh7COaaQFCDUK3qwrKVPHy4
wF3ee9vvpHu4+/qCEI62rqLI6hebo9OdEHuikwZxDekuKGEO8805hoFxNLaRIw64Y83R+jgRlZe4
5jlvNiCT0NtKXWTctNPpYAxp9y+FevvQyfM9fwbV9PhMmlbTjON4Bkhm7X7eKhaTBZJJOg9CzXtf
85jVEJDVHnotLsMamQ9G/gUxysFyLKVoWSUsixYtkERMMZMABlsPZXo7sLF21S3MIZ9gAB0EB3lG
/Hfk/JQh/WxmGxyfvVkR1sst1/HPocYwcz14P0LZYAALw7SWXA9WFJ4yd8z5c5Es11um2n1RsESb
HGdBOSCm+DGIpIeAHcyNGXanZrN22+vhnc0DiRD3M2yQhiizwj3mofNBKAJlHKNphG8MuLhcf9Br
gnoMgzmYXf9nV7tICLI5ZSBodddU396k8/b2rTzXIpIxtkheCX/W90Pwt8F77pguguooiXQSId4m
u1xpRx0d+U228tA3SwzT5xXy3CFAZu9wm2CWpVOjl7ikEmYt6+eMTDTeqyG5en0xGyeURzD2K70a
jnivcopC+PZD6MQRuPZQFp9ZFHgFnT3vJ1H49TcjUCfcrlEVAORW6Nl1CYQrzYK6rd+VTuzxMRVz
aHQNN5qpyX0pGndsVRzbjd7zqLVtLvQ7k3bsyh7svXTbCINXktfVKQof25wZLWwSauxNRJ4lQGao
ZFPFdf5fRBoBerjfVya9I3CSszXudJd8d/T2e6S8CjOPwvU5aewhRar+P4lUzLWTNrz4KVkuSvKu
4N4S8isgFC11LlnA89Lo2XLRpeGIWODSVBRGiamgoNPb8u1mGgABJfGhtRgG57CIsSFOkmwnuItI
bp//40w5mBhlI4wdwK55wo2EzfCX3+/RxNvvc4kdi7Jptu6GmtFxnFJ2Pb0H6+sI+IKICx+hjSDF
Ew1ZBk/hTRv7F4YtnsIGepVj8DpLKqqR5xSEIjnrYztLYAwQHViDxGXnsVJtW+uZTTz58fIc/WTp
9CDURAArzK21HJai1Rw+bUCUzXFEIv/3quSIys+77L4kfGQ8uYImZ1Akrw5EawQuuVgYjaAZ5r/C
x6jtJFpwPCHiY6KoYuvdWSEU6EvYz0lIop/7YfSYEqEOJajYixBUUCKz3wtn1uTwPH5EIvsFeuah
uWI66vidGtE4YN3pelYvDwmfCZ7GB0aBlKvbpW3ozTNEvCY8nW3w3LJKcQWRQd0eliaDyY3mGf9i
Z5GsyYub3YYTuPhwEtzxEYTTzMZVJDiwMhISSWCdKLMhG2BZ/31Fb6RHmfl7k4lfL4DXxovLfiUr
EKXNQI2Uh0OE8cvw0ZOGKtc/f9MpvrQc9UmGAYxnSYY+GkR73CDKJlqSzzPF5WivGGYajxA9kHIu
AikzalPYY6p0VJJjemXJTrZia9ndFufysL+Y9YRQDTT2W4FqSV23bOLTL+phAamEPDr2kmmmO4rI
AUOR/tlRQhJcdj7a9SwKz/anoRdpIT07vf0CG0iiSDjxjVtiGBr4oi7QhfojqI5hPKlFRE6nYLzf
dAMTBAoqqHeebHqwyEfvrKBTCL5E/VRWUn9W7lJmUgg/PEZDeDr7BOxwPkcBO5xWf3zc2+8428T9
Kb7Bf/G97y31a5iQKnWxmGrIg3mHPm/sgsvs8c/kaT6pVO+zMIUh6D3bvQZI68DC49CE8ZuGHVVr
wqK1xPPRYyXS8FbGZzumBs3qyxGHGfcxK3rpz4QFDqqtNC88JRfWiOYHibBwhKPpv/K3A9vQP7F+
/Jw9o4UbUpGncAyW2zh1M0Dlt2h1tSSM9Qeig6/J45FfOsaJHS6fLIm6pcmWzkGhlWxe2UA8Na1O
i0o5PqcLnWjb+7+JgoOOXaiCgMKHie7EZjio5toRdGd53mJb9J4PKjQOvDRJ38kn+gPHMvl5tuiI
wSSQqHQt4/7e8NnywFHpbkw+esD4/EwfqRNhnR7CWa5IWn7pq0h7e2Ur7e4qI0JGiIggi48qtRmU
5zR3FskWzuZVa+tDR+B3YpcKWZmLX/NOl1mEXiPjhLKrAUb5acpQaOwOxvMc5oihxJdCZeMlFaqm
TGYnbGiXfEcoORpE43t+uPvgSh3UqUH0Z0rmI1RrYE+VnO97rVUXm281Jy9HSvEmK3OsfMMSZhms
hMPnSnrF/772eJK/7NQl6uoqbs1FnlIkW1fIaSHuAYrFUtqNo5d6IH6vvcG7fQ4TQpnqCs4x4nZg
TD0LDC6YuWcA314FBLVUEMBQKYWiSoEKqWUxylHtpI8Ib8qqVH8ioF79a+hmqAwdzumHptdn2BAs
AHJC/Jazsl1RjA6jmi/FlTouiBA5KXqiE/qEfI0vIe6Sld7uQW/nuYJ9DWqfoM10HIF9+7F2+bX1
82MDjgyCr44kdqC3hQsu0sGgUIry90ES5KYQL49+BmohSjq2u9mOBAeMsCDTTdWt9x7nom3WMm0d
PWaCesax+f2IYMBxlbizpEPIDLYBcKO4sqnC/18Dkt9MjCikRXh6cBZxBJG8pp4DHaEqmWKKIR7+
tRGKJUKj18BPZPJOgruR8BjmbiiddYeiv0SjjW8SK8zN9xsJ5Hretn/j0cRt5FOpb/6SQ3k8AUXa
tpbvJp2HzXcfO+IsNqP/mjzD4cpLyWh+ESlZf9pwtSGfwihId7IqiUIIem0qkqDbw5DYBmKDijWH
MBr1PcCtRqn3wqzd9ovZKaY8IqXWje/98bUxEtxKzZNyk2+1Khmcx1NnO0UG+ungbtMZe0BLtyFa
YLSvFe0N8H8NSfxRupOLDKdhIgSY008E+SiUjzCstA7+NoGl3qcmS0PG0skjy36J3ZXhM5fR4dV0
qVgdIICwHY1xzKC3ZktG+4DUOcYTJdpZIsrAk2jqLt3Urw2hT4Ah3SWKc/DbA1qbYkOEP4mR+Kzm
KQrXKXV2d11y69A9/dPABv6RNPhL3vAbOQ/k/IUfCsZCUiUpz4MUeBkJglhAmXU4aWVeJdEHHypp
TJ6RINpgXnev5g29r5D22/KNn4mAy6o+jyarxo2hVfAmyYMlp7n1raXUWkyEWs1di1VzZrCb9zPX
COnf3m9mrmwy/BEB3Dk39izdf1++Eo3dVL4OPSuri8ysIYHn1gHIx33j3pg0yrHOYoPr6QFGurI1
eX3avANPVOopiU0/TiGfY96gbvETk61ksagdlvNKWKcmhkQljQGF2eKku4V1jTrI6fApFDD0vNTt
sTurZ51RIX4Egobzkb+NRb5DcM29qoYrdU/234oK1IZf7fiUqePpLerl6xBDXRwuMZVz4/aN5EJ4
m4NN3D4a8pOQpBgmzkFnxEv0GUEGjwHh/w/90v5B14FC7ewVLbUdKa8BjMxcc7rCsaNC9PgCNMVX
TpYkneKutnQHSAjooEJ5i4k/54M1j8T4u9gQ/75D1ZqSyB/aa7NfP2sVlemZMN3oRXY5MQl/IqxD
SBBMR1UcGX9QetcFmAhQzDrdTB0A6KnKWHOjOHYmM45IGq3HDn6NWHlEb9AN3GpbtZcqmp3JeTpq
bdGHeGOd0gPBTLu7q0h820FJ6fERUKxTNKMKcxs0x7+KWVrOFLL9tuR1ohnsIGbCywKjyBkOZCLl
iVM16reaolr4XNHNPMtlTQ31CU6ipC/12+JkyhzRqIGWp+7ZVldBV5J0cRmTNcha/Vl+Xl1NscmC
1Ohy5ghEFlKI5t7e2jTxxNJ2xWO/eDNi8j5s0rHXmZ9f2VoFZ8TmCnKQC70w9Mz9XUR4BR25DnBs
7Yy9cBKXxcg9POJbA0JFMmDGEmGM7H6XuWNJg/UEzQ1TJdT7SK5f51Bhbzw5ODZ4Dj31CHWIy2VC
ZpO0wjQviVblo9ow1XOsZ+3gonbbFApp+aHornixptMgJLZS5M8vXyJs0ptTyqYfP98Ko57y0A3b
gPCgi0IurSTBYyaRz6x721do70GJRXLzB/PYhzq7Ezi3+hwv0J0oFzkhPFmWc9iVEPu1CqYqgTGO
HTzeSBVHN8EMYDF77KSFzl/Vku6ngQmT6fqWUfs8199y6eBnRklPrW1F49d4ewJ/lcJ/M8NwztL2
KWW25mrrgam3E5SViQk0L0R4lYw5hv0bsW+1zyeTClMHKfHOgAB3dRqeyYUH6jC0yLuWe9onKxUd
Yb47MHS6DT/Udmeeskb3uikG0eu86y4/ilqoRpDwx3byQVoSV8W756/ac8UsAxHcYcVQbqY2uqaL
VyBomQ1IUX534PLT7JPzclHxHK3L2qGfGy2XgTmMlYJU1pUdVSdTUP2OzCxU8aKJlyBjtqA2X+nv
CtoQqP1pb0otkTbkpVRGNHY4D6PpgXBZ03tSzl3wqv7kQxvdGss7cxh6z0yWA6HX3NvUR3XK5ru0
YlzuEapaZcEyJF1uziWeCLpqVikpeSTkYkuF29VcDADEDvrd5jw11/9HmZ7GqzOclVi4Kp1t4Nmr
SeoJzQ2XKysIOGjObF1eVF+9576hxCxC4QQvR0oprtU/OVqFrtluw44favYXEt6YQBzZFyCjuLY1
iJCAG2Uf9dcqnb+Dfux6ld6s0YHmtW+YWIsMfpmVRLPfB9dFsJFuTiLpWK3/jOLQi55TZenu3MQ1
DVQGEiJRMnk2DYoZKzS7C7wcSyBhlVq63GaXVuYej4u4VdliC5eSc+Kql6zNM9SZA577aUJwCmOo
1TJXJKLBDeOQaGf+gnhRq5FTK96Ums/Z0zB3pfFHUW1BESvO0M9DaL4y4XHo2DuJXiPh5LZZu5G2
/+szXgRR8M/ML3atds10LVk3vwzA4dx0Z3cDIZBL94mzLW8WBl6Kp2NODxk1DUEqOyb8lS5aBL8U
GKxKpY7oXhcOTWaqv63TShDcJ14PI+/bCAXE26OIv0xIhnRcRExzzShJXwvdgxK+A8rqY3Xatlg1
QkNUQj2GJXLbNDMP1Xc82kq/QyUnP5AMdlhnkK1vGGReeIjJzdhs7R1Tf7cycy32ntwyWsoubgAI
Fd9+ZMWMfJ3SyHo1/6UEJvR2m+t8XKDYPj2OZAuBW7sA9ro2DrHXW0zGxDjpkhg973K+4idpiBgb
LQZIMDsF3EOrb6kvrp/5n8zMPn43uAZyZayRptgYMFr20U5Q7V1MeIovIk208IdqEeAoJMogDvKy
ecnOwdo2DaEXYW2CHuxn1Fp5Bt0HBsmvYjnrfM/APnsurLs887y5IzH2f+YByFxskHfahseKnuT9
earuiIboDmLb8sJEpvk/UF9+iA19le37CU96NiD1yGFjb1JxsqSPjmKj8RDCUP8M5HprtZvnavJG
eRhfSpVUJoMw454mFG2kV30HisFeQAavcDq1GtCTggQzt4uQIUQN7qc6WVX8MXQQp7rm8/2mD1OM
Gmq/yqG0D3zGK4u83w0Q7yP3Nm7AxVcexoNj+cnRXIaPprLMVOyMGbOwcv9fQEqUNqZYgahykq9b
M4NQJ3yJk+OzruqPU1fQohtEO/6gHBx6JgbNpCFw4dBbYWRotcDaJJ2CCq/bN9hXgJSVl1XWwfxF
UOuf3r4jNYAwrlxX6+E2nqTSK3nyyhdH6BzqWMLa0CHQZSRdCI/tfKH4GbtdpRF+Ry1sZgmPYpG2
Sq1bIoqCYIMFH92seoTvsFAhXvoUV/a2EFE0UozQ8j3zewJyNPlhcUG3l3MZ/MF8xXmMOP6sOVlz
otDFAvoCuY/kQc7yJDKxz3Zpj5HomfAUkz+NFoILmmOFZeWOmQpp3mbf9+I4a5XYcMvCUaNCG9Xt
qukBCKNdgvTy+X/Pu2aSAVuJIpj/4zyitD6eiPS+Oht2bWTFseJyvORw0bGKN4Q0voYvM0MWiHX+
aYTHmKAGs6N0JcTruA5KLSmlVnC6TPZl7R8paZbqKvKVjA7FOMXS3cVTzTwOrpCwK/BZGGhbfsJ3
kd1AMlvC+NNxJp7djy60Sq9B0mMl2F9fQJ1fVbtGMx+w5ZyPQf7wLcdKJ/l7y2Av0fdoIcHz9uud
9V/Aqy07Eb5UGE1vx88sTfWozESPAnbJLDWdJME8TyaUJ+2v0pzGOHhkeC2iQA0xiKKkdUAALYQF
iYZHdg5eV+5eebfG3/FLEcELsnaJIQ0WwgHZKSy5niu533CM/uPEBj/38J9X0IkLdSBvzplGKA30
BuvhwInwHDDmGHF7nSOjLYvy3ICA8IWz5AS5EhpxBvpnLK2y97sETrHMgOfaDOdMAOkuRPx78ptt
kj5Fx1kh1oqhv6Gs2vpEZaZS2ixN/DcRFEDakmpdJZ0qLU+6jEdP1MnNOqsHaGGNzrpQ7BlbSprd
LyLIbgYqZBileR9DsRSuJaHcTplGOK8pSyyVj+Eiw2+t7Rt9JFi6mOy0AcqVv7lUNES5+LhGAMkM
eRxdS/1UEEZM/pyLecb6u7RHx1DGwCcQECg2268U7Rs3BH+9buyp64mkp5Z0/EGZPlwyTMiypWL8
JPU7hJUa1QNC9tyL0vXSpC4/HUWQVISfaV+xDTOqytsHkJi70Oz+LSf5eRolXYTVn3rKW7DPq4bT
zMfLJRirk/fIfyUCSwvW4QgkNjFqXd/aLVC4w6MSlm/radoGjkuKqknXupdLNMRor63AmNMbIUyU
4Wk115MuSoN6psjYsYL/0VsPxeG2hLXyAHfHcr95xN/+4xwazU7Q9vvKyPDcHMF4D23lypH86mKp
gMoD+kGozEZ+gWEnheTAetQMhJnAy3n2Oa6iQ+18yhf17Rrarj4z8KXOsBbeCD/jQnzyXrpKhhUV
pQyRWsZvqJ6CRtb5aFBaJyswBujxgYUHyLqi6J0WALpPRtv3jKmW8ujGF5fZtJQbYQzGVlAa7aXh
xGQNvqrN/3grCfhB997s0aLfrI6l7ldbxKAkRG6p79Xn+No0jSIrAhVG2VW5Je1FBlFWlp7h+DSA
6rAwKUbZH0zknyCdyRwzcWv4kwoXukdGbevtmEpGbKXuwv15zhWMWj0Qtcwl/nWOmwp6qyqaMeRt
txdyCDNWiObyoY8VqtZOFBmjqvVD1dYYEMpUvwt0PtM/I5xrCgHvr2WwceDbcQ/WUjyz2aiR7vtz
EpGavDZXhfTNCImiTb2tX65HeVmn/Q9norl9/AISma64XbXd99Pg/A4Mu/K35WRbS5OEW/Y7bcn7
7gyUG1oeghL9hsFLhfws7cTM8Hoq/7VzOGB7AkYDzxJbq7L7bZrUZYJYgsoHkAk6xd4/AUhJKEyM
/ld9dtczYFtseKVl5fS8DTJ6H03HTo61JCbOfe/o0kKl3EFgptOsjQ/7cqe49fSCsY74dHruNhZs
6JjvDm1K7a5XlH2hQClQWtTuPBdN1N+XRPcPIK+AMF4VFtXSld3cjLEpf28jlhD4Cx4u2mDgBCVK
Mk7pJSU8xYlf0vBdo0h3ImAIpkGR6iPzNDbA/DX+DG5iBTFFTcPOrEX0I7rp7rPPj6kG9beciUKG
GGvXKm0caLDvQA1bv1Yta2jQ7cCp6KAEiJGxG6dXoJ936ti9O1c0kupuc8n9qU/kE6om90jZ77IO
G5Wuw6CCpiqUoxXaBSwWGYz/cm9miE+wY/PVWXnGuU0lZl6ADV6btdA94eFVkVKNpBGWDJ42vk5l
4VL7khYNEbwUVMplv/VzOjHcY9nTSP5z+cb6M4iIqryl8Icx+if8xKsJjhkY9byGd/VCDg61njJe
h9cNrHkeEFTu3AkiVTBboDC0s2+BOo31pgwnslr/KdWSZ/zHWnNtV1ahqHFt93DCQb4RM46GNzl1
M1cFT8ajUN2Wx8NIGxjWgz47LfCTwtZgbwkfQxDuXjW2dBxX1DsoJKcxJFeDYVvkllMBPmYgvsTs
rQ6R2GKpZ6F0wpetLH4cURp6U+TSn7UkNiwn1cg7szwGu1rXZU4gCBa9rFe2wByenVK3ZnaiMtQi
Qek7ZyMFIqbtLIWbXlOsJJyt+HjPM+6wEdiAWoIOiix7MO9+ILStyzHzecCvtm6GpHUgiroZpAGM
vIMrUyX1HrB95Tng79E/PU/FYtvmTlvqemx0J0P+deaK67irekNMPsk1pjFMP9BI05zlmyOC813W
lRn2hWSeR//Nt+c5nq7GExlGMksbTZH2Wr1+laPRhLw8Y43W2UBRKAYFaJnhGTtIoAqjr2JV0Nu1
rTcOCsvSLb9coq6M7/WwEjVju0zmvuyoszf52SL3x2jJHZy4Qp5tIN7RpdZksE2J+2745n5MkReY
hdVkidNuQGfqs9/k+LWSTW1t4BiRvT1BrGESqpAA2NTx0NQ46c5RoNMhqDI3CgOAR4/3IHPDQhS2
sncD4QHA1FO8G02XGZ2K4ZJU51in1vJRHYFDQOksxkDSPUwYXHsiBKvehthy55hdDNVo5hB59W3g
rJf5xUgQ4fN51yVPunNcXV0uxksXDikwbgdqx7yJzvwAsfbUAr1VxUIqx6nVVVZ8fRdy0wxHZI8q
JfuXEWHhfm6QlAhTwPuL4BSI8bArueVrt5H5LQ6uWSEb4TiWueBS+55e5xoOAQoTfPAE6d+2Agyy
VZLu5LFd8HoxOmdRkDk4x06gSg58B+6FTbmOXHmTzFHRIAK3OP2/mMLKwiGxlSxun9tAFQaX3piQ
T39H7ADYYN2aM5rMdBtBxJc83NK/F/ib8F06V+RWnO6OsVOd0y5ldIaFEcajmahWZPEechenu1xX
152yYmriVFLQmIO1tqtLLC1d69W7g8ZSLSqChIPF/AzR6m5qW7mcoU3TfmMriRc0dvxuTTzR9dMo
EUHx/EPgD1LawyN10A8pyBfu/fhjCn7sohTVLAl3UQORTXvqvs1hAasMh6G4x8fFWm3bW04UXq3r
c/2IWlhvgrwgmOpe8vLZeXCE0/QIA8tszQPC9qKD0SThQTGbRObXONgOjZsNTZVHDB8mpGzBoW0X
HaaSTWw7gXX18Fe4B5DVbMDgk1riRtIITGZD9YiJr7bLmKns6F58JUEGLOS/dviX5ChRha6COKHQ
tDZr0QCWPNwjtA+Uqouw1b0xw0yWlASL91ZViNtmqc6mgwAnTsekCynKUhga6LV09Dig0/eBy7Uw
I8ghCin3FyZBe8MpWzFNzwyQkqFrz66qjHhPek9I4Z2BQt2yoXReMB2jkPVYYjiwIAoz4P3GDSqc
2K+YyiSRb6f+BtKFdiX0Nfn4+Kl6H8fYvCAjC9DKkhZI9qGz7AyoaFg82UbFoQboTf++E02kZ38n
suqQ4VqtG6J5qJPpzuamawRC3yniol5psFqw8poV05dQwW5fTj4/sk97V4BgrTcVSQmHGq1YfkPI
f8A+PbpALPUP/vrI36o5MKX9Vvoei7vHlXhY9iwxrEuFyTPHtSqHQtaubihqvpzi4uCMzbPMtUlU
nObDPAuoADcxcqThkJRLLxmDWtINaapuG838V+xePMKviFbcjG+8l6ikUvbOQ4+GDDzIezanzr79
v1T+9m7NlNCufT0gdZoDRcLoMwC4pjDsuLgoeF+agAjVZeM3Z7DukW+1xKEaD0Vht83gWyn+aY0J
XUWC9f4FvwbIdf+iekxqb5gjx02EmEaQE8jAbz7xcU2mzjEhtTb8FyEa6Fqw7kL8AL0NevY31clZ
4d+zamVe87hXHgKUPzJw5BBRoYiBXIPQdsH12dU77yks6jCPLr/it2REsqLhPSTXugPOb4BLwwo4
EXB7izb/Ldq9jcPnt6acUXDPdWh8hqlrtLL5F9dOWN6YRkf3nn8AbwTBCWIZxcpCT1X7LlA1KA1c
jiQbqO3c/tEqitYkvYSsk+vJNMOGv7hhNXJQ8eM7wFxTmnJkH3d3cr0JZX+NhAWSbYZAOC2b+/if
sZq8YQH5CKZOHDqzViaOwpEi4Ra0OGVx4VO39Jhezuv+LkD7ShH1K6ynZJUb20vuP+s8otpIEQ37
BLKRsrgdiPqRVTOQq1gGgu/Irz7PpnPqRqgWvRL+qh8uzmwPn6DregzNiDeWX5bF9crEcGHzI/4y
0vRFY2Atug/Sb/CID3xQJOkzbY0Qz2h552p5hIyrLJrCAVdzFB0NT5AUkuCe44qhiY0fpKCDTmbt
ACRbRAzwTgoygOhGD7zQxA180cdDYgH4FyLa8cGAOaZbTLCPOxoX9j+/FHd4ppc0V63mp+hV3rQg
ryIENXi0LRR6bjNCLoXZTJAxCVL+ZUq3vD1VsW/KsM9ndbl6pE+UQJLri0RnGeJlw9e2am06zQGo
UxGrHiJM7EjYb3gGqlKQBQQWmRTrYhjdIYJQUiB/eCrWCgxTDEMYGZaASJGIBUIZUxmqyaNoWgbC
1Waw5bcFLBLvPutipkyFRwPb5u6nA/9rR2x+I0gJUu1A8PWKus9yAojrWANFhXejQ15zHcXahskK
zaOxoCvbZcrP2cxNyGfDMoajS2jgEWhXEmMa/OQ4NBE9r7aBddR5EscHMCF+w7yryzRBO1o0Hy/D
uTlYDxnSjocHasXW8Ss9/2dA8kHFVnEA25PTR/LRpvu9GYE7H950UKrnS/z/AXZogPqPisSudzMB
MYcZoioEkGRCM1mrcLEKRWqI9Zp9cY2zxpRyPokzzdzhW0mWLDHBk98l0vy4yWYL+LyMYnIVSdjO
eQWUy4BJTyYENSBXeaHdMGYM++XaJbXwzP8IaJPvt2oRBnx8LZD81o76C9GkQWwlS7uvcgRUL8/M
BXkQeSRdZflkkyEmfHrSNOUFZ/GKoYb7TQ9I6U+dD8RxVMHqlSmYsiFM5vu8vuckKzfzbOr3c/47
jV3UIQXYkc6vZNx2oOaTmAF2XzRuXR0xwtTitwScgRw/VkOZWu5jdr6+0kHmSv89I2M791qF6xIV
5LjnHI4w2ZRjf/+M5Ur4Vh5ZxQo47nEEc3JhupR+EmtM3cznqIVu9ZyBKp9pkRqFWYI6XCnuObIP
ZsXYJOMYc9Qy1qxULKR6oPJ/RU5btC8KQiMHE65EXXofQUZGYDXsQ4r6xYud2FRw/u3APzXU74d0
ii52XwNs4kd3fjMTial1gj5QkhQVnufuG/36LzStfmtTqtrk5OMJ7NEbtrqmHd70iCF9I7jsDnOL
cZRW3yMgI/4caaFhMnSNp9Bh/a5DGh+ThKwzYCH4HBNprJLqEm3t9Wxf1S88MZJB9OKidV5oCHGA
khqgHoYTZRwdzbrNm8RYrS8H34taNM+E3bx697gysXN7Gcxc4nefdPgb3d3VpbnfDlMaxoX/FFsf
vNIrHMdRYYDChO3/HM/zzAAUKD5odeSzXsddYq9V0BdwO6sYt1ANz9MOG/ed6jhprGENHJW7sh/Q
eXuqVt3+ztVxxXS1ZeC0N+I5yAZ+ig0K761hx7uDRrHtntRT77HgQG872IxkQQQ5uehWQ7qS/WUL
xDN5Puyzws6YkjG+GaTpLQCxU6Qy65vSEtGeVuo7h4hn3coeiZxkDSHFR1eJsqrdEcG31qZPmfOl
RMU7MmWhlwTS85e65S6wyVxBF2ri6dOoA2zCCny2rq/QYBK8UK0q6NLOJx38kP6K6r+aaHzEPL+P
A+a9H0NOE1YoIURUhasyatCHUVplaEdW1XANKGC3Ir8lYzpEVWp+c4wMBO9jUrXXC//GvzLU50+e
LT1Sk8FeGo2rn9ZK8NvKGPkWTfAl4bVbqeblxiCETIRcM7JElnzz4aotx8YbPCHwWEbSq/9hZGSG
MULnqEFUSboyVcMm3e6o77TE0Rng78ptQCyTeAX2jsdVI3wP1t4H2yA1xrzW0qh48Gqjg52Hu1Ut
nzKLstmplhRJXoj6+rV9n2TmiH1oLHn7hECn4SfcAfKAu65BRhGiPDVNMbB6lmdH16PADSYOKAf8
ZJ3GInI9ua0zgN/03LMTfIr2K5xlSkeEbkUceyRJ2GddnsaAhZsRd2nyu6ey8CUVBHQKlJind75W
zmH1mhWOyJEtRw6zxZ0IM1NaaiHRKDXCsImUI1+EiZW2mgPqhdvKlORNilmTrjv2gk1drQzKNSjT
STyVhyI3bVxsEIOuYjToTBaBt+fBTEibgUP9Q+UjwgVjLj+Ia02DtVNhXqgfMGANvLqc09m/a/H+
4moS/PTab6b6MStlWGpREM1MwLuMU1bcrWf28ZtdP17t7kfILAiOSNgdjBe3yh5syNHDUvZJhPpy
Op4O4plCo+I3W0UKh+ynLCZ8RbRq62cwitM/PXtxsaGmjh9fIebEO378ytHZz4Z/qncvBiERM1N4
wRdE3iOX1uEF9JuMo916N/FHm1dW/rGLUtF8nYv0vMjUcAV3mguYPKBbAXrms2ezDivFjhrZVyre
v+Jq6HZP8fG8fFD9f9+GxUB7cQlT3xwGpZmXPJHLiYlnNWfNcQZ2dO01o2wSdLTCutqu+7IdBG9M
D+ErKeIdxFc9kiNbiHE08OdWVw3ZdWkxYnv/fwvyQiWNtuPUmC/4k6DxkXdcIzgV0tF6Iu8Mh2F6
kEipatGrFtFVoU9po0huCtVtBtPmu66rqtrqMpaPMcBcCCNZkc1tTIkEJAf58E7YmPpvV5PCWovJ
dH9xN2c+bp10+kTpTPvp1KGAsu/Rj3AV2XYXa9urQAnrU/dDQNVAx51u8SE/IwI1oGktdAEvkoap
kKNZQqiNkNFtYnVBLEBDtikQ7Pu88EX1OtZbpQYH+lMrRs+Fwh9/T43MQZt/At3NNKtgDR3BxmDp
OUXKxQv6LLFyfb5E1ZIPJb5Zs+ab1AxGy0RBDLKL2yyLOobBKh0JR+zKNiggsg6gUGPyl2aJQQ3m
8XwqOPP7OBQbfTwIxO2wKKLw0khPUeYSxt7aI4ExUxPLtOjLs99y0fiZxwXaWSee/WctiEqUdn5i
YmVKMeUx1tzbIQGzpWPiz+Bt7yOEfq6O62M/6O1khiF52OHZGOG53EHnUAxLptc6xwRA2bJXmMNf
gleVNVrz3LNnWtMhM6O+JPVer5BHtZo7GZteyztlvQwvl3LXdD4Znz2tBIYx20bp41xRd4LfhbTX
jQg9NMshcKNem2/FNd09wGH1tSQVQ1L8a1kwEF3oDALB/8M+JGueCnMe3D7egWtS/FmDz+Q16dAR
oIarFs4vPmxtFoTsyajhlmxv7dCt4C+EaDJ0CqaRJzDlHDCq+ttjZ+2y4JOwvKEeoyjiKXjQW4fA
37kZLqH2fgHQPSbz+oyNblQH3ow3zAKhuvtkYwWodg8nXc6DR1AIcRpgib8LLv3LlADV5AHZ2xm1
dC4wNllOd73WV8h3C6HB439AJUpGz6N9DEHOAFt9GuRcPuSVhRXOxJnbAk+usnYkLt+AVJ5nPoLK
fsuLCvLxyWOcIop4t/xGCVU7xHnYWE9W2ywvj/CrudLShBQjlRGqj9085SJWePARYukAS+cKBXXL
HbH4P/1spN8ADAPUts6xF84tHXIPd3oVw2hhrAduH/AkpGeFTjz7CK8g+po0tEJYJDsCu/ikrAbu
Hp4bNYzJJ0N5JBIfcX/ixmo1P9/KHHUC5FwliZJs1Lvr69AVHWWc2GpsmWEf5MOvXj98kdojlqDJ
AMI0ERa/H/G+j41qq3HUn6Foqzi1k7XT0m2vHnd1rNafvHbcVujpBu9JEEkzNcLZpcPP2Le92cr3
NkeITpuL0k06x89tXV2Nb7xSrwJViSsQLPfWm49ZvphHBfuTHZi1Ycoujfb3rgInogn3aaKHL5aD
0mBPAq1yzxNAJzo66AwcT/KOFSorqqE/A+ySJ2/FKdVU+uS4n/q6Ci79M+iL5msReZjv5I4XjM64
O1ldBntN3FgOFLS/WEDHe4Zk2Xa5r/1G5+MKISNQkxssqxObWP5qG90G7MLfWBZ4ks6oULaRkAIZ
zx3otNtxwfriCxosZZhCojVfI+oibqiRBXLF5NI0knYey2VUicXtvzkgF7R3RqFbCierjai0fxyz
SJuFvOl/Lxr0gEZB0Co+KvQ3K+3RA+WTJ/vu01fFSobQX8svX5oRpYx4U/VCzPCLY8ahBZuVBl/r
7GwiCH8pSSB2Qn/mg+TFqzdNBxUDeo4EwF9iCGAZr9a39lOjCsgT/kpC96QY54oo8UNXcNv/NUlE
8uoYOMcYKgNsH66kDALkWlaZ031eW+20uc0+WtN3rpXXYEygpbH56h0DJRd+cAtKY/+Ljka5BCrz
zqvpW4YH5YYa0D3NRvBKbnVNoIPXifnMHCfYirB/uNDP5UGvviFpDkkqmF5H6ellVEBiZhEC+oUg
4h/rpknMFOzF1g+kbUWrzwjNLaQ+eB1UBrgClmO+oDwk8ItVcWtwAWUh8WdakmEVlqYbBL6U9JWf
UwSA9MCITHfmEPuK9ABz5+4Kjz+j95kpYj6Eu+CCGP2iCa3Vii5pqoLop3Q5sxwC1vtxhQJbcU4Z
l7FKaK2VfCpynyNETYd9wMKSr7495oB6re3YnXERSlfr+BoFKSrZTGG+Jc30py1NrzpqaLkJjH1/
svtdgcZNDN2+u7G07fwyJ588jfqu4TFbHH7qnw8eZQt5G1gn5UvaHKAK8UUT5+i+Ntd4UZjPshoy
XT4ZXWZb/l0afihxdnt62OiiYzYpRumwd4Ek/9cGST5WH5GG3wG/71eHwVhDTA+xtfS1m80amqHA
+t4xX5s3su8bHvS+SWaurDbUVUkYjOg+yKysSeMHuCGR+OyfSwlyArRErgWYmBZDGNr2onSjZvvr
/lUY2fzXdCUPpMVz5eMryAf2rsX6BFCFRjRbvL5XLuasaQRPdl/F0b9HJ6UaxFkDW62bvFHv5nbj
teWcflL0IfChDq1cbdBzUWuTYBhtMgER6Hq02i+RwIqhV+/OuOw26uhZfj74rqhza1xOYOC5dhdW
+Lom98PjIQHnBKTqC9EqyqPgEY2ROUDLAy6un/QUg1NSfWxRHKrN+S+hGlT/vhkZSKZ1t/zc/2GN
bYx/HozVIKKPr2jZ3nGsVcnqcN5lhB8hFmGugrpIU6cVdg+MrnDGN+fv9Pd4L1RvWlvbhU9X5OXO
LljbM8JzWX9DvA2w00/X6j9U8DuXeqI8g4YAt1XU485ZelLq2263eL+sNR8qggdkZn96i8dvtO8g
brwkC/KnjkXIajJbbt7NSvehv88zkgJbHo+hrGHA0HHHz5s/F3ePJbBplRqM1Dz2vgyzViMFTJG7
bRu+5DvGi36JchQIabcAlwnHPtMt3/Yo8BgLZScoHWUAS6lkZFiVjOH+UL4pdNob9CqjAgCjAg3b
8/q4fI5NKDzatYKwpVcCDRxggPat8V4r36Zf+AbafjEtMkvq0rBlcT8pUuYkUIHa40UCEmMofvgd
X01eAmVIgvJOyYGLPbzhdm/A759JW6ZdOfWn+uj7Jld2rfurvOL+kdhK4DOFVFRPyZlHMMBcRRKh
yX+6wGZELs9xfQK7znpxzD7gv+KPwnMyjqhTzsvj/wZeOXyYAurgWkUoor+OBiaHXJMdqcpNncDv
eTsLMSunAMWK0f4wPmquX+fPd270zuGZlS4W0Ii5Yh939frttUP60wPrGZCNIIlqgT3tzlLianzI
vf1ljYzjxo878id9jqWdnPPDDi6oVRPCqI5YIlMB+Qe3AzMpt8DV2aJiGqUESdVxRg7ehQUkIxEe
Gng7+rfG75qS0vx/pILM851MbPmZt7bzQCFKqUqLKLg3WHyn5pqIt6Y2ja8oGM/X6O3/1nABgWWv
iYKCxNCIJUGjOob0O0oFKJSNdSleNrcEZv9wiaTMm6o4g2KJUiPV9zWPO8GiMik4URMI40Cwuovl
sI7xozM++SKpNMOiPWe0R4srDRO8hhOZUa/S/pt2sv39S6dyE2DmBEPn5FeZR2+TNwePERVgh6RT
JvnzCgSRDD0kyKRYYC6rCsfbgKcshg//bf4FTwHPI4iE5SFnWJDdQAHBuUIqe5R68WqVBAkpm7e3
4N1gAk8owv01l6Wfnn3G8RuaEG6rWZ9P+nqfdHH7x2QYIpiylcNFvDNc7iOZjHqa7XyCaLVV9H1N
8pCD+s9bvgA56CHOoIG7jOV33eVpq5R1bfGyCouU1OxPEsOdigUTJaHpT89sQlkZoxacKgTrCfZP
W+j6aTrTADjvg8KcBKzLzaK3V9vsiQQbmL08BhS242B4mNGScrWCR56r6+L2xijUoNCbsZ5gSdon
xHgp0FGB+f92RJ6WEUpoaTdNBNllJ2BKXkGvkXBHEzLXfFoHg2Yje9hx3OhukJVIGz3bsEUuQTa7
LEz6NpLkuHj3OPd0c2SdB+/9es+420V9NgPCPx8GaesTbwTe3esfDvDlfQR7NvZAgW/MeTKwgCcN
T09gBpGNp+mF7FelP0JMlNY1b70sr4hILbD021nOY29OWnvztua9BUnDwEHMhMnRhnK8lR0rxvpx
48N393G+UpvypfMuvYQCzRAlAFpTO1rPOrhQtFDfQMyIDE2h+2E8meeN+SSwxYFEZgOH57vEk8xD
jGqOarvxdr9BxCk8z896EXfxaTR3ND3VEZWOm5PcDutdhoKmdOnzBWzPskNnxVRhPXxGfwIufxjm
n6mHj+RdDYtfkg9d798yQC/WdarCmPdLnf+CV8El8EgPcRo59pP66X70wD/K3SPbIBrgpO7yd9Ud
EsAnQb/q0QpyQCkA1G6prM6AzoqJwSBUHFQplDxjkjXW5fqj0dhQlOjXmsXa3SMZXXJEgVWIp5/V
s5b9b5XtsCASu2AyHZQnpgkdHScopzQVR8lqGSERB1FFtk+2YTvC59BObprab8639XyUQOyBk/ZB
CDrB2I/6AMg3RRaW9EtLuaHNXLgVdAQam5P5amSqQIhqH73515NGYUT/z6YayynT5FwDSWd8rQKe
zD2Qxf9vXC6Q/mQB7vJZUbjhkP8cjdy5RXeIaJulj+li8WuOcs2PY5q/kepqIV7wtt6fO/LXb67a
mViQ5mLTNmOufDHTU/hLI1tgm1iDL5w8MVcdNHJCqS2UGSMyQb5OYafi5HSnBHd9m3Yj1PdQDGzS
zI/MWbA8tAHy3VpXAPtTKvACftA155mJ2/5jeD8tGxxIOrF2OGm3ZCVx4xqQ4McIFDHCgqwKQpd8
+QUeiCMtptozH+wFIINYuP0yGEb+1Kf7bZxL7xzsmk4MAM9GlUu/hSNwPbUksnfT7xYKcIuxYxI6
ADiO35OteuBEH457FaZvXcrFrwmxyCHFvAVYmPy01nxSn2KqSnvh/I/ZCkWeNObmAolH1Wk5ZSqM
PnxjKr44WFH3QZZum2hbuWN+FZZ6QTjuj0aVyocJ3UVj9u6T7GNtZku3J7l1fXS0n6NK8NZbxTWG
xfwWHC/yOwdVoXdrEwURnTCUgSuqIqDnwPmSaRuANKSkC6PVnOlb3idDZDXnlO6/tnWVqj6NjQXU
7bs9Qc49tciRBA43r1t2AedsBmrVYnmz9uK33F6/lODGn+qP9//bs1PlkaR29UREDOYHB0fyd7HK
OLBgGiYj/TAVTqTQPuxx0qldlfEOL54QSQpaVtLJ3zTBWvogSAIub6nuwZMdZSfEl23qeqBFy5d0
JtCI+j8/K9A5hqd0CWoHAKba5VEH1aztS6igwoBMppreVeP+zGCMVhiujzvs3fZlhsuKWIWGFCeW
KUUwA8s7f+M+HXjahIF50t4aWMP0APKzawwfbT5OenJJRGYYP/ySuR3zQg2Oc3sdqhZPnyYU/oKD
sL468R1s11KTjG2dd6pQaWEp7YGfZ79YyuTPqNsx1krlFeVTjn9ZqAPlRXHm3HhA6fOk8kPw4BHL
kvLGgTnVf+nMYCYz/SwsfUUNtTBWhpWSIAuLgZGHuGpLQ3PSaVZu6Tk1hgOjhfGHipVVcDt1w1EX
xBV0ztUhdGTsmHJjLpln91sl6a/q6jeM4B7k/k5pXiEBlcUqi14pMN+dApPkR4EThppbRIgWeSMS
9ODjEfALmLvx7ehxrSx2VqmePFJVTZKPWbZTFYqCdNyavyD6lYjsZNW0+vKyRGkasY5H8vpsXxOQ
izR/3jR+eDR7q1sCXhdnWPz7h+8jjMUMsxLzghg/GXjeHIr53onLCCgNSqHNkcwsHRnDPZfcYncG
EtRZDeCsD1RKI0urM+sUzCatQtumQQUF1gdct3rCzOyh2c7d5SqIV8Caf0n8iuwqWbi7ekqyHRJ6
IbNUzIAMeNLiL1p8rU2/Za3FW66g0vHCshz7KLuaeZ8bSVqLZdCgoF+0HwSffQ6fIyhngEfwlxPK
gu9Ew9IiTCkvmDjrLwcU8t7TwmJFHiaWs3F5IxjW44qL7mkTrFlitqvVU5uBR7iXtrvasyUsj/1v
3eGJoElnzOpqTcnf1P0izx+O3JUC3UFxTXamhX6oLMK8jK69mDMDtmTMRVex9kRReD23dxr9PgcS
B0kEg8NtYOomynAC+URz7zK8hM5Xi03dWdYQw2c+iFFvOC2Un5pV2bPlfs3cKME0X6dmciI3j/V3
0S1cUmVZ2XN5L2BDHiTVb7Tan4S4MOCFt8lK76b/7saL+dajxXbC7FRZ/TvMiyLzVT6nqRZBxaqH
Jd5WHmFMjVM/Z4ZLtEDKtZl12ZV37V6yIIJv7R4E/Wh30hxqiw/RCK2aTt6r7DrcZSUI92GXaKy7
g7lUkt6FgAdazIvNpv02qE6wsCcWs0GBt1CcB/2C1r1LBu/G6rclXtk1KX8Ewx5q+h8usGp77LPJ
emeibeFcjOAeWrJ069VMUbge21EdNvGMLLaKbJ9amm8GjZMsawUl1xHFV1ZXAxzGO+3FYw8tmbfW
DCPHmGJLFyYpv3aSbYMxXPzZcUwesI4qpZHcHNbiBm7DO7uUBXSohZOEp6vEMAfNSrBSniNgutNw
nwlZUom6Ze3ODGDZ29ejxr3tAsRIBjG9VIjStQTyhxGWp0a/erUthbJDJyGIWAAGWrsXrEdmwQRm
eIBWdMJoQVcNPoG9J3IdZgQfwPSC8srX6mBeEzMxAO2/HkuOXteo2yH4jXfnhdYLByQHbRwe7yXv
FcLAgdIQFl3p7qm/YTHypyV+ss+AC+BBZcb5Sz6tHTOzXuY/SpUiwuWi/NqKKjb/SjCtd//hSQIO
WmaV93fLNixvLUB79dr/zeQJVs7BsQ0DJsDgPkFbr+vsiYdnz8qgTZZ0GtQET8Q8TrrSIef52z9m
aeQazgButN1raPUKkAeoPa0monqiqPc0qDp7BwytOm8jaClS+4S9OFmWkU5EeuNVDqDlrTQv3ovy
yM4AS8sQHk0k0CtNzLWardaBGYv4Ec+edTtSoBum56RNWprXepnITYiz/WlIDHlSVJVM/6VkYNid
gjtKhmXlRKwLH+m6oYer0LW5AD7M0OIREUe3gmk1BBJbPa0NPYA4TQBesjhsJwDkZY5bCI0+wnuq
/UPueANWe/s6tAN0G2thgTOIsqp5/9SJ1gI+C1kN+IA3C4HC14W8aXmGq+78OF6sh+Cohq4uZ+H+
swvInmbMiE4VCSsbF8VoqlRb+ZF+EIVl/imya2Swx+SY7TrAcrPBZZo3gHlGYxRoOCffflX5tQXk
b5Ai6D4A2FTKHp/EWWxd5hdkWHIENopi8LBDFVYUwtR5acAE+A7x9i9GysMbsC75mN10lCk486HE
mclkp/AAa0+j6dIW7W7IJlktJ3WWnQnQdeRo4XbEBniLumKKT/2s/wabh1de7rQbNi3JKd0n7pXN
EG1SWSHSU0okty210E/0dCRXDjiBggYOAZRLw1+C2ftPGPEqbqS3/nRi9ZbXzp1Vj9sHWIuM5wZd
wFTrI2Q6Zn4PCq6OVrTMfsEP7pz/H1GK9YtD5h3JCvgy8wmHv8GW/6DJZZ/rQdjwilTM7GCMOUQz
rHdtmpJiY1XN7QVGO5fIy2RR53ykX8yIQ10e5DhM/Xb50l6aR9R2VfQpwYJV9mA/3Ztbwrv57Y70
rrw2QdoQONbxYUG1Zy+naPCcNZ7EEq6T+mSEh7Tx8ruga8XDpWbsoIB8tLmujBiAd+QCLTnqQSWv
rFS3tBnm+P63by8ihg5WQvadx1v0DGi3UikTyfoFCLLQ1mumvlMb5bQf6aDHQr6FTvuRf37Bpt+b
PTbLTRar7EGLe8daFEV7sLNtWtSWQYc+m79diozXQaiiR/52B4IMrrlZ5DBhpUIG23Eayz56U/++
UeC4EHJ3eo6Z2EOXgCLBRlmp6S6J6e524xF9Zqm49C4x5w9RneZd8GkVSJI3W4YqkT4WxDALKx5G
Vopby7hUEeRkrVbOvqTZ/7YHPu2pG7La1Ur55ur5VLoVNbWeMDfRjzSlvHGIVwRwVmycroq5Dmr7
ELIjOFSd2jcEJG6Zb7jKqxENhwCRDO+h8GbhD9+dnkG/eitKFT1Y7p+UTAgqxUvkxE62+FfU+Tyj
TMNppZuV04qcFg1eE3Vj7iQ2XnIPU3P/71Pg4eKL64qcXoEffCVwSNvf1x1PsSaqc66OJgTzBMcd
hcPkViuxJ+dy3kC2REND/hxdZuKBx2XqUHUHSvrrKbvZX96CXwEZyCfF+4ywnH2M6FXdjY+L4BBC
qctfjRxGxcTdFygEp+qGWQLnxxENWrq/LFRnSwSnQ9oCmHVkxh97uIwfcBcgwEEEacpKMwDHISby
jxuFbJGIMG+Z6OTkw4JsvsKbj9ZoXiGaQj6P8fGfdFblV++lwguClESNfZx+NQJ2tHcMB6k/y0QK
q9Epnfxe7rCEuGgzt6KTUNjGMbaBlQbmsytFJcc7UZev5slK9pTO5kU2DnSWklAVVdkU22I7RH2v
UZtGC5NFMUAS5Tq9WhsMAIDSkeObZulNcYaCSrVKelDl9xMWYMeCb7kwUXCKfrkJ0j8S9KXGU78r
NQzehAg4/BowS0qdnYiK/Bq9/y/+6eflGgXrzroqx5iwkw2rAjB54zpUj6fvUVtmDXxIoPiC4qD5
QbaDEvVuosxUAOUF2aXX9KsL5SgYKC9o5ZXFs+v7Gv7k1Q7DlqgMUMF6MKrazV85nmXzMpEGnFWJ
yjKvU0ts7i0VuU3LSVRpv7KBBpkOuRetruPi/cdxMevMkYIX6O7YKgo0/Z24VWxUTpioSiS5YfhA
WzvFY78Vtc7nPIEOejVjrScU8lhfRGhmMx4fi4J7fidI+uuuq2JVvJnmWEgpapCvz2iTaopmeiE+
B6JSvm20VF/M5zgB/M/CBMnt7sYgCiamVneeuc1Kou2W325txvsVeDC01v9RKIiXVuerLBNiN98e
/GUcRZEVy/86NtXFKg4bX5yOmVm9Pa43FK4K2nzCarIHJYjLDtWArIlkVserArsruc/KFc8a76Ah
k1JMVVJU/QrZSyHejRRrYCBiIcmvu5TNoQ1UX5ZRRAsmhQJOJdTb7zzwj4Gyp+5Zf1NKTwSqYjFu
+RdcyPflGPk5OGqCmaGvA78PLAJ3RTk2qydK6KVELdSNwI+do/nvRG+MYbGNIdy/m2w4F9NiBHaH
SVEzfXGxY7SbUt2M/w4nmJiK80nnwm3r8dgehCmbcQaX/vhiDn7h/ASEqddD7nIa/ec4llPkmc57
nQm8Fpp4c0UwtLV0DbKXDQmzAwTZM45lxeNVc/SGCEmywyomNNapWgjGo7odyyJVkNfWfQQWPqUL
iRSxDet0loDwgnUDRUlAbVKrHD1nJkumspmfVx41InzSADfrHe0yroWzZVMcNVvQWDOluRTyOmvn
N1ur4ki60CxDhqAs8GfEUa2URs6tUsciwQ3VtVwmWBs9WqOq5Sgv2ikMOty5Ji/PTzKGtqAgeeaq
+VfKTm2N5ULm9lH77OSK4qoAI751NcZtBvfjBg/1+ooFsX26EklTwry809lAdaXY3gC7mlWrAtlk
sjdjgAykEpuRT6snn6Q0dbpevubmO7+x1IZcfb3r9htD+5o6cgQkINbsSMNLkq06ccc7JPF8/e3z
hDc/vLE6+IrPlOzVeZWr6jwGlDjH6bKE7Nq6DuQPQBNhoeeui6946ZMwjywoqOdWTDVHj3zDD7+N
RD/OxcHPIX/7PIzR6xcaiUhbAhhqepPknZH/SXcSH11du0OPMW8YX/NH24YGSLb8NFsjGl3kG3Xb
rjPVrd5TRrOs3bj7oG0cT4sbuX/zylktS5g4ASlozdHFN6pqn7EO3fY1E2+8iFPALqck3Kl237iL
ska1Ff3pFEeSsF/QUZV9e0zGK0+GQ+V9pt5ximtFU2EznaGh/cp36FGX8TgSqk6pV4oVKlBNiX3U
8L9+mlPFdiCeOjxxVVORu0qURUYkHLkuAbuXAcutN0Bl8s9XIZgAAqIxV8uKJpAGwaRdH73N/8vE
7dOauWPlgpg0SqElCFmIkyxO/FPHZK4YeyY6oxRaHQyaAeQz4w6hLo6fyLXrWYB4tuIbDPrOk+um
Wm5FqImTqHRQzC8SytiYf6DAT+6viFWJuy1bzCbovJSiKdTXFyc8dBlo5zYFiXnvmOhK6dY9FpNP
yCxOCmBsJLf5NYZYcTkI/+HmJjK5oID9EBMBxcYaE0h9fZqMEdqQB26XKaWQK94SuPsgOFTH11pC
7R2mJWzRowncpwoVykL40ZTEPf3tKXkRpE714cnoYo4ZcZbBd2mbmJUV/IEBf8aINSaF145J2BZ6
+zHvrtr0/ZVZ8XjmbSHsPUPgaoN2uBXNrVOm7w9X6dj/lfaiosM40aKsDDVxEMrXSZ13EQlfueBe
Zv9+7GabfjxEQzZ3pJiZXTgzN4lvGkBDPmxqmEQrl1LWp+ZInCaIN6mGvsFSVZC59uS6bHmSo4Y3
Io+MLSjVYWvEsq1/UNGiIv1vxvx2hhuKh4vhEnvWWMUGJuHY7usM7lT+5P8fBbCU57Ld/OgQLOPL
4ZzHy1ThIWXDXgxGLajpPEw8yKIAu2GQY4W3kuZiZeznTtY0Guw9MT8lJkWMczXAff5+A9CHY3Qb
Zwa5AWJRmNjDofaBZOsuTo+uV0LcKi/JYDAkBEG4Bw3ca3HIZaQ9BqGzZK6JijX4e3Uz1BsLT0Ut
YxZRQzPgIp79DZXdlx/tjIhpkUlbPTlU+cLeDdREcb9SvcE1kE2bRT7tz3dFcyEgvNN45a/Ytila
Qg7lhmjQPiQst9CdBAirXYsat8TXNhvOp6jX+DExs+JXUdpARARbtBLQsnJwO3sWj4NMF3GcVrWS
bxtqpGMTY9zwccQenjV4j79ZLpeDfeOSE+7rTBIamEDKbOUC1mpis03qe3WheAIwbpUZTKU4rKyj
Kjd/tUtijVO2gCqjAJeyGJMiLiaj61yEE47MWtKG4osTPmDX7RqJ9PfFixa+60ZOTan2E96eO6hz
ql+IyP73thBgr7y2pdl7xpibBAjktgij3zUMTlDa8jM0BpxIN4/usH0QJlTaE7CTMrHqhJsLVvVU
SeJaNT9MmdsRv9iWJcL3UrrU8he0wkhHjGSm/ts5scbTmqfnrFCd1gfh2MChUdqoKIKBVwf2rrRK
01+Kl79W8w3MYMHb9JbnGBCSt55RxwjvWXwMe556VOUY8UdfHfZrDmQAglbt2Up3To5beUs3HsoQ
6hulr3Mr2SrfGRdhxYh/xYVxECw0IPYXCq9HeWtx0QD/Iv9dVP8iQpSuv5vny027MgyWmfRU93f5
Q2eIxCgP06eQx37Fqu6KQJ7iDlufiNlNKn4CgWDVNWg1eRX/uBxDEQ968P+GUTfDUhOW+oeV0Gui
Lc/bPRD5pPHgOIde9x22NHVMl7Wur6upGWUSUSJJ0LvbYr8dUcq8IA4qPRLnabF4me/Dc4ppwJPS
H2EbjM2L+w+a+4/Rtih3uPlXWW0i5PddmWFhOYuIzjrypSCLSR02M+vewqXFTTdfGeSQl6oogS73
Imu9p/vPE+xOTUkf/EOr++PJ/o9Ke07bUDW4WFqnu37/+vuea+pRWqgXSpBp2V7ldY3arBygdnPh
b9wNwzcI9Q7czIWi3o+D2nZ/UncvKJZUkjFW8IfdVLrRJ8HlBLzb8BQNuVF8qa0yUvLSOKaOxvUR
gpX7gNq1AFOLKBvy6zQJjR5I+EXLA7CyhujXyFHKX/c9QuFcPRREaqlPtl7r1DPKCVl5BTb01u73
UULwxrMjq+k/WN+qkBqLTyPduqaxeQw17+LTpoKBK4QSkFzY57tAjztCfAYAxjfDFHX/vWDT7McY
XZgColGO1At6EB4vROb6jo6pNusOW02skSa2J3+LyXwkUSHk2mqo/NuC+0w/ZIa86kGrbzRSIRHu
IJ3QGJPUvnjNy7geDEE/XCo6RsQEb0yZ7Y6WmxWR7J/Fa2n7p3WhyS55T7KrIiCWUyQlpQkF0t5F
x6kzm08ck7isQJJBK0KTabjicfVMFl+CMphhWDMb8MDHl5gKGvupxbv9AMZrMeO2O3MMMO2TvRBL
EHT+KecxLuuWHUNU8T15MNaf45BF+bzQOybFkJZuOn9yxsYezp8L6O4AeKV8BUFqTIPoQ6cP9/Ga
8wi9hEx/E/vvKOUYeeMMxFSS9dyhAQBjQZq7VrrVe7EqUkjW7rvofZahhA3lWxig9yIyXubeYD1P
GFvpwJPrBU/47FD87iVYaHWyUBVda5prRLpOZbCr1oFK35DZviT5bke7hhI0NQIDioqJDrj5XDp9
naNPyzrX5qPYRvxzY1IhORA2lN4apZFvttoIQkpUIrjk92oZ7HfYPKj7OCZ/HLLMxggEgATz09mv
6Gj9mVbCYFxVz5vrQ/L5GhZmDuvYjrJsKMaUHeKd/VcdLBeZ+bBkWc9UEgjhHanvNROjFDyRmAer
vClkVy6T0/A2bjDcE47aFefJNtXM5yc8+sWD8KPhVi7wfWtEU24WM/BeQBGSuIR1kmKdPawQ3P+v
8/cGa4iamSHB/WN9h1sBf3VCrpKmWKGfSxkAEPgrjSIcINVZJ2Xz1ZccgdjNsuJ+Pj4glO7sxNAN
6HHWMSl4jlmJ80K+B2oLFXYIV00tRHLEaxYzdZZI4ntzgVizTRGOXgRS5ADx8uuZHnmCF+GdL8Cw
Eh2KVf+IAQNej7hiG9uHOWfS2q4Exg0K5KrFyGrYe3SsWaOtOHuL1cDr6oPiPtbeFEMSKDlE2psU
znq3OKmw82H9DUIUeTufFRFj/C36YPjGu/2RP+pT+zDqsfTe3tMfVatSN40C/JWEnTPSdhb5v5w2
hBOULzqY4XhC46urtEmgMzhceuYNHd2lF/evLPd77/6HVCHHhr3uSTgxh15CHS/XldCeyI3l+GjT
t0wl3jlS74PgWTNL3u/KdNZOy9yxPvqTVX8oqZeDCJsZBZCApbxRdRxkH7/ve/sllaU0/OBY1zXI
h6J8bjL21fxyA5HOgyOdoNgx4wqabg2I0xOHIRNRuR9hy7UeU9neB+v0Vvt1DQqvVvH+QJuSVF06
FcmfBNRbXhyVB+IoSX7gbn6vYjk7jIgLz2IFXcCM6Yxojs6Vza1c548s3nOTj658RRiFGgO0JfTI
4JrGoXhSG6J4ub2v8X36xwfTvf2XNtcME/31lUHh9zTkcjFYhn6CE60kbBXEojgDfGoethoPhGU/
ym4RJHkC+vDQ0c+62Ubi6E2mUKaZARfv/sYeKDYmSb4J463WSGH0onE3ACiXIBjTcReOoIM/Byhx
mJW4C5n3G6fytKP92a0vVmfHONzCN3mEpsgS838mJ++NQm3LURrfvjfxUKGm/aYOfB49ulBjNToI
h0KLtkihYOoFoURJXY0b5pj6876Q+8g+jEXdn9x/TsD2/Im1Ku0x2l8zq8dtkU8hWLrQCFla8Bma
Q/BENNCd14BxbOs1j3QLOy3OS5YYwuV3BieLQn3yBAgeH82lrgHGLW7z6lrX2Uwsdh2AIu3I1H10
iGl9Mpnm59sQ02K+b8+K2kpzBPqIpFIZABpEBTV0yC05Ruie6ga97sVnMdvMYoG2WIh1WH6bDPK6
dfabl77v0aHzSaX3HSPzjfth6lwRS7b4WT3IfZYG3pdfRsZMggFGX8n8FGBv3TdFbONKoeLzAKNy
9IJ/h8BGCPEjCJklxAVKxHeDV4fL7EqRVVRGrSxhmY+biv5DFt5Y+992dXOlFHnpvgSLR3BunXSw
HbyCUrmogS8zGf6w5bia5CyV8M+5ZMB6RtF+uoLS0GZN6yWsiMv8EEfnPd+8UE0CWxg8m+Yai7Za
3C1xyfklMbtu3uT+OqNwF15GyCYZzGgGrm9Tcq8hQ/E30Qcxn7rG99cBKLUeFHrydoZm0QsHUnab
oSGvSpLBIzmRv3U8xXpBfgNuFoYoyP42Qf+skvZG7t29aWpKkTMWS7IvUPQD8domIRAfX153DZnj
FVH4IA+c/CLMf7UjjahB7YaY7nCvitKM1KdbcApTPJYSYL3wpojQdvfiHBeEL+9eXqhRRft2y4BO
kgD3bA7E5WXdo3AyYY3trcKVB0CCB0I+ZNJtSwZVJfPWkL20cponphpvOx+ZLUVbWIzr0MDnC7Sy
NQMzXJF7VVaRHEV7HbL0VTqHl/R0axlqf9tTEdqWm4K7tu2fjlBlxmMpcAm1mI7U0usgkWH1b/c+
jdsyctYPRe1r6s7bsy9dfpz4vYeFO1t+YCKHsP2RfBcEb+7sV+6Cph+ijayixEY4oDLKHj1+SbGM
rpdMLMM73ONg+TH1kBuXWqxsjl5WPPZ4T6oZ79NzfQiReLLZXhIU28R8glqNl4VV+8nD37SP54oi
0wBV59RP4pnvXD50/cLyCiL7rcJtCVlWSSaXsfl7WnL6YUrN+rBtDC6Fz1d4ZZSXwjxVCrDnGu7q
zHVyLiKKbwrNqxwE4Hq4ieKsysDmPvd/LSAOFOGqMLKPmUdEc5vJDrbgwDE3W330MDoFLnma67Xs
9hQ+BnFKDvzZxFWIdlVlXaVo5PE4vf0D6bromc0p0TS7+aK7/NVnK1d46E/YHPVkod3dTRV/81+F
LYhM+hqWCphq/HvAgiUKcpW6/8BznSwkZp7LHsvCSjfTVhUw2rEnz/EYwHkENX58ZMlBv2h/nW06
ACJ+/ScHCINeJ0MEWx8Rv7fOKwaLPfWvJ5xmV6Jcbxhck/xW/QHhCAUx2yVE7Lzipp/sz9wVhOnE
L/zygwV/fq/IBnEB0ntIjM2T/pqdc/NIJTbCz2WLqeLrHcU4qhjPuTW2ZYVy5YaK9tBehoWOGMma
UfUTd1ySo2auWj8hWMuqhTuCoLNkVEI6JYYQRXuVfVLrfidMTXWP6zJjiedzZ8Rl1m41q6G67Rcy
RKMNuC9pFLouJdkJYYFPWPDY2Ufz4lz74p4hQ8zHuPNtcg9QQgEZZ193s+9IAx1VFBE3E9sNzyjT
a5MM/YnLus1Myzddy/8v85dbyu56hZk76ZVCNGx2NY+Ro4/R/vgwH2A4xtocbdDucC46ZZGR21Yf
YG6ZZXD+PAZEKzMVvkKxJgByVwPsEGX/ICTi6BTGEmUMSxRtfiXu27geGjAhgGTN9o6CiG+oxA+F
SdVkaBqs4V2saAgI3sDq8ySDftZVn2wkbF8bNQrdOSARGR5xGudFR2ErBvI96CI82yuv2a8maCUH
pxSOCzuM+ebQzTjSj7c3+CsApG1KGGraMbQimX2LD1Zeu/An2IKRWZ22ZMxmOlmPT8sPWKbswByD
yJCFXJWlFALgh1QKrIrPSIEmxPwtpk+Re0ui4jtYHDuJl/HGYx7S5TEyiURugu/gfSBneu4XVL8K
1zm7qkd2QmUKIbZbD3n4txSv3irPe3/kglWeN4FxEjxoNenjjaU26HghRiJEyeJJ9urDJypPPQwy
6tTyMNfi+LOZgcaf3omWpNXom2Ri7yeLNWEJOIf1pFSWcCYDc24dFlnD5E0xmrP4cki+4QrzmTzl
LJDwZaqCsxFsqMdeCH7odPcwxWkPzpYG7kPmsKuXTfOKyoDhgLVOBo7kHalT1taRXG7xxYSYsiaC
jsKzAHl4M3MQLe94AFVlW9h/c8ZMvL7a/ModVGjcWQ9nvlzJ9b2kbU3CK8MVbHqZhYX0goPPoFhj
4a/vpUpjHE5W39guxkfcNENy7QtElfCO2xLKAzviB/SELUShmfrHzHovlDWipd2+XkJ5c8dDt0Yn
Wh5bk2Z0WRk3wXmbWLseKw5RWWUXVb+K9m42P4UJkEHixp5+KtGsHGm5gLKLSsjJvstwWsxRE+Y3
Kss5TSbfLZ7sGge9tiUcgjx8pgHWPSmkgTcYBG6fHPH+i3EYM8gJDGIbG7wbwMOW5ZqplTAF/sIu
mbDq8BkzBqjwTwWnwfbvqDbPZGLLOn0baSE/dc/tIRgRGZUCdJUZ1s1MlD3Zi02jVdvDt14Y1Imk
OARiwuRqv9VreNLTYmXIyqq0iN2qZfTiEz3zLb0dv1a6i3lIgk/1enshr9ZRaUB8RSsSyF3/Zqeq
m2pFtraqvrabxN/ycqogbxxZWAYfaU5xET7cZbRT27CY92lH6vXb5P4xjqRbEMheLZmtjflher1s
0GFGmGfP8Qe3QoB93eAZwDgfFQxhb2d5UgKOZADMN8WzUoTapDK7vwtxL9ZnHW8WUo4NtTCPMQom
2a99cyLWvdXfb64XmPIJhMv+bipeBKVPBVR0x4RCJXEwShSBUZFUrTo71NuT//hHk7F5FR1mB/12
PyqWyOINmxlINXwuu4+0IC4s/9frqQHi0b4LHYzycp7wgUOzqd5Gx30OPdHBGMlcaPkNePSKOHo8
CwQe04UDWSloheez5axOrVjnrx9bLSivRhezo4yeUwkwEHVvNvnonvxHBDQGrmVqQ8io5zVX/CIY
VjhW9H46Rim/uI+rsh2yRCi8R75wiCGDo2a3OQarg+FlfDNhEWJ0pasooDMpLGaR7Z21HKuPOXeN
LK9PD2jromjA+41FH4DlDam5btcvrCDgeT1BDDAaCCQU1lr7w1atQEL06m+nQKKtPQARVyqyDDTq
R6r27t/vvo51wfYSIq2hh5EyiGNUKela6z0W/+H7EnL2/xzVGGr01Y1LAJxoXLPfxFr8GEm3tRfI
5RDpHt77Y7BOkVuO9pE9ZmLFCmPoaNCHJC0j1jLlkgW1L97mtTxLU5I2hDeqWvGoebbZrEjWj6Rr
urrug6RmJ4sZe+FrJovJq+vYJDk2k2NwWz1oj36X6O0yn/Roog0vJbxGENNENt5hJ1O6Jg5EuGDk
wYUmnD47YsD50tQvSIX7fc+pGe7KXZwf+/EDXMBiNt9F6iFuK39Qg7sDNP0EH8IXB7FCx+ZcUfGe
vRSZ8ASVruGN+IWfzzepbYzC5sOMF9sjw6asnj3R6HycZEYgfWK/8YbDfL71xRAVhi/1lEi+t6jI
QZqQ6JlolFeBJ9ca6bIZuk1oiZxrPddFBY1IDRccbbWX17H2HuLGBy+d2RyIb3TALyhCmO5u3Lib
GQwa3idzXXZhLVG2ULydzzwvQ08TrCMxHpdfs15hjsj27Xm48SN8AP9JOjEHgpmS5fb+i18MUa4L
7ShGT6zzwiSQ8Y+cHbdLX2w+Pm/D3PqxQxnA+hdNsJcy/SXlocGynW98v0sK5AO0HQtbeI2VEA/7
ZZbWj8HJdzOB7MirEP1m1ZU/jPfJEpvs3bPvh1CNRtWEfXV4d7uVAt0scYU1Ia19kc32PDg88qpK
TW4SJncPIItlzTERZ6j6hHonrCTmJk5oAWzJmUx7mxzp+/mpNZ8NzTb4LFPkelD/i6ahibBX/NdV
Ngd+phcWg+ujL1Cj/QKhCraSqeD2Nndd7EsE1SdtO8ARvbTgepuwtOcJPFRJZA3ULDT7Ui1I36IW
1i52UQgzGKFPULGPqmQVYgLZLYuCSHLTYfqiPWhI2pFvk2RLR40Xd2oVrC5W8YSrtFPgF1rw+YlD
+YfPng4HQeNjHOmkIrz0ZLuX1ehqDBQdwBzcvdkJXE8NX1uVNSHpA+TtqL1HtIwfA9wDPbK1PX1o
4s2MQSPmEnL019vgh/HRQdMIj2f3PPJ8mTDC3lJl0tjNNJALZXbVqQBLRmjmnsU1K+kg4UwIyKhf
by0aFW41zfU6qIgW0UuWnETz2EXUtTFudO6/KQPDIG7njalKPAB4AEkBpWgZ2r//cJq8LIyK+kHb
1lEf+lINtqJxXJ1+sAdzTy9xiZGRZrbWukhm/rRUCjBz+Sbvb6nDdGtntR3kaRcv7tSLpN8nn9sK
oGKWMGkJWiJEkbnOmP9d3fczgDZ1MbrR69n9M+Ck+19Osv/NxEuezfDXvrcLY5q5JFQTtZbhWVyR
pKgV58cFL/WJRZjWs9hzAVmG8TJGV7ylnXz+w8yYydFY7cnLTyXAV6cyUKkw/9iL1qcG6+S1lUYY
6JrnDebnUNntykXXaL4fy7+fY6kRGa0PC0H7L45L4XBfah7WP5kJoSNEaM0H983Yytxa6eWK7ohu
5LbLiHhQNWzEaLItyOPVj8+AuVFYD+iCMQsHelX6gtEit7bcHTcwdz6BN3CJ3KkduBbsitq7eFkw
vRrbnaReiAxEJI5uPXeQLmu7GCK3yrGz2aAL0oNdMBGV0vCB3SlwDSRZTWmgvWxJ5LSAtkMvZFfv
k3npv34AN16PY1PLRJbB6I0e3HXq5gu02adbYoX+uw0M/yoexBqEp5NTwGRHUfjXqa6+MDUxs0/X
3Q8PzQtXN++hOMnDBuuqRshu//yAXp+/ZTuxVo+52IefaQ1vO3RZuaM/p9IkvZim5mPLR5ciFMyd
Z5tR/AS7hLQq/EnWLHK7t9C6EMqNuSZY4vevz1qNWN0Ni7hhJG8nU1xAGw2sxTS+TCj1P4HBIinL
OCJzV3qUdnvq7livcr8XiOYOnO21mTucJXy/lHaPiawEP7wnylKErzxRwL84dYk/OheLNAgfL/jR
uKpQgeuidXh4YSUXoGo62h3UN0b2j3+AnoSADSe6S8FUsYK1HJZCqW6KJxiqz5phIxR4/5A56RPC
uwWvWE39P4dZNOyjA55Nba61FnIQrv/V2exAkgHavSU1GlPTsmnublfX5x3YVCCd2RF5QUj7lQN2
cHidfr6XXw5/BeRuZ3P68AXbGZOy6Usyo8/ObbRmLwgYBbW7OnCDmHX4sO3iey2CVGmgLcboEZgd
AxtME5CbGExvtMlN0UsJveTgosVy8EUENBYyDr8fZGezRRql7HZckWjsOxX5wIuSedelb7iyRZxb
bUfCJ+kRFoP8Wq3KdatMi9145bxq61JpO3WJyTOqrWEJeK+W5Chnl1CHkkrZkZy4cWpj8EeksN6T
qIV5nDLByskqWKrA1Aa30+bjqzA7yK0EmkqwOHbdfcO7X1/MUzF2BjGFLJ/qdxUwKxAkPCjoig6G
KFWQl1W1VxQBAD8I4U/jYUR7jqGg3aEpYiQgjmIj8c+6DnEPE/LP4PihfJgVVTR/W1UB8RW0+MGJ
IJVvwUmESscIQoosgoWEznWK0I8CHLQuHBWlmNUEL0+HBG043GuPGfc44IlcquV7P7ce1GpTHM19
47RG4qc6hTgwwRcItTIXM/mRFPXDi1x/+gbU7TkjM1GNFZQ0hkqveQ53jAI3GufVGkiueRKmPUGp
gfDi8uPXOGWkhGT5opXHMGaeLOuzK6ZJt2rrKBe8dHA2CSqjFsA/hljels5qu4MeN6sgGJYlc0ip
u7QoLWxLNyFOvWbkPRFPyLENwEy0ddJHCaVMylI2UnLdBPvKmNsIRYJnTCUcnEb1F3UOy/s8KOla
3NTfZHrelrS5q5EpWNWP1Jub6OCGti+DMYA3uSeAWLd3AY76mSweh3ed9BXkhfv3ZOgcupmAFMN4
pGyqcrUemCKiCeBp2IemppNqp2Q9cu3+igud+Q9OMnt6qAtk/vOFsSBOG2oCoA08+jawFj5xA0qW
oaHwlWfuFxFfc20FosAv2u3WoGdjFsiRYkQ0Ej+2cpU5rQskr6mRlLDCg2QB73itAqZ4aH/ZqWVz
Vy50ljfnZZQdA8ORZ+fsIafOZA+fyoyZA8aixmLU93u7s+PNqq6ySAQjjRDhjvXD2zTGQRNY9VLM
/vTGdqrYfe966CYYzjntR/JswTe2+fecTnh3yRlWwck8HeoYgmadYO+c0yL4FinJg2phuJMw5a42
ZIYT0L04SPP6Ao9AGwN9+SwsT6gLavRhltrbUjVE/2tgldwMyFYmDzR8i255w0cr1igh3sy5yLFT
duSTFBOy9g/QzYSnyFrPebIUGag/6oq131w1z82n1sG6onYvmXmcx3Up90GvlIVlc0f6BtbVaO8j
uYMJHU1uLr23XH+IJ4Va8EvXOgVKCZyMaLAHrTUAwRGNPJNvkr/UGzIR540bqOD6NJnargLEHLT2
Q+V1a1hWelHnk+lMd3+zfVXybTPl6mI6x66t8r9VDQkGUWKlwzvkgQK7zdFUo1Yh6kLjmzHORRzJ
/EZ/RHzTbzWWcK1HiBYnYIn4AFc91QXTDWhgrNIABvKS92IGv2JOnbEfaQkwIiN5Auxwx0MTS1a4
/PQ/n8UEtzDU+9lpp1Wfz9Pv2sWpNw4je10gjQ6OJAx2JWZbPkDdrkb2HjwYConOJGl9Ebz0srNx
bIgDueFOq/14YpIm7/lz8qCmp4eLKao+gM0BKlKMnhJdHO6oAXkK7QlgspYvD4h0uQBOsMY1ZkjM
M+Zltek6PefmZ8fhUlGTpgrQydfZxa+0yWj18FOe7MX14ShjtZkF86JBws7jG4+LTe/6yrGzq9jA
9U5B85nRP8A3pX+m4gTk8do12PnEMe9HYwjbgW54eXjuInCbmm7CwzHuznc4lsVc34rkTouzCv+W
bhCA4k4SCzMO+1uRIWRTbedHN58bbaIKS5UsSOzW0zQy6p9sN9znvh56k5jGxgSDWqRqas3+RkiC
+6JReodsOYkVvIJfLYOmw7wqVAf0ypXkraEhsNCRLD28dI4ObGA4/imYLE+s7P/hEc5BTDVXIX52
bITcmuSjOXJyvYAfp2YWMYw2BCxtlSaCJhCs8sCpz4TYnCY1qix3Nh08pFVklgGcYdbwTiqzfLm8
lthprXOGvqKKnyxPoT08L6rc/f31athtYZMfMI8aN8+oPrx+jHe9Iq4cyVEXQrfyH17BSWTxmpvQ
crYOF6ukwYDSnmOBAjSdCG8UjHY5l1YzVqpXH18M1GOm8zLuqsLVLkdLhub8s1w3J5cNUxJTfj6l
6gNXYHX+8hZySJqDT+H9fedh8sOhw4wD6mavoKzb1wyGjPkqpWecnc044P0xCIh94G+0ZurhwWBO
e3eUoaAfULliLL9hwD457aLD6/KoVbFnF5EwTebodGuorv465dnzrh+ieodJVOljl5OfP1MsivBY
2+0n/UN1NOMTBueGYWQhTWPLxh5WvD1/ANsG8RheSNtOOA628Fid/NrUQqn09COP140Di4MBMgmD
VNmdlCsUYndVEfjmkr0rurUiSwm6dsP9W2IRhRRDOEoJJ+HqEX/YcoGzd1+SO6fzAaMHSA0W/meW
UWImNXUmUBtwNjJYDJv1Ml/pmElNdIcV/QXEHbSPIeTR48Wg97/dzNPlB2QYkeYPfb+kfxvVY8he
E++P0H8LF/HsRbyMLtpTE0oM2MvUN7jSi+Dv8T/KR/lIMuuaOZpOWknOimMENOuJCa5CZLLgiyam
HdXMJkPI5aemOvfj+2eZxt8sZIKn3YRFV1CISCmsbIoUunH6cIz3zHYKOukOlwCR/p5n9s4JVuIy
bqJH3WdHV6SYNQSNjMxKHBaxommnYlVrvqSp2zJwd6u7eO5hCdrL3XUdAFKftgm3kGPUUVgzboSx
RU9z1dQ2PYe6DTXbMm6/FnaX5wYiI5csiMUvaOF0itaTFGwGDF8FdKkzcvbhz4kxA8IDZXuvO5kA
vAtolsAP5wJAc9jttKyAyDOA2TyMz1szFUo75YeMwjmJQh1IiQfsy8zxNvG6H+a89v2GfY24reBO
CLTO8xVp9r6Po6VnpTOLVIRxsQulw7RxMUQWetLi9z/XayqnJ7e+ejYyRgBFFj+KE1WBBAYg3ptQ
jc9gcwGRpDigqLB1IIZp3g4wlxTjX48PoXFANFUG2hdVLUVqv2NYB0eJ9lQme0zhcbyypql8Cv07
aLzz2g9wUPVsimO4YMYh5gpzxGABIF0essDHFXNNJnziBDB++txUB5wdJdMeekK5U72FLXcVVHIZ
KnWVRf5K1g9UZu+AYQB10dPuZkk+Y+p5V9FMj+SIBn9mikOQSMj4npWwhTSn35KSEDpk1b6G+xXI
RVDL9RS9j7WAUmUPgVx9hshJoLAPGTlzs1XDpBBuz9SOLbi74qGGOhngCO7Ob5rkNLVjGBU2mpLP
NW/UQ7JnLDPjd0hO3pj6wNnGhVjyc8LkKysNHRxomT4/kxOpFinHiko68qwkcjUhahs7kb8YjyX3
b+LXjZnk0jFz01q6wsWVQFIl8H9/qfJMrIWR5bR0q5FN2aiq7vQTYpVKsVZ8kdft18A8I3SOe+KS
VsWrFx+0i+PZSUBWY6NxrVkn5r6sx9sVZXT9fHJGVFbeXlTy9W//jZsUhLMnXL9JqcfAqSuGX33s
Sa1lb+ohyRe1lBzZdPEyqCcSGCd3mZLXmNqGh/Ob9YrO1Rv9IXD609H1rNZWWGckw9RU+YxCjV9W
2Af121Bkes/mQ6lmqoEgZUesrisg9JgjF10WFFR3yvrz6d00QCMSKNr/Wdk3lExsn/v0Ie5HUSv7
0Ww/2ypjZEO1hRdiJfvJtDk2JohskoKmoZiMx4hwUWn49nAJ5tFZg2vanNxdUec2u0VxYERk4CQ7
hUxNNOr+oum5fXXexnOLlMZk2kMzOSvY00YbR+bvkJ1hnhIYUxbfwAT8EdmTlPLeVJptmsW6Nf71
Ow1bRh0PqAXKi9T/wbXe5/bFiCA9F2SV2uM0ROGYA4bHUG/xLCeXYhCZNFkQWOLs/0LPSDb8KytJ
X05cTL2zpPOaOAi/nH9piwpxZKsHm+nKMm/FIEbHux8blGksA76VZTsinEN2CFor5BhCmgxmri6F
b0Dq+aNQqwQ9ZT5Ov9bEbD2mvfGxAh9UdAjpo2u7DgBaM5HfRRONz3fVX+9RPXIxA6MAo9FKsCBH
SpZX+D+gBVHegyXCarzNAkbKAeKNSHedaIKYWJnJhgl+QXnGGDOcV9LfIMaFFEtq+6OYirWYrdBa
BF2NJzl2K62EUh+KBEC4JytGzBveP9pCbn3K1CDFf0CDGRlNG5RwG6BfOYEespIAdlkO6ZjaVLK9
kZ8b8l5JVO4XWs9a0LbSs7yPuTWSByJ8v5QWX1RARxBmmIaR91oJrWwMu9tdZPHNFoeYPKVSbRFH
a7Eb8TMV/DzoYAywQSk4wFmjbSgLA86opSul5PM9fzTqr/OzlWqqT6D37H0mh/vBHWOa3l5um07e
Cvs4X/+FYs7SSzyfvfrleuIFh3QborzccE7jjKrJsjvTgf3SokXchZO9Gilk9XITKIxGhcFZc0G1
ANLW09L7oCsspeDVtceZI0a0VShs+6c0+YQm038OHNIsxH6MZmQ/4wt2G5M4JW79mgsBsRwbIJTO
9B+OZoYl7j3w1EO9mFqCaA6KjgHIiT3IUQXz95190dCj29JSkJUziR4qkQmFzzEcrICVASGWUrXj
nwLPYdZVzL6VzJ+h5/tdksBOLX/44/Efiy34yK+RoR3e3zUBlfxIgbziMrCa7uy61dI9f7axNNP4
265fC3Bdvfz9SSVZnbiQNmM2u7GdO7dZq7bcdY7nccP1OuWo1iHjRufbEJE4EQs+8SCmiMymXTjG
juFb/Oa49vBHOVF0HQBJYK4PK2jFhWGL+E2mVC/eCqEValqM9E/rkoeiBUO21br3FZnG7kVATSbL
H/uHx919ulc0llb3VmpifsKYg+IL0rlakGFpUKx0XFskPZg+deQ5FipEv6+rB1q/szrsEkA5AHJL
EmKdgXsTlfrZCf9YRFRp1ocXZ8TKz5CIh8Dw9YWMYNG9PSnnr0OJXqo+YKmNSZRC/4i6/4fVBou3
aUiQzn632EXiBbR7lnNWPYbazYZw8zg6cMwrMhR8OtFH12DkQ2nANCMrBMBY7whFy7RKP3RPvk6E
kQo2hcDo0B3qHoe13zaFkCKb5lFJ6a7z2PK9Y98Ae4jldjVf4yFr8/CA+7rzYlEXckiui6TGoWyg
XkN8kLSaRQHZyR3rzdRxnWGc6ghsdpJm25/974ybwcICtVeo469iAzsoegHhUPVFXd/huTAi+dxh
mVRrdAgp4Sm5ehgQnBPwOvX5BCIbBKkrgL4WgcVYkrxedF7lAPREWYaR3g0n+XGulsDKSBHXV0zC
P350hQeAVgomOcAi14iN8ax4qhi2XplAXd2GvMokOPsJdiyh8ExtM39ykESi89vm/NnkkvstyUdq
kbCx8IRlG8/tf60NO+ecFGq8XO9jWhR7bH4onWW2CFfHIg3Mvc7hqQEMS/MQ1MozJeDMqd3DEqIf
EAcySD1NYeW0lbqvr3zcDMpGVA2eBJsCDZUF/WchBbqoanhJQAz/ferojFoRUjiTWviChAQLiXd3
sUDUgv59EQcA2gOEVAQcpXzVDUv+8xZMRc7lF4ak9gVe7OWGxjEYft1MYdOYc1hYTV32myKpo7XD
ZSxGe47i3SkqG1CccXi2cdG5NSZKWK/3mprzUz7nh1KCshk04qZrQgD5lyyPCiCOFkFmOKg8xa4i
XBE2AT258obz7zrcHVc+Bu7pkO3x3L9BOIHrwU/tXhrLkcUMFOg2P4aRQ9jEkv3Pr/qtjrUgOTjz
6rQjUlQQLmFpkRWKQGFnZWUNKVimVhlrRtOh97bTIgmHbLIDHZ1K+1Ia8H7wdWRGWZ2Sksm9dkXk
mLGrC8m1GzUCBXokBgE5qNTTs8wND0cFDqyoBQg0IZhMoMWBeB/m0YlT9Q2y2K3az2gUpop/gSPK
SBj5q/PE46f0bPMG2cH4JDtGnrjokEZrvsnzTkdSl5IqXj+lfVPm4PoVsk73xqN8ZpdzFSqh68eq
d1B2SGaHLXa66DgGPcPxS6qXM9um4TWIgz65tpr20ME6lPkFhvlPCqRzkR5Cnfqc/bdh384FQw2g
pt6H09wdSibd+cZmWmCE3SvKw+lPABhg7uYxrvXBWkXt60D1xPUoWAkAF0xLTfeFIPToMTVo5H3l
6OKIFU4ABRkOJaS/pgs1W1H9rxwoleQRzEmTZ/npOuSx/duizm2H+Krj6c3xSzkHFPCFvlKxdFRs
8p1HEGTNfg55WY0kV/KUqoYpk8WOS93+17Z+6I83KcXLOxQni6mZaAOzwtU5K5rGtBeksv9pZv4V
edIiFa294pBbddKwI/Oq9136DwDLFErCaFvH1WWjF9oenguLrYCxrzlWXOwNtwspFqEPF6zwEzk7
twSAEQfitjVAbCC7IEAOpo3IoSmRf4J5ZVrkiIUzDwmztzYN26HQL5EB+/JPMfT1jSy3B5KI8nAu
MGGFcDI8WvbuH+6a+aWR1oqNrR6G5ffX6rbR5YEASDcdQjjxHul9b9mpvNwku+J26iQDH/sKUcbg
c/4oHvsO4Gg16xBFTFPJv1Wf211jx/ZknIz+cnWD8CgqmbU+Lg+mNPTVOXdJF2X+F6WJAcH5aEu3
PjnkxYNVDvF55FgdDOV2rHxWp2dMwnS0o8Hh2J3Tow/aU1HBoDr4Vz3Dn6mkG6jffDu4T/+Inpvh
IL0qE2ZLQV82RchPHiv+ogVO50essBtRHw5LiMaKrrAQoSl7b9f+mOT3ZnpRBYXFAnYYxunm3uIV
LrOcPf/5P5Igvw2yXvjJEulbsDTqun4JWzPWJiiJkj2GqdzgXWgbw72Xk4/iqqBx2mZovOBeLgY7
+PLRFx0sV7jKc9myCTpl3TIL+rMCogtBRVJghIWkRQc61TEiC4IhxsqRS/npZ4kO/3o8UW+4U9lY
Z7vqRtrg7T2Bm5nDZpeq/bkUip+xbFNSezgpY0ImkkXOOUgP7/wqbyF43XAyiF1tyf95xING56EA
tJDYKsJwl86rzzCPj3k3Dz1XsGEFQr2OYRRC4lWO9glj4P7dFaySYYuU4jvrMyBOmUK5EIUPmUZ7
agkY1R7ya0K+L8dDsGn0gm78n1Du6/ZNT/241RHtfJMrprcVoF0/0qe6CVaWLujrI30N4nkrYSzz
ikmz6LrVKnDoCaSyROsQk9JKCSS+xWvpSKzjL/RLWkqvONfaqzlGVI5oPSLwM+r0bEDoG22miegi
VacPTLQdY6deFrTCMvchaRjQrSIZKUPyhXCEEMoIh3p2QfANpR52Qap9UfyvLLyOWd4kn3LD8jjG
sRcLqD5zYPUbFwAaMXD7sArQBww22GLcccXhKpnxdZlcGcW0UXnoathII0bCsbeyz4QKA5A/SmBQ
4sM7NH9WoYWVtGhlIc+SdSEq81MLTmp1iC1wkpXMcj24h+vRxpvS9fhOAdJt9TEgHxLkVgIf6o8l
bzeHH7evPkth1DRWm835Z6UKGP4h+7q75oTSdSKgEZtRuxdK5dIXFn811B5Aif8/z8FRAuiCIDuK
K14QR5ULWPJfMrDpSfnwV31mSuJYZH3FyzdyjxV8KrO2zWHHR5XhN/jAM2ghNM1tmpBc+OAyCl60
aVYzYRKjpxFWaPfaSg+DDDxDLXRsIFKWcGl+CMZWOuLDjkUMzzbmg6ZzoePgwRXzsmgkv0BjJHBu
AKtPGe2HXysIiyF/IiI3Sikez71QueA8ypXWVhVFhE+eqMWziCRa1tLyP95CfADFnzzme0T+Mc6m
l7HGCxQaGJzd242CK5WJ9J3drZRv/Y59aOVQfQaql0U5AmplssTPLSwFMNlsu4awWdwUTka4WhSe
B0upyun9wArRvm/uVOVMoNfqhOaqfQRTMQ5Jm5EhI03zoDkcoCQSgpKGyiHU2nkdtLuvcno9P8KA
UVVnd08QIVBuK8ycUmHynyqDB/U3jWOoBTLCNOCEk+/Zj2pxGzzQu0b+73TWJ+EEAhFYTSrwWT6z
JcurHm2lNwu2oTZ6HS+sL4ds6NNuNM8gChSmvwQ22CcPn3kuUohproEePm3ZyQPzKr7WDzW2aOE5
mJ+Qf5dkAMrfydGKhwlYk69YTVdnHQofrJTh9G5g3oa8+DGuzup6vtLgNKDGVW8TwYcNm47ISTcc
k7SFXqaaO6oUEvFsy51SG76JXYe4CfFTkmvtq3KWE1bwjVGHN4QdKEGnsM0OvsRxywmEaPKgIxrs
YOq43QDQ6+HfAATZYJXDWOI7io0Hd7nZlKC4Ue9GWDwuDS8XsBDmj3AKgBsq/71bI1TzeYtMN+EM
4UWaMzj1Owa5/80KzA4rpmSbF5Vq62u310hcUVtPeOprF2wbSUtk6ZcIzVoi4O96L93nzmrUt0yl
q9siJreuVCMV5zDxiKwv/FNxi12zjADSK6FnGhfxR5smUdqMgttKHud4ymoUPT7eTlPnx4/lfDzo
+rWyCws/nuLF7dqq6K3pKPgZm5hpz1DGy/aplAWDONqTgjb3Qs3yf14dWP9oyuzEM3kQx5kXyNgo
FAtsrjgNHVMjcTA1Ku4eQ0lpYAvmv7rLrhpy07VejlBdJz5PogYVQwF/D0/SYdWYflAK85OoppFX
IM7btIdh4PAFYqThx3UxfcgXiNjPV+eztKLMDRFFIqHKPXwISoMdoPJy0YcBHuHE3SFzBOQ4WJpd
/Vd84cAHVhBp9H0sWhEDysEIZQs54y8bApAJ8FFVJyuJ3ZmYCjX/YE99pwKiAOgWl6ZaWeOvBNkS
ExazeRY/jsEVryQ5EEYQW6Ol+4l6cj5cIHVhzLF5Ai93cTtLWdGs/rRTCvHHbn7QGmVCedmwyR5Z
QQJ0FJCMVJYayo0zbRCK8yHwtNURtVRl7Lbd7pjkLJNF+lyo5ziP6ys8A3qf37ooix5Q4wSCf2fO
ClAE+L8z2TOTC0b3dQBAoDP0l6wfE+0U5o344Rk2dbP3dBCNQ5P/QPcRuIt/ke6AEbAPXTMUmvwd
aS2QEur6xpLQjNYQCOkckQe9m4Q5blQbWRMccOSsN1tzHtXG4NdtOKNozWIIlLF/JB2ZOi4+8d6H
TAZeGxZ8k6jiJSezXr9/Nt+keC46U3uSi/9MeRdV4PEbvwZV21x1p0AXk97DgN5ylq+aUtNV7U+h
pM8GdWjvrpEgMdeX2SIG/3S+7ucLrAfx4ztPKliW0JcRj71LJalEaDCOz5aCPQy8a5ZvyGeEasxo
sWPEwD5yYtkX88f+3LYXhH8qfVdSSJ4JcywdLbbhF719WwGc7KJ1/gCFn2MIaGpFXN1PWku8YoBL
vFZOg9tI85zMdNQl/rV/WRIEL/tfWn04ACBJgdX7giigaVGUn7daXh+1ovlJDB/I/QV68yaDptqP
gqbhGEitOOZZW1yDqSN5EjczOjW4FBunj4sx0UYSFr4k54oETyUsIsEM/9zHCdX3Zsg040o8j/to
2d3D4gulEpaCJyMLwvEpsjTeiug2brIcUBuXMYc67A7J4G+6ZbDAg8NOgL/deXTG60yA6j+F2EKD
WTk5fc2ICiVdU3S4p86pdKeEgDVzpxTfbl89AIBNELhZ3ayzaZ4dUcxA92OmZuqIeuEFVP0JSWP5
dN4JPg6tVQC5VgTYIHt507t4dIGG7p7Q6/2YgV4b8zqHb8Qdt8fZytdyxYw06DCjlglv1yFpLHW+
/Zkrc9GOj33qdMfxvhxvFMCOjHy0avveidcUzbM1kUE/2Z0O+qhrCojD/E05Y6aEAw/zlcRd4aA9
deSwIifupt7JE1iLu4ktSUTmx801oBZvUU6rPAWKHObL/RLhnQlEGz//Xyk09bXTeHm4TiyfcTB8
KmTZSqF5uVDZxcogtV+7s48AzM/bGaac5m+ZvG+dmN83XhXHHjO9ztFMKeEjVPxxdbkKxcHcwaiD
55eppr2Emz22Nd12UIM3K/HJk7IYx8aTvH9KOTe1aAvxTslnr1YTQkPtgfRgNaKLYseXvoxNkZAX
f9xJfzMcPQ+IyLaLcJjgGAsRLpgnBXBZfAjXUYu+mkbWosOPdDTpS8cdkkVZY35+2zrVSEJWT+VU
RlP3rEPReMyibPKk4J7q1oZdVLX+EzEJLZ2snduGjKRbEXdgtWY2Uk0Zoh2zD0z21UjhJXRbptbF
tTUqeofDAGKTNvRHfoRrDtHBdfAROTy7yPORELRFe/9Io4U0/vNPTUivHHj32KZzUmOUGYt8flIh
HlrMs0OaoEC1fyQbxvKoUGziRycECfwPkdBpVIE4HvuyCgQjJWLS0vYy1iS9GTTy2vDN2VO/olol
mbBHUr7cZbAeK82Ljr4PXfv4Vg0YfVQ1b6AVpppqpB36sMfJLPzFcTb6WnIWFXyVhTYCzhTGrxs2
J/Drlx406s570qnR9M+RXfyN/vnCm35Oiv0hIPBqsTf7c7i9HrPlRdgc567OHb2fUKBr6AS5PDx3
3OF/ub7TggSSTSOtqg6cYnq5O5EwKO8om4ePK3uuAUPkTw2pquToLxQAdfXGMJR6lrypiVDJ63aZ
r+jtg5wmHv1YabNIWKmvOqYyCmgErJnYWuBPvb59P+t/ydS9Mf66+gMWNfWG9QfubpR62naGDZNZ
1LgOhsY0mSj5KRPZwuFBaa1Xu+2zOiBS8ydlVe7V6ccfyCYmXZZ/9n+Fn9/mN0rBsLFCG0QVo1pZ
hopdeYfqYKhnG9sq0SBnbwNyL2nceKEmb0dXBP1pK7NNCv9/6mloXSPase2ces/VZZQO0mGf8XPW
2rkgn965OzDE0l9sxrsBSPVXMdBe+EHR6L0wzbqjeabHTwV6UITJ3QQQIwb/ZhUaSwXxxQsbh8Mp
Tkx/OOuw6UgPztDqbd3bif4y8QhTNCmjChjVBxd/IAA3V6Rkw3bNGNbMDsk2JQ/AqyBnu8tQlJRL
TPcLXupp+RLZSHXef0msL85NePVdCuDS0vfktxCsB5EpNaXPbWx86Hs+8JTRXX+/GCKKZPAsRCo5
BMWczEFDZOY73WEp8H7DOurOMIKuYm30iu8gHvION56EUA7JdUxymnmYX65gTtCLy0t0LD8nJgFn
b1OHnAvTvB671bHOzeWqT882oJOqxYT3/A9hd8h79jShAyQRtOXtejzZ80S4IRHVsvgkZt2eDR8o
Ts4EX/9l7Hy3GDUilviumNnPwt0Kxun2nJKKv207EQx2L1KoXb+YAe7Q3GvVVDCY+ncW3D4StFeY
mO14hKiGkoaSV5AExWuGi5S1Iwi5pKeZlxTCBufWFpPrfqSQ2nzVQ6ggLfOzmaMtbVxC60+Rnt2E
dC3WnxrhYsraFw5LiKpQftBF8Z9q0CmvVSyCyUU6vrrmRIql1Q3yVYTI2Q50yyotpkPmRd6OK/iU
pYJ7+6zN5pL0DClSKIcLGlyYct7bRkenXccUQtwdc3jSlRw0sjO828ZqrPRYdt0+G5p4ISFLw06C
FpMTsfT3Q9W7eN/PSsSR0HpWT0IrnFgcjmcHt+BBO/nYnQ2uvdT/mKV5h/KYIBd4WjQSBzSqRPaA
Eq5UJW3oo8CPRG0ZCI8+7oNC3IBmKXyIJdPYeDyOVfhcXv++BrffezM1Z4GE1oZYkrTwnL3jgM5N
G9RrxsSimVD5KLx+Ynq779xnxLhPNTjgjS5z6WiIRgQv02+MCOp3+GPSxU41njiFlRh1so+LDAfw
3hyzUm7deZp0SFZIVbP7/IYKknV4VWbt6jcf9mXzVn0VkJiArFBTUjAqIa2FfXgeeBQf/KlfZZOE
2IS2iT8GBRi2Zhn0lp9yZA282/iscQNZVDZGl3MLJM3iFa8CO6Q8CF2bkvr9EEc6TUHCub+KXGPW
69NMaFW6YaLckoQmVbgncshe7RSAiVzipA1YmgaTo5/fvtxC3pU6g1CXaVVo84N8kmbkeoVYj6Zg
y14nJXpev670StkiEB+HtMq/lbwigVB3pTEyNVWk2Iu4Nv8z01MkxL5Alhi2F7l/QoE5KTRCwApU
6pEDT2Qo4P3ku9X2mwlYslXfVT9N4WBoeqSPjj9Ds9l08yo4h9iS3VRP2EiXrABgok+2QWjap25N
8eFRjjEoz5TzDAxzHuU+poNzFVDKl5Iam/bhUh51FBdMI+sc52lQ6EcnRuPfFjPe/GJKX1qisBtN
5rKsz35AzZvPswJ/umQIWVukh3RtoM7U1cgZ2ge/iftZYZ2tXXtAclRBXwbykHB6KkWOm51abu/x
sR52VwjitjELYS0KQyzweHjbqG5ZLg4i3hG7WJcTHQ/+HCzv7F8/bk0dd/vp1Wo7H7h06GtUB/O/
GTFDzMfra/uSpq79QfqPbrgBLRoWQ217i8hAeI19RHtghow1tbS8MUsJwtMRPIQsLS4SHVGT2scP
j5G2bOgDv0MCP9Cr5SbHlrcuIniEaGN8jhe9ffQZDTddVZCIaWmN4lEWQK24UaKrPth17Uzw1Xj6
+PzT9QCQ4DCMoyXbqy7eiaPIZ72lqp1pNWF7uykYb0eeD+KsQCgpWzm5k+KTvfWgIEHh4HDqt6Ck
waJ3LAdbw9o53222XZ9erbOCmjw9bFVSNBTDOvCULoTcRp/fJCJOEVMIy0GIUBBVyIHiEeE8eAe0
hAHY1BtURFo9DRWeE/YovVlZSSMcxF15jp1vMp13UF2hGugdlEb2NdQmIH1w26AVfXx6+dtuKyFa
7I+5vK8+9CYtwcfhYBkS1g3eSs5Vy4mGCdrGdpcNG+9aVC3mNel/0AUo9ai6Ab/ImtmJagy5p3z5
Tfu6EZ/NShiGuXiM5QxovlyqeAcDO5Eje4+fJ/RHxTesdAt5MrXP3kqTFMsTQOBk6F7R8gU+rHDm
7Zko0GKnmH19LmFuqgoPgcmK/1V4vJYSep4l4qXdAP/ldYZ12nu9OK/lDM+f2vTMAvmI8kgv6aLc
45MpbhnAQpvFbrKCWsb1sj/BXYA5klvN/SeM/HDMkVYtm4a9OlmTp2lwA5u3sNUD+dlYRlVM8Swa
BDgE2sN6+YNcKi6sw43lHhWECs0I7wBytad56xI89GA41C8m1oUGsq1JC0Rwk2tZP++umUUa/o9R
GrWp6ZLJPNWEqHWNyxU64NoQSfP7BYjWrlQ0m6ap0hdwOhwyunRSDw7VnTvm+nx3pZITkd6JECxJ
yd8O4fqPyIdnbKcDTiTb2K7eConjmWdVXLKqjii1ZHKwBbAyhsQM3gLvXzcLXFcaGI/OfAsRDx/9
5Oof7qnKUt/T/qZLeGcAhQ5GwxqksihEAeRYwcBN+/1Rq9JFKxC9dy0jQm/Eq27hHBL3l+GiQtrz
5F0J50b2aSBO0gF4uKN6+xvXJHia0+TyJak7iya/zxKYnSObsTvEhyTezwUJEMFkgwPzdRcpHwo0
Wo4k6Z1d8g4zMh9lv4Og9yzPs77E6pCQrOeZpO4sbX2b8fJCENQUkgTAt0YTLQXpXbHI5+wOOUQK
AOmhzexZZ4Iv0wMqvfD1qGCDlPcjGfFYJsKUVtY6FtnAFaqUosxAvG1mRMfLNWH3T4UaIwkxjdmc
isumk9uppOzdL01vyb2vrH/wDmHU8nP4HTaEykQDU0klGIlj19aCWgf+kOA0t60MlWlM9IJi7tIn
7dafXx6mFCMv2RE1sUOOt6UOIKVKjh7FnIGYImxNqAL1YDHgMZv+bBNu4fw0X8YteA2HxFn+LrNx
eqGwIhKaAnFFdTeZBISx62hw9I7C/e9ZwhA9lNRy0tw4SxXifj/U7x8RN3zR1b5/C3zbJpP8KTrr
/H7Ny1qq1h2fFVxhnArt4ZvkYb7cDpwYPkkcYqKP7W1B5otwvIOeys139AEfEU9GTkO/KXNQz0H8
RJKBMe+rNunI9exAt8Cfw/R2s7ihdgAVYnP2cHkUC2vt+Bf37moYbGbaGJ1MM6kseQjF4hgZ57p3
1fTKE/VveY5jQQk3vbbMUqe57KxDVhBlrQOACfzJ7cnXcBOas82nKshNTkgUvPXVQV7t+molljCq
dyLbfDB1tH38O2fLihjsvTJxRlJXdeG56cYzN7Rn1RiwQLRYx0gSN9ftrg3VtuMxSd8Ydw09CZCq
zj3V/Kj3502WfOpOHjoL9f94OJ7nRndc2+UCzSl8LYoPpGuHLrlhpeQDwxOGyKbF+dBRi4n6oavt
g8pxsp+sIhglZ0zawWbyMDNuE+NYeUrptMEPERuVjlD7YxEtqiQE7AxEkVMZsV/sutnZwhZD5dEg
rxsCIt9GPF2OIcMtM0htuxcLTroH9l3NdodF7QB9cmn5aH3tFkQvZoF1PM6SRiiPjKhFyleB+fgI
Y1lM1lmOuHE8J8H/7QMq03M3p8DLcLNP7xTkQJdTopwBkZP6vuEX61RCkySz+SRaNF89LArbvO/V
GyP8ReM96QeL7seIQFq72FLbVVwKF0Ust/MXVD4447gl+uaIP8wIdWZybk8gpSk7CFZF3mYoOBlM
PdEX5nMD68UEUFvyubcaNO/BXF5G63t92G8Y4RtaNLrmxO5ZQI3Ue3dqMFulkWps9dSAhrIeoHMw
fj06rGSjpVkP4aTt2kxqUvsC2rPRX+/xxrDyTG770IqtocNhY6iIgi2AQMvgc2v+K9ZdO8erDtVa
xWaKluREXiZ5Bm4rxuwX8WEiJBehPINFoLKQJyKOaLanPcBtcy/kGs939ByuQLAdWRa02QeM4BFp
lbl14fFsmduGcdHV4SV/7BBAVQHEpy9cBkq0R2BDouS5LsVZqfhPEUcFkHgfO5IlG41IXIDXEgu8
FmmZw7QreiV8CLT0NsaMtZgrJL3cmj+Mymo9vhYPYInIFjeVPCNvSh3A7PlA4JWH6/nGEmR/Gp8k
N1qR348clTJ1qeVUTFWahnWcS+StXk64tK4oNXGp057ROSDTlNgE3yTcQV+On9DXf0YfjDRDlh8S
AWF8kzU8MVHXSpG8S74Yz6YCpH8vQnPmn+OhrWAPmquesXQiQVtckdH1xoeWhkuvjxAH+MWj9XkS
itSYmnsecFDoEgFnD6gbTtV749BvfupHTUuIdtPwxWoSJXQbmRnhXM6t87Obp1uhJkrPSJZjjXYC
LlRzj7fHNNYiamIX4fnI4JucYS/u5nlGkwghknG9p0TEMO309UPHIevFzELJru/ayag8YZfyl/1V
KixMmtmqoEuxs97SF2BsA1b0TQ0XXM/o5xH5kIyJMlA8/iyAu/pw8l878ZWKw6sv9IPKCXOrsqvI
AfpZwe4BLp1WPeMHuFWn6t1NhXbfSIQ18w3+Kq83jzPOy+u2/EuJyYV9IqmgYAO1bmyrwpCYFjIE
SEF1oW/yOWcEIx/NU0NRylDDQTHDfUufn149BaBN451pM4AjTMLbkJTmMicVjrL83AGIzbfE7U3B
8tped2UEmi4NU99R0vretE54z/37vyX9mkDOb9oQ+O8Ny5zvJYIUqGLnCQeJRAySTREPl7UiWeXf
0dj/wIUKP2a6Albxc8GJr58tGzUVj9KKlBvcLiuSORRZNGBKRVzr2Xa6V90O2Dud8bvI0aiB01kK
/maV9HNmd64qlJgnV8YyeUhuXLmKX4curXjcNNMC03d+H9ph/Pg1niZKC0qk1Ut5sXQsfaxMSsfK
6rCyc0oX1nc/k/snS5kTbGBrKX7+qeB8/EXCHWmmDuMODBIcd8r4Dv+NdlJ14IRzN9zWrlZVeMr2
PwLPJiizSp9lyxAJfttLD7dWEXL709KYKJZ08fLt6Qs5jWwgM0HmGGJCapLpXeSFFrIU0+EWgfxb
YGOzU/X4KiEhNJ8WMd6K5HwlsL9d0bcy11Gs8fUdaDBqW0EGncZ8xg4HSgPfQmRySwiLZMsGBcRB
9ae/kNPXo03T86JQDNSXE0QTB0IgYHVDHmpfBgwAWN7/jamhF8Lfm1Rp02Nyv5RkZU8I6xTjNngL
cFCjxY6B/IuRXVzMDj5oxjbydFNfilKs6wqZ8luTzlxdWmG5ORBylqLM6eQaEU0qiF2MlZZ6ulNS
AW+urcDaVBGfBbaj0z6Mfnxv8nKPlKLmc2uKFo3dO6/3Tl89m63117bInuQCVYWSfsDnsmYKN/3w
nXoez0qjDtuvLYnuo5aGpf+DrTepsIg3HHNCmjVDmfLO2bQyLl8hsURMTqGVigtfE93eFiX1AdHj
C60vD9Ip122Vw8ZyDyFSqIcFtkePGrPnPsM1F+jPZkZsMat+hbsBE+jZhlFr2LaAYRasw3qBPHGw
MPYRrCmMCtw4fWun9yqNGw3s8PivvsmxSNhm+8eC6N+moWAg9nDXSro/a1sHSXyCtB9T5TSt5buy
OE1UuirJdltBzcZsrV0Pzpp58s3MTuQeaX2kQijYj5sAbiASwOCLgX75Lum+kIQ9jgotwMRg+Bm8
azh9SsLQvTpDG7zbhw0ht4OtLQrCMdxv9mh8Exl1bNrbAwb05PCUGIgHwBjKEt7ovZklxbPXygDV
9Tvb7A4k5ZXJbubyXI+ZoQv0RUBJcJVCEiNjALEXa1Fdhk+qfJ0FgJrbwNMbVRw0OVKZxcsnzdzE
HNZtA3IQ8l5zfFlPmMrmJ8wYDLOqhVSwDmZobt7FilHiDLl4NFQT+kdtPaHaLKQv+yGGnZvZdvXT
rio3mzPRghjJoUhRJ98ZCB9zk/wy8gyfXbkssBEVXn/98UpnhoeGkY8Uei+JKQ6RQSIZ1PfQQ2Lx
I4/1JX/SfbHTfj4UCoKHxz3yntWAnZ2q3Y5b63fosmXqM3+f/NKX2/nTd45AoPzsMUkOpyiMY2FJ
3xJ+M5KXd5rTXkHPaKV4Uy7gblD4x2eaN9X6ag9tNrgEY2QclInVE9M1tro0nYCLT+akF9E7CkxO
Iy5/rFNU/4/iTJB/8ZeV67S/7zbCtaIkeq0eFgTI1C09s12WYg9xKs/kMhSJJoi/5bL22t2EnQU3
+SuhlnqGc9g49FrMbuDX0QAE873IcVzbd3GZxQJy9J5ZSX5lUuJWwUyVCUp5DpVzyJmL5XjjX9GF
VQ+VenICg1hV/hqp56OUroDE7MKIh/vprGV/UUXtC1nud0JX2nJpcOuweR9Td8WWwKaMz2HUyFtB
/DFMHevrHGi6SUi8g4aVLAYcEYCcpo5BNkz6GbHM0Fa4Sn0DH/rwOIP8NSGWbhKVK1DlRF40dGIV
rPskbM3hcXnH5bpQyrcjgjWCkXAkqKyqTUttim2xch9IwJ6gnoP8QxufhGXgBDCOf0J66xBhFRuQ
2VMrlN2WON1+sLYW3mMn6874951j9vFteWEw3Vv+yYVH764pPyIvXzn2QgNJhTWPAC1uxO6Z9zYV
rKiIov7WbVTOni6TDfMqQ8KqXo1hg53kE91eDIhzi47wOCFy9Tu+FrvfLTOijszOhCWE0GnWRpwE
RZrJdYgjzBDeDcSoHEUhSw5XNSH6N9jLjBJKj0u5ijaVzkPqAyHWA/jhmQv3RVeIOFn3zxK9OuXS
RR+W4LePJVq4tNhI6wEOJdZr+uh0onjxDRzT7KPT4ODlljmI9iDjC2DdiYkNJ8RtgpnMirS3AF0l
u2MlY44YIxPPlWmYF65VItGKZ+KBN295+6Gxe6vFUUdpQa43w73sw4H/wl/Izph8051NJxgsBK/C
2xyAmYi7d5HKcfmb0mZxf9ZY/bR6i84WM8xsWeTfrVow7DLhGUDLA53nKv/PvKK5DwQ8EvN38A3E
nbgyx3Rdd3b41CvjZDALGXr0tjjlEgXkJe84pADtd6IVg8E5gegq86MvqwWBAtydVPgB4+VKCRxA
SbZ5wF8k5t6qcwbtQmC/fps8cFR4lVqvIMG51e5zm84JfsZMmG+zYz8tS4hUUQIrApKDtVr5dWGf
kTR5yg2hg8RIduuV9JBffC4ddHtBHBVkBAj8y/BCjmdP6Ej/zKq1giBx0HpPPSyUmcmvlUwYrCXj
0LhrS2YV61vuieCWmvBCILKeFYbva4JGSWJv+/h0ktVDJ1tqIygLHnTEkbLGSH1/QTz9c5X+daCk
ZcmMf9V2TdA+BcKtU9bJj9rYyHkZgV7dP80ZHxgc7pAEJ1Ynn9+UaatzD8pIAHA9QONLZuWQb7aZ
5iNYiz6Q3q2w6eQWG/CGndlyHJwpwlzl11UJN4wSmxO1TOF74H30OJ1glI+gS0Kw//TLDWTDOFhO
ARNh0OrUZk/5Sg5y6jiHUjwzVC0zdhZz0F3YouVJrIdt9klbwqwwfbjGaAAKkpxMpFydMz1N728f
7IL1t35tnf8TfxoGzQ4kUvN5IF5QXYJtGlavbyHSk90zv8y/pDlitv0u6jS6FEqdywGHRhn7u6vs
LPOmXCUnexdAMs/wC3wAT+PAhcZUiP+QEE9bdq4N8FDh9nHUDIw60a5T3byxSVknW/mWoBYrGKCz
is3OlkKeVrDlBO2K+ohS3e92kuLz749jvTbmJ/Zu8pmbCoAyIsJR9q3sfxHaKN+A097cXX4yQt9h
ddoFUwKKyyQhP3tJxMdr8/RpxS/85UD6etbPCgI5xN5RJbddy366D8MLHHeSHoMz6jKm9BZ7Y7o2
VuXvEaLnYcdec4uQpazw17xvn3IgeWPqWyZXyENZAUi2uAHfbfOR20Q+XCa+wWT6LbXMbinJOGTH
t5uWN3+ddoRzPiV2d1NmBnTsBQB70T4dr1dGFZNgzC08aMe8rQ1dMFW6+8Y1PzsF3LtgTaiXQiv/
w4+SEVmDUzbG6kZe9uWSXN2I7jM0cdLNs9RZ1WL6/cxZJnXGGP733cPXXS06g/6F1ESEDorPmQJC
5n9SINvcFHCI4/lC5kF+X4g7xHVoLjWsK/hPgKW/q4ABVtcr5as0nVZDbYnBGUHWQpjz2KgINMAE
5EcfVWfTFxYrcHxDv3p12NMPjbl6+KmQy+7q12UwY9PYnqN1m8s/tb3VmqQvTuwhf6ANNwjKc7j+
qk26RYv7R5j5Plp8c4ClLUPyd9RwPKU+8MWa+bnZvKoxUYltdPT98AqT/dOTX6ldSBWg7ctaELre
6bsHI6LTIQBW+BOF9+JUu9K2PnPqjVP2M4liQU4T0qMO82WTEI5KILLSp2lerEw0dPG9/ZgyRpgB
Q1jlnFqZD/yL3Pva2fkvIVMddEsNQhxsdceOIcIooXmXr6SgFSGJ+PUCjk5R7MoC9bJUfCmFzrdx
jhT2opun/dCphB1grH0sM7g377+kjpfv6iUPKy1rbS2uT2idUwJjT5X4ahkfvIDQSNw3kplPqLV4
0fPsLSbX9t2lWdvIFjd6ydtL3sVe0hrx6+77F87L+PnbErPZ+2i3BJK0NznKQIldIg03W8B8V7l3
zLdK4uIYn248/Rl5O+QLiYEkvVEaYWvsXjhTJTOizfyosAc0wF8N/jWJsGnKdoihi/csV02NIH3k
EwYkFxxr1TndoQRxK3A0Zbgs8hfNSa1YKB0e0IUe18NNyB1WiZtXdq35mETUc+J/ZSowCruUHE8o
+9L5nL0W2lsbLC5mIc0JWGJbmu0STCrvHwn9IQGVw91dk6ecUk/XGNAnf65Qst8JfrqxH+HLwul7
zBruJVMbdxnV21q9nltmyoWfgUf0iwcVj2b3c3gB6d3selak8/MS/wpObxQsg7+Ds52SxcPWn+C+
xoUP+YpnYBmM9apKYw3p4dFy9KpKZQkQrRDe9FthQXMg6utvNEK1jscHBKtszpIcAG6CK/9DtsKR
MTk0lRbnFY2Rak9WwSnzvK+5mjmxAhBYiovHkeQP8y6yQoWVX9PaBlOi8v2+B4kI/p7FRTDFOQ4L
3DHyZMG9/Oe6GG47G46F1MHoitAoSGptnrCTFCGjNPPmttdJd9h3v41PfukpuPpGmKoU3Wfwdp8z
mGeXeGa4mIIWh7v112sg8Pue2Qe24O9VkmI0FthhR08Sc6DVO9+0ufrHTS6k/+htByGQmr046UmE
2EAVR/ga5fdC1YjFYENIg59MsoCN3wveHn5YAbhfS+WY6IGlRm0B3TUcdbxzDvcn9N962mhwT3dR
en1P++qPAkw3VLiZjWHm9T/fdPncj8cvH+kI9S2YxuX6LYv5VclwGhqndh2umMQH1/InQbMG269I
X+pQnaFitlaj9wFoXcViDKpnruKEU+BsSvdgo4gi6rjor/LfkYVqSlghtyOKD/pkhTkYzBMQ8ckQ
iZjUdahKb1kG4fbyPn7Pb/I6ccgx8x3R7WVH180Vj6ABrPLHD/c3WHOV9kjasWrMBoY6u++ClsXX
80kmGd7tUhLZhOi82sF2Jh9qN67kZN69Y8OcBQGykWTLN4Ck8w/iqWVF1A27JROsj54u1yaNEBIa
L0Yrvjw62PM51kEHggnlw4XTLvzQwlRZduFaH0UnC84ZVSttIbhCK/AXg1Ck8a/9c612vsMjHsgt
YPfQLPe1PUlREMQX7/zmg9qnbyck/vwS1HeSmlBd+cyfrX2m+H2LM9GQ4PZfWLPAnh5LFpyNwwC6
k7RzcTNVSWIpL5XHTYhCP5Rmc4B57u11ci0mrOiqh1LkJyE8itW8YpPBlhKAShVzMW6/PCGS8IOf
1gN80B5DXvW98T+DyakRqF51ZuND8ytObmkqyFHo3RFbLpNbIuMW+qZaRUJYIUKEGLqX4t9FPLOA
J/0wQJWtHEinjBCR0ZvJd4Fj/v0/NjZQb6bNOLONJzpfVWjw8fLBiHSyHFbqj0NtatctcD9HiYAi
7gGCv0KQ/jasaWl/QbwxqV7mqjAmYYAbaouEWj1D1hXBOqtIO16vLjPy/SVitRuWss9trv/wxuVR
pAtTuHh9TdO1kElj8ax4ZGkCN3BPyMoeBk6OAtU7qWzXl/cJwJjQr0J27AKnAKes+uxguasBR097
JgywBVUGcrkwpwuudI/LIbcQWwjLhZZ8YXUToc7tUdMNbXqCyoCSySKnn/5hwYVAq9vYpDyIURmd
tAX8lRwi4hrMJzWjX3LleewgYqw7VyWG10FdJ/1Lo7lRn20+s/oBLfzVAMnWxnlNUJkrU/4YOXBa
gJrh4WdUWJt56VTkGsXiyYypxaAlO3xCmwWPO0j4C7Q7byGEmj9goZgBxrerx4kYZ89wGe4Q6Y2+
L29aaQ0T16wni8P3VSb95tvRNZRq8oTZQ/0U9Fn6nbL2mGzn38t0LMclIp+UoloABpV2/qvkPSLj
yYixfg12MamTVWaemxy1VoVRqt8aiAN5obeIxC1t7AHvt61GUS0VR1Qnik0n5Hfgv+05vBU6Ym8J
VLKqKKY8XjZ1hGW60b/0i5IpFbp3/1qfeYdC9l35VH221+sReVEJ8abPZsB3MNwxA9vcadu1xs/K
bwqmCk2CuZCHMoNhe+E5OwSr1Muy0ZexxAEFghv7LFzhfE6JnRu4A2SsUpzsoz35OFsrOYhVQGKk
lnBXGJXpoXy4It93qOM8ExBjJwowSg5yA2fnOQUwesax3TFP6TYkM/UEJOX7QRT1yZlqCx3cPLfq
/2A8ySnkRrRhDqBtorw7wsod2hvZ3O02wVRjByCEeMiiOxBIWnqteKt4tleabA6aPuDVQzv7umFt
Y17nn51AnkmKZktEzsfyBZ/NLSlKGIgydo395VFC9JEqw6YyVaBWDSy6PbVg1+8m3tXyF5RxzcKJ
6a7f9ze3KIcW4Pxh0Zeyfhc4ZtfwuOhE6rB1bcukDc1gfT5+SnTE9W9cDQn4uq2xov2mN9KQBGI2
5xJOtlRYljJyGZGZHby++EujvGPabo+6uPWqQx25+c7Qdg2OYbyvPo/TNJ+K9HJ5JaeBdcp+9Ri3
c3h56ge0QAfSVAyc6oTDXlpYbbH+0BiShfgjuSbC5GQ4oD68DnH3pdn7C4h1LocQftOI+K/DjQbJ
22E6UxXwx7YS8tIW9BEisD4UZB3YxUcyrHXw3WjSHspoViH7dgiAMUXdyZtzEIGZF1rsRamsb8iq
RVUZkeHjUaIpGpbjoU2IFMa9vKPu2mKL5xQI5R8BPOQPt9xT3rcdJVwcHDhDQLtftGzPh6UZj4SY
s2V9iChFkahNvn7ms+hhEjnYkpeKXFQEbR+DBK16esEaz0uiTTjfH1W0HM/filtPEdTtpeP4NQaj
k2VtHZp9Efgd/q9NOUdjo+AC38VF1r1XnYHVoQTcNB+m7X3Z2XXyFTTGLn7mTnnbFitBXR0Zo7vs
jpyYTZIrbLPqpUANmC+WPBeSBwac/kCbgSup8Mq3dpOz5J1iqJbjHRuGfb649JmBFx5CaIg84ns+
liyTonEdofUadEkyhQ18dKpdYSWhiYVog2zw1xjdbDCaOzAMdfPyE49s6iy3HgkBqlKM+3C3XFC9
nyeBOxC+dggS90UEYjjZ5aUqlKS9WVGreKUTtCYiGzoJ/8pKgXtHrXMK++eEOvxeq8P+siNNxvKL
SZmGTzTABj0S2gNmNaAp2e8e+MBzxEoOdbgGZYp53+n/Dmb35cIFBAhsocbTKKD1Gx3Gw3ylI7p5
Vd78asRbCWw/+2Kp7DN/6b+kRM8Pg/O6h9kA0gU9X4t5vvnMVbBmuvqzDUYkalvbjFcOy44A2x38
g8WzuBjdUaGeNR/zBpXuU1awd64prYmmt/gq0PBjvo4hkQj6CqskSOr+7KLwWmMlodLqMSSTfDxb
wWY/7Vi47NhTTpbYcht8Tehd4oYezmsk1HZyXBw/k5b4kOvcM4W6VteJoqhJK1UIJ38RyqEUsHC1
NrNQZg43Kkert/PVWLGvGi5Zu0h0q7Sp7CN+ZULM0nhl1k9tS5IZwGm8FnHLOgNIFEqoGqCvCt58
g9TzjtWHPtW48mbYqnynjMICDa1DnBu9gCqUN20d679nnhtkN5dlAQ5F5Ns+qn9opn/ZFM75gP9G
UMEs8IeToCQK+M5pb5LgJHKL5FIvAAQjmJ1UrfzYbAXgSHrHj2lilwuTwr4tzIlP2xkFDH2whVkH
oYOfc8TeN6nDTIi8VZkKWJdCHXPeigpfcWLrrCDtlGGNHN3/chG4AxV/CptausyG3VsFvn4rhv/K
ltninN4cZJUGPszpub2nxp2x5d17Rg+1uXdhdg2YRdAWKZJmXjLUbeYBXmGSRmTrLPZuUMIwQg0L
wr3e7VHTZNXoIOhqfnGtjWu4uWj22PGKBYSgFrjCDrh5LsEOrQfgT4tTFeHa+dd5TTjzHfGhasrS
QRXm/45sQGENQwMPXyqGP1+56DtLOfoWDT7DSn7mDIVRd61UGO43LEoa2yf/hp20qYYbwhaZGu8E
QXK9RDsY7DrFPaamDRvR8Chy16YRhNr/qgHT/BoRXtQuHMfBg0bjhMquCxQ8AQ6MICk6w9LhDyuM
aydY4cA2ooiKL7257TiWHu0qkjRjJwriqOjj24iIhPrhnXY36Gv3hshvu/UEVrc9lgW+V64q8Sjm
t0Pcb7/HRHkX/uHB1/LC1a8wQy9u0S4nlrhTYHrf56CLLzftjCKx1TtIcxvsZhl3k8uEEa9hbPHa
Z/Ov02Riwl++RZC0eN/vTJxVR79HWWYZFyS90Vw86iWYNQy0Ln69W3aNFz3jWvkCE/Jv1ghUlwcM
SZycEw96eiL/LtBzxK2O6mEHW/V/vKopwn7KCFYevTWtlXQLLq+dFsvdLJ4lglap8nx6MwIVDWE0
HuoHxTo9yMW2q+THkArho/1X+6XEvd10a5tldnaZOGlN5vISwhpm6Q3f1a1Szs9Aw2/nyXa5602K
0eLPAlphhy6dmLlkROxOj0mQCb3lAOs6ES0TsBXgtFswo4VsA7emPYV0CyDiMt8cOuRd5Gb41R0i
rHAJNJpZL/sPPJ6PVuVz/+38RCsBPonrI/gjgRDIf+Akz5sWS0qKiJaLpGsQ8k2nuO8ivHBzJ9eY
eunCXmQv0BOeIBCfV0uErI8Gl0U8XX2KtoKACSkivnkdwAXc03uqlucFpxWLenzbv1Zr+5ne36Ay
mJ8OtTvZ2LaCGpZqnaF3HbGze375ChaczRu5bFLboqDaVZ8z+cOcPBXDuh1oEE6SEKSoihqZbMLD
HBxQXQCBraEdGZiFRMGISTX/ApdctL5RoxcCbLsyQcsWDAwp0KdMiUYJ+ZdgAiL15fo43m4foMX1
GB1wS4GnxpI8k0JmcMZ7VKqaexk5l6DE7baXwblX3HtQydqwQaQ5sRFWzl/mJp76YtFfkqmE2aMK
SuNxQMC7ltnb4eAefsODi3I9jH5GII6t6/9zB/YtFtJnGg1HrvHnNrdoNQ4TVXNINwuZ2Yf2sW8m
A06+n/frfa3VtX5FTOUr91VZvRgEEijBSOy8/Hl1BjvJ2KzitOjNbNfaubvILcL8bSL06LukviQ4
JGcsfPQ28wj/2vUPxEyTgi1/zgqeX8tKT9DxKT6uQgozygxYIVl6Bj2p++KDP75jAwM3RLXVZ9gX
Z6AnlAAEMv9dZSsPaFjz+yfjSnxbsFKRkwLz0Gt66Z7wvKxifqKMswUD3Smro0ejpu535tk93YDi
m8hpDtC2QmVIRXZVfQa4SflQk/TEFDE/HOvN5wJPxzJy1L9ng2Mj3Hhmn2YylGtCaAfUCI8azdc8
zVZ9M4kGKunymnxVs3UGE5swln4Fj1shDAqMhKftMweQH8SVKrnqX3O3GohpnSrccrJmYOMng2oX
xQ6YB/2ckpWsTb20a+SqxPEznKDzE4TXbAu+WCEXGYub9LjfLg/b0Kt+7h4LgeeqOS/flaYapi7Y
JbuXeG0zydxcI3rcjIfrgutUa84RDNeSR8ykFQKG1569Ce6HmcYPnd5j/Ah8mj3qkPrx4D9itqKb
v86aV2Sqw16Qw4NXnJEzl9rKmK5arZbnhp8clyGFWLiTiMkpH4eQiOxeHFlRGkATw9nschQolFW8
6Vd31qNk2FHC6FXTHxoCb29Of3ln20QhZ3KIvNRBUfv0Imgj203jIzTUA7GoDVBRg3L6wwbEVRYj
ykbfVzvxDZLgiqJJWKfd5xFkQnJZrfU9phRzziB9gsHT9XIQN5QU1Xhb09CyxKlREJok50f87+IJ
oq4SeSQS3orx6yWQrUsINT4nu+tgB+AahfzvQKp03jmm9nrt8LxEnGgOxSkeRLmgB9Ntz20gL3Mi
Qoq/A75151TJdutRStixUSo+KmJVKIWr28CgoSJbjlbKIx25ClGTgTbQ6vZdhGfWLckgFQit74y/
NeXdzcMKKnvh0+OXxGyVdQLUZpAE3JgmrNm2h2uf+t/bWDDmCnhXBmf9pFBsG0HR3pVPY5a4m6ic
CYKcIMQtRPkT+g0WKw30+ZkHQ3wv+T795JLn/AUErLuZZgPP6M33eZx3b8nk94i9ggd54p1n03NC
Gz3Tzl8QZ6QEfGpsnNbdo9sZhQo1vnVsQZdYQSYc+xpk/BPta/5fRAgtdou0Klff5TYGZPEbn+iO
KXLbnnY6WLqCtjX3ehNETg3G8lMS2itTSy7KFlRES0xFQBkAcZNt05w4q2WMlu23Umg+xhg+zRhY
wSqxe+sBtrxPpEZosSnH/Wuz46pVG96QVW95Fpf/wbki6oPFYZAwCtOK9fobRfazo01yFD7678kG
f46NcDmvaXENJQnn7kaKMz4BJhaxvKmpCo2XNFNUkWRlU4KCddQxJ4rCPUe9DEGLsJSEOytq3vHz
YRCgg5RgoRcAiERRYQivdDo43Dj2cJ2L89LvMP7nvOs1EG9sp3K4KX/FYei99B9wtVe4T+E7PXfb
oj7+7oAp5CgFD1uGX8jyrlkbVj6YzHxXpY56XgMub6vaBlRIf0ks/CIfk5lqfku+9TuK+h8aITMV
7KbSZNlh/8UVYJzpltCIk2yP4Y9tSA8qfKjlIjTqKuYbs1YK3yOylDgEk/X/VPqrfWJt2QeiyynV
Cx6b/TPC1dRv4r2ne63tfRT4MWr3vTRpKKj/raNQasNxdoD/f+cKjqZb6LA74Van+iW6UJkSXZB2
DprWma5s1CC9YoHRgWTgfVupRQ+F5lgOT9qLTVf9u0QE2j7PXauh8cdAFdwrz4Wkjfr2QIh6Jf/w
R0Uqy3e6QCLflmZl48W2KvxDYpGmNP7GN/KyAdcU3AjLCiJYgPyvCebPXajJ1B73PowbUBdd4Nxh
m7U6C1JyQS1zhUAcSY7Chkd4ysHJooXrXvDgTeoBZyBiC5nIjjTvjBI1Uzd1FBTDBSiRs+yrpBFo
n024Fq+TMEx+crzMJzy4N4Lht14HeNr6rPDWI1UIpsKl7gaCONicU254tShBB6DnLnmuaN7XU+ju
/jY+cGaPETHQ/+uwnySh2fxhv0oXmR1/3VkQnhFBa7dXF3RJD8OnFs6yttYWadKaRupdvZc422q2
SoMwbAqtoeUdzyZ4Dnip/aJ+IZkDphhwKWvsMqPFTWsHQetl2BqaN2Rd/dgIppjJms99J2FcWTyh
LvwFMfbKBvXtGeQ9fEB/838nmkHTyztpDqkhDe0kvDvp/9M+cc8E3opZ8QIt2oxLinRrE4B54Q24
MX6fC8oRluoLP1d7lObOS0AVnPrbYjjpat2d4LuGjYOaWDd4B8i/Tjk921P3Gam3otebkp42rQUo
D+IU/CIIiu9uBRRld3oJkkT58bhPNGlQJKalCI+sV+IurChsXy8XequxZTiyPYd0JE5m0rJNitbA
U3PmGpEN/0CczXoU7qMo3iWNCnSCANXCU5jBNR3Ly32rHTz2NbWp1XxJvztJyz1gNHsPlA6wVRo0
dKws2sa1SxTTZ+5wTaeb99I2x8u1VxMntCPuFh/4zV3tS3VdxirtFzq3v5awS7bvsbkfrvcoT4EL
UgmEn787vRHkqdbZSO+Ougu24V/9mtSq3gGuY8/xqbdFShNyQED/5Zx1eHP2+L/6SwvKOvUQHin9
Q++UOj7IV2nJ/StuwSYRbWtSAY+G31VD34I4vcpD5Cnda/ygDbkNch0NZoYOzUYX8I8ryCn6UzX8
abKyISajSlqhv6w0jODAO6JvHni7gVXXVFxT/XqIToDTCB53NRxIaPl1uS3zLuBbVE/23BL6oNcS
rrBEkeoo6xdLeZ66O19ISmxDQ/1oAPFOL+OWTSPsjDa/CNr2pXaz0djIhlKY6AHigd1NsykXPahO
Lw3oxVczeddYCos619R2QOszN6gmnvniHb+QMjK9jv907zUCINxR4vYzI+VovcA6V+ogQJVXrNbh
xRUnlvcsXP94ZHRVNy8IIBQN8DxwbT6ccAJJ3ndeRnIzP6Q/GWQ5KSAwrXREaF8ngp7GLw5oIb+e
8hAEGznHuZA9vcAqD47Zv0T419zrutsaDvtYXL0MSELi/N6GRKs7tJcI42QDiH4KC2c3zrzFDScH
aJaqm2MtuQ6UKTYYHY2U+306N/dQXNdHCo5OenbPJMe0TpggnAvcZPaLypmBqeVkM30oMHiFEph3
f3IHpjmijL6SYVefqcWKW2+TRe+QHngvg1SSts5ZzI0cFZZGx8WJmd7Aj4KcvdCZbkGwPmegGRck
7JdXn0AI9HnFuCbhDtUUFY+wrCLA42AlA1c6nKZinkwIfGEfw62VR86FZOJewXzjTQORKSqHxkkS
wShjReq3ibXstme9CZMrvk/FLr0nxp98YxaB5kmEFlm5T+zST0ZzQDfspUyFh5wQoeTaonOdjyza
bx5trPFzLBYuj5HAFaqJ1VIT2WhFK+F/CgLZpqvVrpZnETJ8BPcZ9GDChzc5ufeJ39GzcBvYSwba
/flb9MZtGAFBiZphxfUdTNl1A01IIL0JP/P8qrf+GZLH71eklqqusk/QLWbon7/X3h3iEElR0iJ1
IG11k/vJmYT/fNfLZW0i/CwFX38t4X52dmnPXl4YJcbb3uY+Uo1s4mLnZOA0pNDe87Jap9ZpkFco
qK+8nxO7R3yjW0cEP0VdqBGLdS/p7E0yLx+toIz9/MyMa8SARg/fNC/XIj2a7oNtI1NdN3I4HNcn
aMuCirbjqqNgBZSJLqwGtzHI2a9NNWa/6RfCZveeutRgKAOTTxfN/1cOrz3BKrCSGcNowRmJzRkM
eF7qew2kr+bO9Zc2bfAjWT3DLbp2q6j7g8om3wAjAGP7Ruof2QpSWjtYrQCZcKYaEeVqN1yjsA59
u0YpeF3ZY8r4rAQHLBM8fDp1HFDWIufaZw4VWBDwZD521f8a9OyOlij+KKwuc1Hitb4jsUu6TI3b
4pnC/eaGZknPm6PqjlVDgXY2Cz2FOlfkgIAfyOFstfIOT0kI7vZ7gZX2qdPAKf3zZ9JU8WDKY5kK
GJDrtF9FlKuxnxcjeknPemSlpX3yimYGtCfWmr60uRbVhPpjMvY6iNyhs06XA+YR7U06fsMBJC2a
dnmOsGg3P7aksfaDms8KTFnTMy3JcZ1CHe2PGq49ajVMiaGDTu4F0WXhvyUcqbiBsJpvo1dWYepH
3mCI359iB0xgsC0gGQvGhpCKjNdplaLO06Ts0ep8dHK91l/yCr4XnZvbtrr/mCu1g7zQEin+5bZc
ggrVTv6LOPFl0pN+jasw7o0FIDfcpukGAZ63HANmBL1y4wodJ+XQ3wM3llicXqebB9xGMHtDPZKB
IYp3zEMiPgErgibrfYZKrhGsMvqlHV0RtFbQha1aPiMrbUsjluOYq8PN/1HKuov9ut+Qc/Bk8OR/
Q/sTdI3wG4pAhZVXlV1GZUtYfIqs1yyjVO+bjMY/BDplR03OMIR9ulNKkqNrQ+H/visGwCzAjnlR
W7k917hU5Mv1Fpa+mT0s01DPVoTCbwmwWm8cvf2fIoYQtuQqax+g6oJ02cU9zEzGKGY8IJKdSOF6
yeb0A/PzY6Zf6liHnUXMHKC0LrKiehv3zDn7u+yNrAJ36nuLqxc7jL2/tvJVEziUHQEiBCWBIqBi
Gb7CiUA4UYcXHtzeg3OprVPfK7ZVEEasdgS5KG72SX6O/HvOc4qQYO943cM6j08Vl9nmymGYn2bA
Fi7zShwJuMj4Mt7wTe3Dw4aIDogd+yDIAkgBrcpOAFnAS6KUu6iNDUNGHXciwPqYLJNdfX2iJYge
a0RQV9g5ghL7oesZTU5Gg69B2XaIsV4OfL65Kafqr3fj43g8V/gPtV5iuIEDEi1AoAHe5MEaDK3W
hLYAmue7D5RqNMeSf3QZ38KcKdHOkMdo9MjV9CLjQKythB83snPl3+zH4EVun0J1toaIRy7l/Eu0
rkA8LJo3MJ8/9BmfQyTq347rnnEWacUwWwcaCHUIf9oEjo3IpnPdwDbViDBN9qQlKD5QPb3vdkBW
RIPGxxzuXRVV4RzbWx/Lngwa37dsDU3H3Y4rDZtRvb0ve+hztmQexUFROTVNOmzzIqnUBDvf3cWS
h7jt+rjmT4ghjhDxQqq5mMQyf1Z/ja0WPeC3GtsVlF5jpfoxNrh4k3d2ZGJ/TMQtUh9ApDZp9z11
y8SewfZpotNpfjj5smWZhZtmbbi7vELwCjRj+7R+huiOs37ypnoQsRYH41YiDy3/K1mmFbTUC8Ed
FXQN+BuIqLAPJCOqeYZfg6HH0ITZ/FVc/pF9CxSQMK4+jOAtVypyB0mC8+tUar09exAGbNVT/3FD
rcmJcjzHptzGm5RLPqvkFstssroRj2MzH6QXZMIg+YChut4/94ikujP9pMkn/azXpaliJpVWoFZ9
xheQcatBYXc1VDcwJckjHA1KFuMl66k7eIDgcP8y5KdEGDC5vEJbxAbRukc9Cq5zPhqH8aD8C6B4
GopS+lCPy7/yKXZPTMdAyfEY2hgVA1ykcAP767K2ZiL4KVxgfy52hIyxBvMgA937Mo8NuESDQ6n9
gteR+Bk7+VKWsCI27Y5QQpPDOIurdz9tQrYwzvkBH6ba8dhyeVebch/UoSAHNwNWoii4LEYdkZdJ
SU0KuGKQNYIIbZ+E4anxoM6Dh9YjSQKwox/L8weXCOdG+tlSXSqepifTsYujAtCcne44vHBLuK34
QxN8MTZRScFR3yVGAG5JtzEkvxMmL6OV6yTfy3o6At5JzbUXQDYl+5JZEVu+KRYYby5vEjfl8kcw
+cxTBjUO5rLlONHcWng8ZRa1+1wbQsfUCJ/w0pNkwP/+GYHMHLTQyYxwvG3zWR3vlUkH3VydX6Im
RRNvH421a30f03UDJUTDq86ibr9DnBiiA/D2RNrXDrSOtcTioc9EhVjhckuQaR4r+IXIIDW9atW+
QPyE3ALeA1EiRCpm8QLhJ0+SM3D1+FQMQLUa4TP0jpPdJ5Kli3cJgYDvXdBhpa6+tQLvPnoU3OdG
HLgZxo8yeugHaO0VRPYnEFO9YBUYeYmiClUrZMElayHXRQiIljJA30cqzorH/s+MBm4Qy2oGlqub
M8stcs0xyz3Tt2m/WPjITw60rJHpwUf6SfBqaaNzXoA00IoWA7cKY6b9ltWvPOrokf6bfZ8FpRQ7
Ir7+Bs517UIt/RnxuL31zOalKcPFYQsqy9nWPUzbtSc/kmx11s8BT83dG3XBKAmOyLxwlfeK/nWn
MPz9/Rc9XChOZ4WrcXOAAMmhrb39/cJzQq2mBqdaUMk3UkLclu914IgiSrVaWp9glH7SAOWngMRD
usP2NLAPyLmxuZiqNP+NHU8WqTWJKh0bp1m0pj84U+kgFqjTbgj3zfAiiiIXX/6SqzPxn+AJCgFw
jr0TKDyPjGvtH0h5T5JxI0n7C72fHplNOaoUgceYbAqTomMzFa9dv686ToiFAModxmYI7Fs9H0rH
Tm78uUwNzYDTfKCX8dFPmPqKSURBV+tzQkd9RnKm7LUD3uQHh7cg6CcWrarP+FhFEUq1Jzxu3Gb0
+dnZxjIvOfahgGZnhxsS0moSlnPo98nQ8FW6FkaZeAmG6Hq0Hb3is3HtdB3rBwoKFzu1md89e31k
WU20R2r1M6AN1u9Nqh1/mfCP1w1SucveGPJ2+V3H4Te4vkdWd3GgANm/wxVfCwxK2ZSMquA0Q1Pt
7NeOZx39n2he1xa9EuiDtgKYWlxCpVNn0R2Nc/wVgO/+kxcJo323En9fw6At4zvq3mxljehHpegk
jtPRU9dC4LdbUpfUEurDHbaL2mN0H+9Uy/pDFRVjlQOOwbLuH7iCShhqIrgMI9Ikfjd4TqCQ5yQS
aN+S0TiWee0gGatAs6emv1DDEMuta02X4AUhuqh8JDhnvyJPDGm/bqkmB2DVmYJRAiDPhlzXXhu+
Bk36b2auPPm8JfQ8R+9VuZT6jVzZZIKQ/mgsjpUXJAAaIWo1MzxfGUYYXJpSi7v9+V0WLX2Ukf/H
ADk/+30eBfNUVpDKHvtfc1lyyZ2F6ka3IyI8ixhRlpQnc6cpQLr1I2gC1pTdDO8+D/zorPsN+x31
VIA1gTHR2Ue5H9dWUxOzBfsl7rhWWfmUx1uQKOZ764LaGMi1fP95+jHDaGk0sCQ400uqbW7hi6PZ
fYPhb0XOCZfkMA0py2xxlLEEpqqqxSFnKGj3nyNT7nWDexVq406HbBDIpj3r6fW97FyGGonYfe98
TVH0og/xZtn0M65wmnYImK9Y/UZ3IYC6u1ER8u3zHDjfDYAQZVO2jYUkHdndfsWl5f9xtjm7aVwk
Y/vtNHt1JIrrRPXUb9K+MSsSzYN+ZV/nyt2bfC78r+GZMIGhMd0vltBzHdrzs1FYxMGzdXCjn+qX
fMwGsD9CduqJrGMIXofVD+jI5JUkW01mr4437A8y8+nwZqnODJL24A5UY9bzGJYyh/F5QvnMClh/
hffB7TerU+UsNP2mH4N40QRxbYZQCO/YNySamG8QH2qBTEoM1NkGI4Rn3k4kLAhUC7V7Bm+9Wla6
+rSxP61QhxHF/+mWGZtZNoqNm2yabx0a+kIDxi3RWhJOJXNd5c3rji2G6Q0tvVdUj2TV9JCV+Y8K
XheEWvTJ+DPHc0yGycWBjXTGmjN820LkvXRG4RjJAG3cylTQ7gr8cmQ75cMMMckLx/T+AkchHrxD
RCWKc5JbSbG5Exr04UponaG9JJysvW1GkrLf1hV/QznZzFTdtK2tBRaSrRVd2/dIfy1q8ygdAVJM
rxA58x90in6AVO3xggwl4PjGYlhL+4OkBL6ocMT2slSNyVe5OFMN6xMfH9bEGe4QTyAvUSqhZMqK
xEefPexiiTCpnyVr5OM7jnPuqi9smMhVUnNYs+DoIwVGg8fvSJct40pEdA4oMzJ+MadPvwKtZDJG
5uZKadx9bq7FA92vQsQ2cUJSt37xproiK2MSb3+0iQ5jBagMrq/a/qpPQ8pxjuMdvsn6Yu1r34Wj
5wj1x1jvpPwBpkksEwk/OJqfkF2tS1OaY8ZL3meGPxV50Lgl8smb1h+2usdRL1bJRSISDK6vgbSg
FRE1GfRBydhAjPaM5WYrA0sa3UGKiGGVvBCBreggEXvNLMVBuyCo5E9WkQYdS55yUjSxbd7AWseC
l2AMb4NPTmFJwtn3QoHBzULIOlbkGaxqK1u94/I1J8AOQG1sYU3RVIctbJabLNfAmok8JzQqVmcO
P62VsSq29NMK7M0nTctsTKEUG7xlExET/XFy5ZnNHdkxbyloqoHhyI/3lkp57IBI/hIL0KkDA+Dx
5qNodvq6EFNfY7Ne6P+GQDovUHvKVQrRTj7hC4m5slYEFKj8ML5hawr8OF6snl9/bBFrr8tpMbZz
PaDWlBDQfsDBNtNfMidUcfNiCrmoEn9XWC28zN6781LX++5drLiFzMoq15MY8lSuqq6jrVgaBJBu
0ny9AdUO4yqYUP+Oc/QFoe7r5CVdvsiMhjJ6TQ3Nwmy211thXauWnfruK5IxkrlmRaPd8sYW4VN5
iUTMi5uq9usgeUFz4DdSXRRXKlVzqrrWt7xLEW1ziS37/HxSWuwNiRiQUk4ada2o935eZd/A//mf
sl8bPwWiT3XdwuQzB/+nc3Tc+KKweJXHAh9D42f/BejZH8O8YXpwCWhPmYaTKuCy+A6hvmOh8BpJ
IkHcW/5huM+twlShsnsmgnps9LEwgJDOd5Ojoo+zxebKtyO+Dng8GFBOOhsW2xI/DqiTuq72bo7Y
6NLqYmyUTuxlUdiabkCyLtY3YGaVwgfVLrI1aCP/al944rm00PiBbjUmHpZG0tPYB+jxJL/UW6Iq
xvi6smTuA0MdqUU/veEzBljF5rEn+03ucS9sYGY/sV9h63aMSM5L/8d5mtQP00OU6L9DSBGxjLgW
Idyr3R5hPAq2UrKf7qM/MJgUKco0d81YWkxY7Wf8tVgi8aUWuIcPW5VnDCagN8X+3QHKaMQpnued
BOkhWvVextsAhoO8qlXgmDNKxXdl6W1w92z8LetqV/1An/GRD0tK+L/uuxmvDoPUXdVczOZSETy/
e477ZlmqwoPCmyOOuEzNmhDcwyyPgZ3WVD8nR8/3N79yzNYWSfUCUA4M8Wm7YmHoh3T1qw3adt/R
N2PJGVG8325cKGmKImYLr59hb7FL0Lu4BGY2zP0ux5LfYE+UZPJEadYtZzps7uagiPpEDRk60usq
vFUMNcdCRnn6l4CgCpfHaPbNI20ze93k/H/j7MooD/z+2726lq+sVd9WbyHDsNa9JXeDVqFvRRCd
EBA5VDVkA1zkCPW2dJjbD8CVlv9U3C1fQomongRkvTMtsBB1wKYbPM9rfHwMKLKxZHOQM1YJtaal
RikK0F42DkfbFhJqs+Yv2aSIxr6HJPZ42Lq1l6WmzjXlAoFQ5Lo6LUwwYMFd8keB+xj+ne8UsVlk
nowpMfBP3D7MZDngM7OWqRn6telpKmJ9KKjH2aoy5SN/9xlK9vXfpKcYS8WD67Z1gXjxvV9RxU+4
V4jS0hAFLbephDkn8Xc0xsIZUW1Z9qeeeDMdxwwKGs17+7ZPs73nIquQEWXdmvNJMS3wRQGO5imD
6iPQ0r6Rwb8xOH9FhIiIzS8byS6IIUQBbKAMmPAJ/YV0M7l1f8HS1f1BxZaYI9RCTyoa8y2G6xzO
d/y9rx1C8/cnPOwGAknH+h2zGnt6r+spOF6pabYIQOVfbIY2kCJav1SEnfh/CEbQMg4Spbvq8sxK
7Sxbr9vC1Prco0Yu+EwvUDqntTawps9tOXDnJbqCyl9cd84U3zu+eUgmqBzoTkXgvt3wsnQZh0Dh
roH7qaXQu1Fx+n3n9Wffo+BEOW2g/9EqKrhUQmQ/yvYdO/Y69+/mRBumirtt/S+PHjZ92gbJkoxd
hM1MVRXIjWHfJH3VhSrtycmDR2ZuVvQK2JGVjVZtdoaJbTVq5SzFa/Cj5qPD/lXep3DeGx8MjB4k
JUZwWhqZ53dI+x18yOYnvYqVJ5tjtBeOd37ixmUyMj0PhLDokbICTLeMtXFdk6Lg0dkg1tzRL+Pq
66WfHtrWOk6oAtutx3cSphSelsf0zPMpMX8DPyG119LrtHfg/mabYRlAEDt1okf4Y2YJNQ3S2s97
7stNJgjUrqg6/OoVD5Y/6CNc3M81OsNfeQDc8p3QNKgfR39yqlfLFcZ3vtHB+n4f4XmUyIelLzph
3f/J0XzvRJpZnhl0jIPJ5R73w6M+ih6d9zHgJeJYvOJRmzKmWt7y0oZPIRRH5+X96cuubYNG1nrI
eGMI2wtKB7yVWqg7uvzWn/ShKtL8BwmnBoIz457aZ4LjIu98mGRUf/ZJTqTJnAisl6COV8HeIj0s
3T5OmdJ+vUXALF41GF4siBTRtNPddN3DeUO8LsqFmWgSJvx9KXy+CM+se8G2drcqzcpsibqNmhlT
X3HXxpaNA88W1oVJNecT35KsgP/IxYuEmZB3zQEpvtWiP/at5KQLGqQ872Kgi3P3HppBQiJHy8cA
pRLr6ivm8KbhPoZj/m7nsCNkHL0gL0CcUcS1kUEz/cntwcoohwKpU0/iokxP7R5gy0RvNqB2jvVn
IT1IW/OrP0of2GPmQzG+ZdPd361xCwhfDC6ERmSHzh6kKlSEJZ+FGFGGx5xbuZa1K2klUVmCCp/0
5tvtTKurdRrFOUAy2Ys5kvnRHRQh9+7PyYuDTzCNoCoWLtUUq0N4sotxl6QFIkBP6I7T/qrs1NHe
1hT1gzYkHOhm1Y6b9Jl403rw9uhmWQAb3sTbPXpzqpOtM7PTzgZvgstP2LtTyseDH/7Hb0Si9Cam
WKYJKIh+FPaQHHN1VG0we7HQKn1CjPn7FOonnOua0GVr4VdMwXmQh/cf3Rz27ZVgl0qHWrFNQbGx
7Vp4Mjgh5StQdQ999UIVtrobIk0aE4szskMFYdx2VVX/at4SMaOhEcbAixjgPOx/2fu0dyofCx7y
41QwrWDek2uGvH5pgpAulhJ39b4/zbq79RZNTC8h077DPlWdIDboRT25kf9MQce7BNhtqs96WBCH
pLVZjmCIPZnZPhj9ty8oy7kI5C18YFtPdC0Jcl2TG6W8jNB6hA0sF6LKfl4hiK7J0LvfcXtz+K5d
78axccGCwQzKUOEXZeHy6gpY/zMzS2UWngjxokRZuKtovOi5r7hYHkEPLViAw9Ixaz01ngMgBpxi
vrVE89Y5rr55zecctkgF+S/htFEJCc1H1BS0sdM8hWR2RXNghzS07QQlrWBRRii+dzV5vsY63dbK
ddYBmd1MN8B0qTk5XEIyvcop7cPH4l/A6qNxXjSBg7rbqx/m9NsHz16TrXqP/iVDpku6PSz4+t0l
mSUhgfQ2xKu2Me8bEKPMWTMABD748WtPTH5OoSj28dubIWd12DUMtL38sFzppcCUPSwz3Oj42YwN
A1f7+zZdLOHDZHQAtJVGrE1Eh7NxTd3RMWw6Mla4WizWGOKGJkN+D4d0waU4Ml0BZz/Rg6ZZWT8w
wlq0Nv/xWh01FiDNq+MssMNIg3Lu/nHc908cCspjlF55zgAMtpSlluCoxTBwJurjG68+ROOQPqJX
ks1DTgKuYOV1uSwgpWO/sPPvgMsKiAHKQSIYVkKF0IFdAYmaPUsQ9BtFfSuyOXDbunOq8A1OiLFt
rAcdIfKDwqChKQvio0y7wb9bG1OK99YHXNrZ8iXbe+vN556NX20sX7HsBJqZ9MSetcoPg83b7cnn
S2qIpsRwkbPr23Q8Ud7avOKbsgKcN6pncLYZko/QPbWMN/XNjf0VPZLO+/wXuMGTpJfYpQAuOBLr
I1OiSYQpYHgJZFcKf+kQA/7KOFFkzVqJNNGS3wmciKU+ItYqcRWYhUXOZw9xzOSPP/F/S3N3+nSO
ElN2a0yFi8j6MmiqCc5c5E4bsW1atqTsQfH4ASwIpIETADCFg5C1J21k9EkxnXUwCEyEWgxRVF4o
seFFX6iKorKPepVvGIJHIeVXhvReYltjjD06tVgCU67uosS5kaOc7Lrw6HjFaelzXfmxtPOFYtSf
hb1dWUG90rspu9BaLpZYmdNOZ1m61yCYmSlVO8Wqcc60OdfYqnGB7JnZrHDVMhhtYv/GXpmwioC3
mfQUmiV7M3L/Cb6aHmc1lBgrJMOcZLwIleKpFn6CYJsEDq2JjAQkIUrRsSY2Y4YarFaQOLthUfqu
LEsexYgPle1TdsjyPaFNBRuhYlglgkrDdfAklT6HYoX6LurokWV7fSf32ZmyNcUuAcKYpmhWZm/R
AcYqTqFhDAL0uzZ5ZH3wNXfgT+pPF9yBs/7rHNNCa1u45IL8IcLrbuoSa18PPssMf5x4Lj2KMW/G
s4iV4FnXDTqM4AM0Jbn4iISphzGgIrxtI+T+8s1aDCXoxgAczr2T/Xtr4x3xAH536U61BSoOh6TK
R/+yYHG/71RgmwTTaHaKaAEJf9F6txVGiMUo+7QS+ohwNi1N1xX4aG8Pst063wdDL2Q3i1EzW/Wq
ulOa0Ckna6SDuI1WELZMHpUl+YJp8c7VL7oWd0PBv7Q1gEfcJcGgcOy4Pvl6O38ZLDFC9jHvY7ZP
vBjEPKVXVUrNquPkOyHtIVekL5Yw95/Mzjr4WSiRVb3Odf+14LH076ytd5zjkW/loZcdNlgbjDLD
7/2HAdNHBynrk/FFtwApih44HfXZV7LunXEs4GFJ2vO3XB3SBmVDEanul2LMAyEGkOlYUZdM+LB9
WFaaXpZIinJe0g6KhXtI+g64SqQY3SAss0jRdoclkIYPUAY4KLCHAxwMZP5pMWhAj0PV7UKS2ho8
XADpmkUwHAKSjsElXO9gMdfPO9wlMVyXp0LWDbnLy0IAaXwT372hpKx1KsYzFLfd+o4pleiBT3VM
/jCx6GpMMHlO6hlbGnOBQZG8a+meu6uK5RN7/ACsEAUTHbd9nddCyo2dSJyJuZXEKUo7e21ikKsM
Us7e9NT59nmipxN/rbNI+CxRMn11tiLbfMNpiKliOzEBwGZSUmWp96jGtjMoKTk77QtXA8vfigfh
/3tbjfLKfS59uqPAb57/3vJ/OvFX69VGJN0FXywGVt1xjJf/IFnkyUAFV4+yzOenij3mmxlxXVe4
NlyDtzuVOikjTHtTWh0i/syPG8dyjuz1u9PUx8IF4BT3ZQCeEIPGeI7xrAiXqOSyqkZV6h03JNJE
bOlEByC3N5AT3pvDe1oiBMrS7XVioNlIGI2kFCEUW9FB+qx6LsKB8b+guZI1+eDRbQPThqP8i1Zr
x5FiMsSnx/93HP1Wqf4aBUjB397ALRNH6tYkyF5M25TMDQ5sbSRd+qFpB2lZSZh4RLWk9L9+MQ7j
7bduObf1i6gTXh2+zcjWYd9nCEgbIlGFdcQOzaOPZA6qeu3hU5X+X2KGHRLYPSRwsHVqcx3aVWWB
VcxjDYwDhD3lOZzP3uv2Q3RSFsLd0Av8wuzp4j2bWy1+3ArSsWYD8nZ2JaNEyd1FYhVEmh21sgXI
HsyNC/W2ZsNmPh1pqB1dy13+L3PzHY5PEyXC53q0a/3zsMHyHskIBrzv+8djYJ4OTkrqFxN2Zgok
czlft97YH/gmk6nh3aa+LyREkBD7NcTj6ZYRDBAVtXI0BlcMS+pKZPjRYYHA5uvkcvoPfuB8ju3r
5mR22QSRTugmhWr4z1oMAPVYa8s7MexukfWz3KO46Xrv8pwTYkSvKPKj0si0jzs10Ad7qmrajfoX
S8XYZ4XVdNZ6bGA2K+1xTmGXHqlx8Kw/l5uADLPA9/LeirWOQejimLgkcNWhpugalPxw1xOcKZTY
UTNtzIablgeDWyAZFRfc8OugyWSsh6Vtcx6NheFIh9CRMkXyN9CsqXuGG6DJzkntNhwITUeJfVxK
n27Eb3tYMtIT/IR927Eq+rs8ksoChcJD2EGzp2VdzFjyZsjUNKUBF7LG+D+QlYENL9PLowGVoELe
Mmpr3OrOyHx5Iz+8bihHmaYfNG6Z0dwRmoqPR0Mz0txItJTT3JgxSMA05E0501mf7IFj3pXZ7lVn
p+YJE3pnSWcaUP+VxctXd+yhmGxUA8KWgZhyX+0pk7rGbpvvevVG2oDbBhXjNQLJBfz8o8B+MpZg
AYbKe228Bnps0+Fi/QigtBJdvkDXFupcyEQifzSJygm3BNQIiXyqndSjywzIL5+2uJxSXv1KLKDw
Puwx55WNrD8PsCQOhsT7/9tqV6Ncjp3U5g2yF5PydwXgdaH+Gz30qfnqeCKIwlJM2a5U6NIgB52H
u/6bUCQIKcSTyYVx1tlqnZWvCrJ/vadzCb+tQ82759ZLRKxCAznMoe3bL/Scwa7h2gNQxal8FTWl
N6rsxm/frDpe7GKnoeVn4wTfuQqfZTSC4H8W6UBPnZHJA/33Z/8zLlLlR5gY9AqgO+DD/ypN9O9g
saNvH7mHJWrJ2ed6KJbLSqCYXEhoOIW7d1qAfqTarHj1lOtEGHHbG266wY2oApAZFIZkyRzqQoFs
PxrjEVDwlGytiz/o9bLN0yJ4K4E6NZiNACTyunzjhDRw9kyqCUSVDbGx0rgeUyGPHErKzZfkGQ7Y
SdHp6fFCRo9pUFSE1CEaX6zC7sqqxpGq09yFsnxiV7NipBca7FY26mcPmW0/0ikTnnYxblQCNa40
pQGa9nxFHxU+LuL86Rwoi6uZvzg6ppm/Fv5Phbiuhccb8EEji+NH1U1BayrBceHDjLnFGKsg+iSP
0nv3gnCqcnsIXWhCbumnkp7VbCHqyLWx40papawvC2s09mfKJfqFT4DE8k9TRXt6hbaYnH2kbk+J
yO/hdtSX9CdTFP0QHmQgg06OEoZgO820k4CE42FzZBrSPpFGF2I3k1gAnjESLOPUUJee2jivRs7F
4tJQIQrRZdTmQgkjOefQ4pykrtuSPtHHgzbxiqGuN1v/Q65KAjQP4MV04ZHYlvbn4K+GJ8Sn+w0Q
m84CYqdjz1giwnqq6nMOnscKFxoSPah6ForyVmYJ83sEslPFs4069APwqSwyF+JAEkaozV6Z74B8
IRSGrwuCpyTpcxbRiAsxkMFMBwcWRf4Zamg4xjC0iSf1nXplG2Px7Ce5RD3yyMYYYnEZNaK+L0+s
euLivqaVvhKtCUbwQJS7lRU0RqQSv9IVfQ3sPDa3XCcxL5W0n+7nTjHOnipn+wpsiaDIOqZX4niT
TSLmmNYZgb/0CRTQSAF99mewPsy2fWCMcFYrE8Mh9ioHcguJMSmEJl76GcikOxH59duHgdVshB5b
gkWXreAjrgV6R43qKcHiPprzKk89TfnuQiQnjFWi7hiYHKxj8rc/Xu/DmgHNPhObXHVYe6+b9quJ
VWKgLeBvqKGLd9eTdXjztWzcrK3oQufXOtJxh2fqi9E+OUIlVY2lmdr6bsKlHqG9jo0Mw24bAgqE
QC78iYfzPGBcX5p8RFq8ZzkfSAjKq63ftQr9ln07HkO8iU/VdTAwhOqE+Xod2HO680OJXYR/a/Lw
VPEIMqoagWJpRGHQgf1M+EF4LwyhY6K+UTMLwRraYOK8xylEvk9fJgWMs6DhULZRsFtnR012+x0a
XjRC2Yx0EL5GSxLvJV7PNjTCD6YjwdPRe6Nvjyg5OrmxwqKhqGJE+ctcOb0c8B973hDauHXXvp6k
L8H4RtOCDtptSPR0VK5La2EMFAu53irnLEZLrsmssRWzvUPo0a89QfJ940cqNV3k9Fgk/jHdmcx2
30ePPvvRnWEyc3+kEnjDmFVq63Vu5FlnWOpvOMe5J3y3Wd7qqJCB+tt03Yipa+K57cfsLuHRo1fk
sVMg/M1Rf0VpkdKuxqRmCKhF0c1ZpcG5dk60gzCOvHRwhUzF+rAT9v2PBLOcsTGpg1A1G55pTJZz
dUueRwtQgx6jlXQvhQGmzTdtttKCKXrSb3CACHWyNZXyV/OaIJBjVEIdRkj8iTiiHG7OEYumPDwC
Lw1bjmC26+j0JzO03nHYpNZ1SgCtdzx2fBq5bD4sEVK0HX2MHbwnM90XnaqPWAr59n3J3NWzI3hu
TDYUB6SR81DCN/WKJzU805U/BOKTNPWhannFSgqtfxqBlPXUOsgv04LPwVKaG6ZC9JDZhGwPL+Vb
WEZcMqFLeTfTyW4OdoJIE9YfGe0UFvlpeCvag6RzalZtozTkQ0te3y4yWYk4EAx41ZcdegXvbaoU
QT1yFRbKxNgosBs5sNky9WKuOHZKFh6ZX3qygCI/jMvuPtlVLpcGIq+1Ha/N0RyKO+E1WN+WPbMc
bL6XYcg3q0kxM1urBLFoTxSThqC7/TlT+vrFrUWA6cclh0EMbQoCgagKJ0H7rVztaUYwXGHZj7qy
XdgAnZ4oeOSR/UIE9tDZxA1A9MMdcw66YoWjB84JU4leOeuMbzxHeBFfAdzXoZFriOwu+R5CYhVF
Xx1/gEBQVcYQgFaUkfBaypND4aEfpKL9UT8AWnnnAzro1XFwejivtIBPi6LykvOP0SkJHmyQkMro
gdYx7h2aJiNM8oqiDUqk7A6vpRbfElSp97Cex61rlaYmxMz1CaNPgOUqZseaC9/4L2KZunxajrWa
nTwAL0ipZQXqb6WKpV9kz4o/hpzoS+KnFijk6I7QFwYVcwZd0q01mW1GX7HDc8te8JGYOfItiOf7
M+RsQWLsIeMBD8ihCd/dRTj+AaFkpztyhTl+hmhoOHSBVJV2YSNhl5KThiUUjNIKkcutnnBYY4Fy
m+peGUjBeuT25+sLuQ0dRTBMJvGoYJ+nOqzuKoJ8d1hi53rPbLHkyIb6ges1offz/40/GZr5VS4d
9AaeB+X0yh+ii5ojPfKEMlwnx9LRh4WMWl6P7oLVKx97jnUvdAjFnmNDRLqfuPk64U66H3zXsgyS
FZHrkWHLdS9LlSLdL4helqmbAq6P1FnN4VRZUd9Bnh1mQWQ/jefVcdhCMFi6wbfOYI2o5//Tk1bH
mfWfcRVds5DW4tnrba4PXcjoxd4qo6MdsSr1r8KLrIV7mdrPWxm4JWq6sPhFKdquCk8wRqGA5RNC
fgQ/DvPfrzfSmwWZPv8sCj3DevztxnhpQDM8g3W93ykxa3UM1T/mW+aRnb1wPcwj4ALzgK78HrDk
aX5GpQucKKYB0E8Le/WubYOerj9aB/RHgWf7luSxGe5T5S4eoyzBtzWma2n2hR8eUH37+2/SXemK
/XaUf7Bw4Bg6ABeikyUtuhnYGCmbW1nwcq2iwCozeJPI41SOIOObu7eQL9IYe1HW2WdAf7XAUi9V
H6WVrmRj5gvOmZ1E8od7EsONoobEl2u5VWJAGT3q3BD7U1oLeRCw+bc8+WB4dFnu9Mz7mB+HwUhf
eZRUy5/QGZstKm0T+QMXjG10qxY0Su4DAsn3n6UgRKtTMasxJO2ABjQgKji6h4q/4zSLMvoU2+il
JMOowBrnXygahUvtnL0d/Q7nTKczIM2WLP6ZQfDtKQPKrf1Ngc/H20Ip8f/UaSy3pdjp9aVfVFu2
pM9N3yCnU9YsO86QOskjjT1UbNm4Bdvko57sPG4L1COHLoQRrwrtOHsvJR0cMgcfFD3qG5S91m6H
U+kVi5bGn9CVxwuDbptiUEGfSd9e+QsK0My0dfmkK9RJ7lnBLaKuTFIJmxbUvgNxORJGM4VytGUx
NkzJQ2enfs+1CDVw5PwCDfRd/2ZWkepC5ronXiTLVfJbi6zWGj/0anz8tEYwkcehiJp/p8tAA88+
0SavmqkKAU1y6fQTNwJGMH6JdNlxaqRC8sbfeBpJUqZdPUHyyg4eRjienTW+7HEfEmlGdQINzb7P
z7pH9nWykufh78PaWalUpFNVNXYTq8yiUBIPB93WoAyaO6wS/Axhk8TR47Ppgiak6Lfzp7dqi7WB
pl/XPVdggiGYzxlG38r7ZVEe/F8PQaLikM/J2CMgElOsZGcnZF3xYGwsh9lJSWNqSO1mK1S5H2JP
WDSKTplE9+0WotCu231wohRvnquGZn4BiLXx2RReaBo31dXsGgH0w3xtLpoTyYrnd9Qzl4RUSZ8a
bkgVua5z6rNWuFNrVpV2rCxGBZp4nKBrhwwTp3uM2cnb1kXWFN8H4560aHCVhamTUqnsMtPjmbg8
8Zda+ijqFDxCTkvkfhhaHk6L1w4wgMV50PQiPtqFucshOJRJBMnGf1FSTdCTHjlgyDmrg7Ga8pVY
S+0UesUhF+fEvn6Mrn4lPrZHGKcsTmI5PxN21KkhY6PURYZ+J9iUJkOgkVuqns/YZ9gQc1lBsccm
2fL9FxetSNqPnVmD95dB+/SD9EaaAN6FfrcRhaEwPESQKue1H+C3bZCUtLfNawgt9wiTDDjwFp6M
Xh4S7P9qih8yC98rG16uc5pJYPA12znypSE6VSpztsbRU0KbsaQX1HAZ84A3BshLPCcrhOoAAu2F
BIm3Db6tLFEn7mzfU2euHjJzONCw9qgbigafJSfNgF/KYSjyTPzT80NAbz1oPqhrXr8+ig0SKLTv
svw4l35d3LlVdOYOooAGGB+q/H7LDJ7ETHtbHlakDnfVUNQcPAEtxx1fj83Y+ALeqQLEL41uGWF5
Osgr5ZE6g3q5alWY+jStPnZAwzxsPVAIHrnoAEfW4TU1+jNohpEOwq4hqjlk5DonBI7I0kGbXl42
zeI+kE7478Om5w67xfe9OElTnPbhpF7UDJM/14TJ9mVR42+fyBAGP+k4GCC6wh1c1MssLIgK4yzL
Sp9UxZxReIl1T5qZW9SfdrjNlBsT3H5qDrii5E83t1WdBQsDCWx4Dcuu0H7fkHgjah4PPtixdTh1
IgR9sdQwJSREUnKgnAScvoJSUDMp3UJj5PKZ95HucbEk3Fax56Oanl9DK/84pYvm6UIfPLChLj5+
G1h+mMC1noQHIUrqK4xcjjwi/K/3qT8uaPevx+U6cD8fnPyM4BuNaYg+WLTr4G0aPQGBOCxP1ohm
Nd5l1XMJ1goaTs9fjep0+GZpl3O/yk8eriwb5Q6wN5SBaRT/Da9GQvQo2tSU0DgyW7ysMhJ5MRKm
hQEoWKSp/BmKOYpcSpwQhco/HcaHlz1SvjdEBCHPAzLHf5kkT6L9HYqgnyzFisfSqJI0VeX8Pikw
8l2oM0BSqmDQ9PoWTXmUIHSG1IFyeVPByqggr5LHZ3Vgmias3sicBT62dBgr31CUspNgFANljInX
9Dkfs3gmaq5RuoFcFXgGlX2/67vib8TULU6yfuaeFx6vSPLyZ8PxB8xdTOlaNZHk4lfFk+/vwqES
oJ1fLcDx14E0G/WEXmDtD85kfHP1hS6/2Pg5ckUBJnAIBKtDr6SPSScKuXUZx4DnJmWiM4a4VUIv
SrFt1X3bEY2vSHRRZ3TIYNA4oCyZ3c4Je9dAUfkp5CKCrsktWx5ggAOi0r7F8Q0VLi7E+VQUU5m9
86yfq+9bNOE5whHDTKCYf9o9eYVJI2Xxj8ovI2bOtW9cK26vgBnTsw0NanQGEDYKaxQazqb+wZeB
ly8+3cblX2vE/daL3b22YsKMvX5KbG5Ns3CM/pzpJChEaRZejM7MzFaaX3gwuLdLTE2mE8VmIpG+
dW1sFOOQstSDtxkRJSGITyJnAm0EwLTkDtsza8BwcK4SOWf4d5jMWmw9d/X7cXsOAJPvtmlToBto
Ix3IB28MPlGmF0bom4nmYgxEdHhof3mYEmqqXB/6VDeTLXyyl1muNm9VsilMGtQVt55dfWf6lr5u
NCA+rRG2JmrPO9lae1YE99bToO2/pGKqUiACC9arrn59Dqkq88I4vn+5DaJ3JvpB74B0XP0HkWe3
dbdZHa1nQ0MQWFOWXuBL99kAySzLKxSNTVtBuT8fsBi+9q1vejpHupXKmOuLFF44N/i1s8sjlDNX
4ovMGrVUEbYBKPqJymzoOwl3zu8dhfBp6XJ5K0GJ6lVsRVlh6uFIOf0igFnWXwkrNjA6rYpcn/oL
Q4u+tnpmCIzSseHTjlLZ+eOArGOFVFZX1Yw9MwJDl9pgfQe1K20B4HQhpUeCgQTOcn+6EiWF5WY+
s2DNm9rd5BI/2uGLN3TN1oMnzp8Ho8NnMQU7rsUDyLGLbdXlQqAGrFgWyUZDeE9yXV5b967MlYtg
ih4/RnirUph27Ci9j88b4d02DvOQ7qBRTXBlujcbi3/gLpQAe5a694/5hSO2wHJqL/0F/AF0KWe1
1V+BavU0AHiRHXrjlThByT+h/hgmhb/zwFzYzcqoClSWZpnOXjnn0TC4TArE5xbOWl0kZC1Y2AyY
1sb8VrtB4qT+SG+Pbwc9Pl/ntaeRIuVnwO9MZsJAPNaH+qPCa6RicuypdjWP+2cZkrKU4vu68Mvp
dZ54raQfqVBL2IH7NvJojuJrtiCS9Bee30+tTLNWGf376/XOZVZBSEC4AvRx1AK66TZFcn0WUF7r
IGuiL2IoghjIoCc7AgcOWrBrSgeacKV3lTfV4vA7uvn8o2Bj9f2y0CJVzcukXH2wrb0Li7QPMX/V
N1xfUgKm+TV8Zn89RUSAwBs0nGyB0OwVDKf17kmkxMS3I5knJS2vb853qHmqfQCVy1fB42yGk92l
WrrIXgyOzPNg7ibdwQy4zFhgHbGfRI/veA3woyMElvq01NlWL95DB10o128a798aaoBYfWH+C0P9
ra3IaRAqk8esS6aIYdXAhipzyl5T7OX3Df9YIXEtxo9fEq6K99l0YoHgbPSkh1iR3tLLPJ4VHyCz
HmWu5w/qePZM2oe6Q1w7Sg5vUebY8Mt31PjQFjFnINVa0wvtb8gJL+eZ5Xc6BqNFmzsU5U8GUtqC
JFGqstahQtZJO/ACS3YR+69AlxKoSdpq9YzJFfUXgsiPm7nR1rRJ9CEf82Zrxdxt1+lAi8broY0A
OZtFRia6a/mi4NNDm7av+5ILbeXQaqJP8DAQLiuDUWXo3ZvaTKnWRQTy6EBhjqidjB1l39wsdRgW
73/3O/Afiu6BAC3uHBa+HBt6E5TzwYzFXYTJCM1JcR59VUKiYdSn9+l2c8eLJS3+H3IeHoEzttD9
ldoEe6qJ7gxRZE9a8LeMgwSotbbK/bqnGs5zI+Fl05II5BQT2xrE9YLzLuBsdcWO7hMAr5f+ZYM1
0c+fgzUtpmEvzFDyDgTqwKOHqkVxuUGQDtMaUhvbA3ARH3VoCySsUOlQ9OjZJaPSw/qCJ3o4jxd4
s50ysQQ9RAK97DpQMw7zAR8kWN5AmwSTDWRy0GgpgyHxLGOOe5JvveqsjO6vcgfAOA4kJwA6lH/O
c15HrZmVao5z79HK1NsTfT3ZpdA02z/0yiUv54zV9+CSQ6zJuHPrvvEcjPnEqnXdGloExuNp3sVt
4u1viZd9NnVVrAE/u9mD6T4QokScqWIKRhQEinkcmOBRbaVglqMetcKapzw1scHa8/yW6bg7HWdo
EbVAmZkzbnoEkx1XqCV4IRe2LVV0VZy1f/nNYN+j32E/4y55279b7g2HdHYgI0AwLMcYO87GT7dz
aYEeUmoKOwSKVOc1W8paHTspJnfCqbpnzi3cyAIMncBMr2nUx6T+x2VoDmgpT3cU26kmJy3HRfh6
cmsQGGANDFEfgN9B6ib2Wew5Ydp5kea/s7OkOSwS04Ctq4r/hUrTaMN7RCXGzHl7r7kvfgk8XaiG
FZSKIcowhsSpy6pu8lVATc8eZTr/HFGRBo7Y+6FAimtMAGYsAYPnnURuJzqLO8Rb3LzvnK8PWFJz
1KlJuqb3jmmHsWfOHtwEqvwtzF2TQjH1AxOJVZzgfm9uNlpCNdPT0/ePiP4ZA+xerC3Ayq3K2zOg
Q41MbkaibcEVDfhsM4NuDDNzA7SGS/itx0Gdx4upfWZ1NBBAIESlB5vEoZPxTcciFqDnoph8kCM8
R0Wh7xXIvN61/7DEFNs35WHEjlQp3tyD0Q6dXsNAhEDCnIKBLN/iDNcA/+KSewOBYkFi09ASF+Vl
UrwA7WdC1XJMJBVoUSWyU10/q1yVMedVPhlMhrsvljCkxB2xquR3mjXjQ1Ry+ZzB7bzFEBBk9BHh
ayIdQc9HARkPetgabUmr1hsBW51/q317ToV++hlAwRRl6J6EtYVN/9iHG4Xu/f16whPZPpnl32st
0/GhVBCgxCNCdHZj1xYZhAzaOhTSueOKTlPEiJnJwYOrJ4siE0Le6g2QB4H0iVTOA31apvMxYaMI
uoQ6J01WW6KPPIiOu3tbt0MWS3kBqP+8/ldwkDARrcXnw2dDL7nUFwlC/slLAyYydosUY/G57E1w
LPbm6RR881RLgcn0czhzo+SD8t3y+RDNBif9QSwkg8qVW+4IVtWhQYkJpZWAh/8DUR4l7jewN4nF
ZwPAzO1EJ9EkF4k88ctH7mlT7A+dtuiZW/gftpqDLICSQmYCrGS7XdZgJFeN1Lz8ePf3NzE/T6X+
B0GT6jZIkW/LEtKrwDnB/+Y6RHLLAQt122gRlYs0FoCG0tCU3juVb0LR42j8lOXnjUoFDztSYD+k
KKg7gKXnzHCl5qs8FaaUPLaDMr1jb3cd198kh6RNYnYjQunQ95Ie0Yd9TkdGwQlbzTAROwKeipVp
HBbqTpPgr1dKPp9wlcFhl+G62PBrUIRtqLPGXnbVkVnLKYCtMmHvsH7Ih1Z1hdPFjxPHc4QXzE1v
ixRg4+zhmk+pYeprwAaryxK0Az/rLaTl0Lnp5FcOqwWgEeWDmy7Kx60gLkuOCV3K2+FihzgwaOrQ
tVlgH+92gEcxKCFUrbnpG9kfl4whlhcGGE1iJVVr/6ubwhcURtf2mR4XVZaGX8itFEUDyj387ppS
ueswHvOnF3/Q+2j5PIFOt8L8AMSosVemQc7g5sTxp5ZQBIGmuHq84d3SY8p5+20GNMxfOLhyxCyU
hLslRG1DrI0cnXYZMu62WS7eQ7ABe4NQA8Dy0Ewx54FGqlueyaAXe8TdTm9tg6rg8brrvS+jZaTJ
C78hCjMOCe0HEecx05J2Toq7G+FeKG7OzWpjFCsGFl82ohlztcVzwBQi8OkYe53a5Iqe+3Yj98eV
jgDIz5AFDoYSj4d1UelRMuJ4VZTvRfz3Uql43AHBvpPo1nJld+6gvDGyrXxRMlnqpg1SM3bEjJjt
22cdhOeeo0YUK0prC7RGMH6FXUI/xX+6D+o8pFD+OEsYEgyBH+H22RZwssY/fsmlXaaXsu1ISxSV
ECBDCe24DBsyE0e/7kW6bdNBHDXCVbq3ovcKvLDfh0xjySiehQ1G6HbbDMsIlArJ0ZH+/MRm60GU
KwvA4vLYpZtXw8mz+hufMlFAms74lzqYsaN0Asrh5KEi82bVGElwPXVM7c4HEunlADLB8LKRotx4
cgCOk3+ZtcNho1mrEpIARf7Nmvm5Z8HmZZkQ9zMMKng/3KXo3YAOYEj6trouVyi3SaKI6XfmZUjG
nun5fAeKcj74YEi0SyMCHSwSSpB/aqZYGpHsyn+bUr4if6D+UcDBCBAG7TKFixKhjB1nif7Ll4Jb
iv+YI+ov4s9mOJ/LXLgCcUO0P0as7DoDi3DyY4zi4m8lS+DKrmvo9wY8YgHj92KBZVNDhl9wx//Z
CgSGHvKxtwcd7ZHeVIGE02NCIoeTDqwg6sHuKzZ5JyT9qqtcYMNqxKkuS6DzxcCsT2TnAVlJbC8J
jK7MdrvgqO/c8Oh4GsFv3vtjDfG7gtPDSk9usTUTzj8aGdpBKJ1ltw+SvZYIj6v+PfIFpSxL4ftC
WsbynNHi8uD/DODI0wzM8+udWwJk6JocT+wDGJY4r2A1LqprniOpNYOOPmkqTAmVwJ58vPSBdMwE
nqK5hbWVTPvGPdxent3/dfTyBzxzZzZydgm0+F4ACB3Yi1NbbO1VK0UsyIAub0ugjAw5745ex+bn
R1lwe9/auvgkyXZlfxAobpkrQRFd7nD9sSmEdWJymryembZRSOduPk7g5iJbpK2MYgUIYBEYorjJ
Y+U9g6C+31eEWVfA3QqCri4pzmjyb5xZZkM3mv2GsWND8N8Rh1mN2yGf9xf2qbevX9u3WLuvDLmp
Sn80AyJecGtBbcVBjWqeFVzB3EYsrC5w0TONi/1DFwJynMZi8sE8NPfx8ujXRGMs0V53AK5ezM5g
5uZeNQ9cYZ8JJQYFke8HommLtLArcfx4SECqFZNUjvtV0DR4atOAdlkCJAKlWnGgdIBtJXjSr1Gy
9tfKrCBKUJE3SM/0etbChuWFG0EjrsDsoT9Xqd1acPf4kM8eJYQhNlRFlUkey86pA6rO8MUgwAha
F3v/ak/Pwjn2llQ0+4ElyLtevhSYkzyh+rYIunI2huwVSJQ5aEe7yHXuBitilbNSix1Ix6oGRJQI
hFyAum1ht8RICh+QQUKmGrAX4k3QJUOFvGHM6dHuARoQWQTQjBi7gm3KHp9TIedB64pR+E/+p3zm
6g2R11gT7vqDEu1GaEQ41vE8npHP1AyAvrnq2DGS2H3aZFAXCIK5ZHrKZxKB9thDyLRnD9hlbJpm
sk0JYtSKU9ao0RqKcH2ElNnH+2tM+j90Oxm0mlGpIfbJIh78ucjhKsRvcFQNjJqEGinqnfnjbpUe
jFF53BxTeMymiovFTboUOB5HFbUCkSJ6LDjP0uHPOZnEtejZBZKQchDz/MBEKxaGV0HRP3VtcyHV
c6emE8bG8P/M687dYbtpbREkz9nJlI/ovu7M+6czF+h6oAYnsj4EcUZTgVMAWrHUp8qDQ7VWNM37
0sxiCSUmgBVXDr9Qzl5AQLaXeIFS7VnnHvB3+VeF4IWQGMutkpswAT/tMTko2mo0ya0aYj/Sunry
Vo4j2Lf5mvOQx5v6QpRS/rpBaQlz+nMCsw8WCU6Y60K9/rGhs24ADZKtKQcpM4vQXt1GLqZAOFm4
GjwBKIoDxmwJ/hYL2dqCKAUe2j5/OHDvR5BRzGzRy0vkhozFskIkQKyLdEpM3n9f8iqIUp0FZj3Y
eNxfNBjbGX0RgTqtm5fU8FkagpFMFNrdePOnJxppEeqPa/b9Fnd8W/27bPDgv5+bRxyjYvHh/Pye
NdNXjGj+oSbrwTF8FjDdn5fxoCZ/Ih2kwEIeiu25QXOqdC48SXC7O7z1svDeC1AZ97WRNk4pdven
tLeB/Wr+DZu7IcBUmoAhDKmKzW+Eo76jfjn470KQg19u66YaE7pChyLX/k+ZMVP/o4hKPMT6i9Hd
XqlmrDoRf//GqrD1pyk5yGjrKzKgcOpsMtYq60UfzMO+80sUONJyEotQRZTf0t+INP5faOaAhI/k
Vw9wysePh7UBeJlP3iGVbmoOSVeMaPJLTCYUoctHNxyXDVggugXpKa5IvlV6gyjhS8S+aU2nbiNz
k2M+93adc4jhyKaB81JCf1jiqXPPoxNX3NgHt+JJ63w3Pjsz+GW8cW5l3KU7otnUfPcLFexQdjEo
ht2HsJcd015MopMNDBjZwdGPOLJwYU3ZA1sxh7Hv2Kc1mTEF1Tn1MiASmrFLPvpv8gxkuyJVrK2I
4CmgsRWUKjWtALESrmuR4Dp+mXWKTZZavd/C0sMimLhRvvBzi7FmH2LbY/p9+dPh6OfxJYZlqEig
hgfCrnpqIYfjKD4QCu1nKV1XD0FhXOGyEkoF3BhkZlADUsRXYPWPFdZUHpzIM2++lBx0vriIB3VY
e5G33zmYlhn8ygJ3p7MX1ag8xXdcjOdYkk3M9cQCpBsqahI/BUlLw8V5QtmOZuMLaF18W1mUL1pU
a6dwxgYweyXdKmR5WLQdO/kQI/8e1RwUO/GJbMucgs9Akc7w6aw5ZvdszFwrQvos01gvdJfzFukj
AqPcH8h4vw0f/GUzKCGggFUS+ce7nOH5bv/fDXI0ESSHd7+OoePPq3YT3RrPYPINVMwdt3lHPJZy
csP7/JupGlwFLSeT13zUkWKpFTRTblCPngq428GfWnuW87MnR3clmTIhk11ujRyjDEriclf7Yh5C
2UiNHkz7p0wP9llWEF3JL1ICDPNkscYocrSPXADaIzTQmR0KWcD3mhm2qtssudw1cXW7orxGCzWI
HkLKDyV0ce1colyJ0F/bF5SgM/d9cTF84cAxY4Y0d++bDsQeJ5I5VC/vYVavE7VjOovXenizd5sC
DMy3JtjyYoCWBKwI/cVGskrLUABH633alewaGTGOyjfKyjr2VcOkBWgNsxotYRfUsI4tGQzk6Ltr
CsFQbexbnQ9qxsNNiDGm1vTt5ZFpRw9f9Ghkcislh+rChEfbVfQSiX90TnN8tHI9ljlERAPgYTAX
MFyEV8ndJlUQ+yodWkn4DXIzwA2VB5zGUXNp6MIJKUF1DrRa4KJWXNyoxuwLqbiHUetnKpoaYB0P
vFm3OCUpZ8JzjslgvwvRx6V3dcbfPA+Ww+y17+cywjVa7SR2OtZhgmIFmm4fdoxPx+0ZrymK02op
ABMLBvcuHMqVvihRZA7NWS8RktMZggcA/FzzbKq2Qq+J0Rgw7dI3wPX/0QeTw7XR+ToWqQYuBGjN
/Xf4Ya3ncmHC8dBDrivkeS8xs6I/A+HEoVBmjoUbRrlkth6FRefTRZ5zhrn4VpmVoYNdy1qGXGde
2qgGhND05/qPFzS0wpRQRL6IJaukjD9VgSnQbFlRsiY8DYOVT5Yjord/1d69hBXtkFBhK/IMh4Ba
8k5MxwGdf6xvxkV6J8+8zYZLpwvCxargPt++rwsHCY4PPaZhRt+7f8I5S7WYxdvzJX261vZw/+ND
7hyfygGhMFYg0oEmQ0HUNn7kfzKWOwcBa+uDBALMVrsZpjB42cpWZypvKlXgsQBA1YRR2F4hNg8q
mm7Aa155X9t5Gwow3GU81hguAjoO+Ai/uY9JxSxrSFohOUbDCJoEhH2zhpwrEe9X1uTRv8Juvgb/
eVsY3byoHZrwIwqGpQr3ht1xgNbFeKABt7C9yrQBMKa4iVSF/ky1TmTVG5f4q3dZ138OIwluhai0
zVmyWzeDXIlw5Zp8YHdqv774UKJ/xMt4FKcqxmME8ms0Hu9g/ykYVqOZcgDi8wk+pu51AU0YKAQQ
L7LBAvdSA7nbJm6EOBLYQoStRYmoIssGzZQJ9mPEckWpKnS8/MmVh0dAVvtTJZGq+7V1XO5bYPFh
splAeVZOVA+V8pdCV3a77u+T2jmhrwL1wjmvRRPO1h2YUcRkzV/0h9lW980KKOzrch+KqqgfMOu1
A/yK79hGX6h+q+XrzK474YCGumfZmZyMZjcQWo1IyUsEQKX9kcQk3xWuGcSOXj89kW/GgPlIDJXw
lRt2madBrfi+Fiy2wve6gvWyZMRtFprWo5y6pJB2wixY4oR6C7+kms+wUGsKnc9XwDo5hkepQrum
qJbVArTj8TeKoACYgu2+e+CXer+njck8PDjQhU8GnPiCplHCfzYacfIeOqVfF5ttCZgx7su4Uq74
UoymiZYRFX2sH/Nw7fQaEYt9PSTJI4gzRPdg3NBjr2T47XqlPUbToeak+0RXXCsSCR6iLJyEytt6
fLbSGyBOw6atj0xZpe5/qq67vaIM83N14sDWLdtlzRmMlnFJNauwQUIn5nqZWkUh0Vo92rLohcq5
9yCxhwwGXk0J6rsrELZ/neHa84Od1Z4COgtx3H6IbJyhRHC6/WKZjhVOJO5hDDg9jFSkrpCS6mxv
7ci9DigWvSwd+1WQ1cndujaunEFmJJbYJbYZyG6+gBNHrznwbsYy8HMQ54zxXwtFSsOXJieN1mqO
gJdhfocyaeN0AB9q8BnN6TijThTgzDT+YEqr4J1J9jbqwnEv1g+uMDlxG7FQYpu9xlK45ljNEndk
kpGn1lAp9BVGhw86UER6d5Czp4omUFNv0JLViaJi0fxTz8V+2Ij+gMiHEplz5e2jUJCtHLmjGY4R
1Cpz6fTn7a7SDa8UkM6UzlkRxnaykwT4uCxlzEcFgD4K6Z/ZbKOZ6qBJFlYCN5UXx4b3sCMFOZO1
kcFhoE3gTFYHFi0h1YXGnGbynTZKXQh9MxMgULY1hYlY1aof65qYnxzExE4w3BhTlgc6rd6bKrLd
YQO+wwrqe/FQJboXEHeUhmvQZxnxx9CgO60OjoMjIawJ3Z1Zvlht4s559gkpfGzKJNSgqgFSqSOT
RV0l04K8iSapMIxnHW2Lfei2pb3Fq3Wqmoy4PA2HGQG8ELUp9NeZKgZ8MUmgnhmKLwQc5S2Y97Re
TZfbTbVgoSTkkUB0cX3642tnZlLxcuhrrusyxXSYxk4dOPb6gSnoCSD7ovZVcPcIO9nGHMqnJ6qw
efnI8lrJRu+g6hMr/X4FuJIXNc/rmnlFXNImIfP1Vnyqhux9BxVp85tg3w48ruRzhQQWNXS459LD
uk61KQ6eEYZMLJT8yPH6tUdmiYNJX14yEbKpsRSia5ESF/VpUuIFEAXbtpAw9jvorzp07Ox+nEVT
MSHOxFzjwT3dadQ6QmHbtvySsKYan1YEaQYIlKzVzVovLNbcjXQdrTAMuW/90e4oHrTV08Yweaql
j+mFh3OpZsnRTfCK9/7am2twdiVCDXt2xBOMuvV9b6yliaWvimCJ3NVOx26IL4eUb8wBlqFRpgsj
DA93TQAG8sJzCYS28gor4DywLatvZmB3dXqX6olZ5caLm/i3aB0lqsHISl/qTeazW7xYIM30VlOS
a7DuTGYG1/yMvx6Cx3oMUSkaiPClGdLlyINuoYpye98SkuGBhhek9IPjSmaL1lM6LKWMiQ1kAK6V
RcYuSPXrnyKciVcQijHwPa1AoFHMo+bxEb5CYFzJt9KObnKQdf1YyVRh/kGesmDx6ba57HNUvfsW
YIdqWwcoX8LU90OXpcoIrnz/9i0fH49fIvelsw3mEY0xZpSJ0CDrA7GCsXf/bExJBrB9GQpAdCjj
jqAg+6qOprWKmF063LOTmH4h+VB/JJzjPlo2cuAs7kTqtZegxOWgMh1xQ0lGPaYcFmIDC2cuZ6JH
cYgHjuSL5yqYlLifZoW0PwkvEpPjco7kQkeAqT2ALDgFSSLoPJ/5xCVOqHmjaDHWppMulyafbNU6
q786pI9HskjZDH0mkcQudOQX2ft/hTtDOMzsf243VnT3HTuoAKQM5QsGryDP2Pgx10XhMDrjVnjy
n/vspujFVsNKxSXTtebWrStrROeilj70tx9gCQ9nvrobjKJpyICDfTPdOiEGbE8+aMJwP9fmmBAp
ZoLtGpxXF+Jcj0C29lODobwXmcmeHr+u9uBl30yxnsm17alf9he0f01YxyhyPYwoBME3lx6W6jV/
/cSsG9m6vROSHF0amnIRB57cFq1B+eeluGbvup+YpSpZPdf0CzvYKaJ3lSdvS/qbwyQGB6juPg6R
OcmvtKEdBsuseR675hYYbvC74N8DGH8nA5Wlvx1Dh0AEamtACqD8oZ0axcpHkQZvGTlFA2NgL/Ox
GaPiKnfOIe6WDQOLL+vXdgScfNv1/bhz6kydeLbbcoB4tFYnroxGyysp3pjWg0ejG5jGt2Za3McD
fTsLkCPBUkOQvvnG3gQFfcqKJmqbuXbdsDe/iEl1Xq8mcKwwuMprtmxSeEIUkuBOr2s6RFUBPxL6
V4Cjr/1/b2cb20izmy92m92HSh5P0RRfzFuXChx5NfQ+cCpQCjz+qcIttEk0PUjb9nwE57ALG66T
k2p5reI8CxqpDli1vyj/nQW8QTMj1sunZlShAa0vfCWkUYN1rCpnO37rNbM025PMjMByIkpRu7hs
s4VmTMuYWkjdkCtMtrgtpC76Oxaai8RIe8Ob9kGu7M125d5xqLTeDV7MDDf1zuuFimJQt55Avra5
LSiuZUl4vhEI0cmHcs0XKRTqWZmNbuFmF7eSsciHSEOfjDeQ5ttdLJoNVNa3HjMfu2hiAt3LL4Kg
QMTdBSzkTJA1vD0k9TuEg3g6/hWpkwygRAkEarU/iOB7RHcK4lid8XHlNSOo2sCIBLs1dy7afgm3
ma0vGhs1yI4v9E2GuB9gwhqfQD87G3eVb/uum6NEqlWuftZbcDHDzKTt78bzsclWMZRwi+93AHan
RBlnKOWYD5vw65auOCd2rrqxuOMexdMt5PwcR4rJlIQ9ujxB/EKus/gJiyiQJ5V/AHNsExlyXg0q
AXEf4vEVIBHFqqrXAGeBMyy8q2B0hSzBcIaSajpPzwDVpBCqVyDJPX0F6hyM9qcXQ3OEajRUJE0R
XcHvT+qwG5M+2UB3S1XIGmz2GTkryZU5pUd913IUnvel6M3JvU+FkgnjMzWDIBX6Ns/zWFMIbV3Y
cQI+9Fj0RFkCMpbdWIDjgIs7ROW88dMzapPrv8lq7x4Mfm4vVnljFVYBKd+8xBK3vUAdo7ovgB7V
AvGo24cxjnXXNihKIZfAXZDHrmUBWnneuq6wcjUQLXyjElBofO0zo3Ixa9+slt4kgcAwzJ+fIVN8
2ImuZV+ywAyfbCjuL0LN1dxy7++n4iOQwm7LiTAMYKTm2uxqUNf/vL4xULKa0mOgUtz32r/Csrqe
wyqenWdJVjTQAh1u/9TenX2ktmGCrGcjdyhOknNrI5xYjkjQswHN2jUVFqS/RDj6L8M0KawEuYfd
32LnumeMd1cpDZ/OX216Zn7yFZLkGnp9MtqHw4t2Dw3x7XPwb+GuzQpIfTidRhH3OgPAzZgV8h0H
BIOP7XwxmUo2UMKf2sns4r690NlLFyQ7iI7D7mjN21YP1+E3tr1ncbIIOOskjbBzc4mFNNKlAkG5
IYKAd0mayVWaz3by0akrqHGhYMcPW6ZkpwYDJWozSKABBVL5VYmSH/zWQG4R5OXaIuXB7GxporV5
Y7UDq+/Fk6O7LXowO3pBt5j0BIP/bP0HY0qgFhAUnSsXgE11Q7WwqF11IJVMgtl/kicINYZjVlMU
wXkGwQ3HA4k/JNk3sTbS5zVeyoav+myZIzQ2jB9JjNh/SHR+SVaeXAtogw6tf5O6BcafXPlB5y8i
j5O/T7e4BDxZ9K+h/p2CEw2lPwTt91wV1S7VAD79tx2L+eLL8vC5CIa1RSOqeQb8ttG3WmZys+g5
YzLPk9eGxmPBuxjgSM53NIAznqdVWXAwKm7RPAbC9Mmf0HlPtvlslpqVZzNVyyoU361cJI5nWES2
S3u9GrKAgcP32kvZ6HP1xXhXUzreP6h41XCKsraLay9JZ1BMPWwwJsQDKRz7oQEj7zfShLQCJNhv
ssls5S8QM6adkm4xpL89kkL1wWBsEHkF9cOJFSvPFjYJXFosiuxjan502tXRkp5YpsdhheF0y/+C
8BoshtF5pIkdJb9s5p7uvEFPLax2K5HS6WJWoVU2M80cqmwtyB7UkzbzIiuSGNIs5qIYoWZXcKEa
bkR1yw0s1aQoZsQXuIqp+ylVjOJgSNGE4J31QFTovQja8Q1Hcp7Y28u1Q9+TpziPoCQdsqrdqRwh
DYVyzjSn0pb+23n1lkItRszx1rNL1rgvy7thdN3h95alNz7N954nMDdnKIZtMBH5qrGxjmFMWRyW
/H43hlx3SvotGxm3gx/XsMatZnh2wwEJvcJwmQDnp86vE5Zi0bUechIaG+cTyskNxljUNyOEUFz7
DKTBEwl7EqiU6DDYCbpSEV7fPDEeldMblDqNq37xcVXvmC+GPxD3P/wsWZE2CoIs4WEuDwu87JfW
4LUBxa+JNm2hPKkAXo/gHl+h2q9JOVJP/YEZrOO4ac9nWpmkzMKHPzUnxejRYDlYprz5+lv492f3
Z5IkvxMmNyXzHtzIdks+xrbGkEtESpCDo61weAIAMKbkIoAzReYkKkX3lKfy3tZlTbWD10bjzBXc
p84xcXMfcBH5cfsDCt+UNZ7NDZEasvFGBMjSjaO5kDu6KRI/XeIuD8c9K5NIoFrzz1kc7thTFb6c
axCRmxN5uRRRUQv5V5w6+V3FqInQtIGVpx3g8RG4QJB1H6lzO8/w1hB+v/YvXvcsrttqA0K/4TZw
cQ7hbBPHGXhvqhvd/xxeE5HdZDgwEhC9pdN3D+5YT0WJUy3uU3EaIWxY/mFltvm5/bVHyTDwxzLP
mbkiOMy/n0Tt/wCmhxK+zb4whhZ0Aqzd/sjZJvXiNlwMFnzp4poCPmCSocAYwlPfhsXIYuZp/zLc
LuVz8TA+x4mGToei5SX/TqHEOUmdHa7aPmznPYThIU7RlV/lS2sDUAuWLqk02le8yOsV79Tb880I
ipToER3h/eTigxCsvF9tVbu+uFcUhfqS6VkOvb+J1e4UKhi+V+T2/i3Y2g9k+IBR5PfkzKncipAt
FZaKfJnrfNl/65ztVXmvOURn0ncIJwBO0pRnzOKd17WfeacS7zYNkXKEWpS/T8wW2++1XU9NRG6p
b1+gnFHdYrg5hK1K2BVsMOMBtPiJf0UJUZn7AvF7cpqRcfdX9mYgI7St+bijOUJ2bfwLkce65ryW
E3EKRgOWhgILCRZcbWQCNCSA87w46TMuGiziOjRVW38Fz3tQ+mgi/IBx31CGYa2Wf0D0lGtci8dT
cRula3RfWL8p2Z43l2bqmy0T6hV0h7QF8xpCeYDE/f/+fRJ9QG1g2MQ9QPnluggU7Ph7eNQAvxdI
RphgeDz7PYKKOcFyHL0HB/eP68iOcLMIF1Nv4DiUQEA7Z2LSMciAhFgmypPnDjoI2pgXuhi1V5E1
lVjDMC/WrYaOdvuWK7tG206FEMZU4vXifc8PUGI7eWorAjAObX01vxFBDBtSL2Kd2PsIHLbw81WB
KbO52qWWdKrOo6bxmNKSQomxiGyDDQq48U3iosKYOTuDUclrCh1xtlvjrBhvkG4QkVuvlbkdZ/2r
M1bsHTRIX+WbjbD2POEW7Rl/84B359qTfX8CtKDqid1QwvBmx54vX+MCanV4Ir41Cq0uL2HeqoJD
e4d2TCjkHmgSJizm8s1Bdhd59zOfBSwYjZadItkVnbJDtW6L+1vlUgsq0u0Uj0QcsRuQtWIaAbmT
RiaS1W9A5PgKU9QPWAblrTqfgTBr8OuyWCHh+TrHra/Yk/YYtxhEwWS2D82dS27TYtkOC7Iqvg2S
+pxXfWZYOca/Y/QmMcYlIzVefNIzywttz7JwRVm4VQ1Vi5DyLKe0NCkdmTm6sUn24+LmfQs1Xa2q
N6dtzSSWAfigNC913+bOF4S4DDNVFqdq3xs3ztQCbQB5MNJwpC7mmKaoqlrRAUN9vJUsQ04XWUG4
PdR5a+fvMJSMgT5in8SWqhavD+mjwDij7rKmEB98oBhSQKugca0W+55QsCC4ODavCk0Pw/CtfFo+
kkfoECs63VrEpiFW0aKGDpKo3I/qiASK8J9bDWGbNhEQ7bzek4ywlv+hHwKqcBN5vIcVM+2azPt/
kJgQc2SGElin+0w7LYk5SzGlfq3BjwRSU6UKte0OYsyBF6VCy885m6IGH+onXsKAubuBQ0/RgesH
bSAxeFHU/fncYRIyBmRLOMS7P4nVULmu/slqWwKEZuN53sDwZJFv13iIrnfSo2qUF2dUmQAU9pVc
YW6jLvIYHF/99nsfn4zaBjw/IMf/EQ0tjUpcVvvovIMeHCHJ0hhd3hV66dhvCaBodVuE5SWKhHNd
OX3CVnm8h2xHay2H47aga7pzQiKcODyJq8AD3PHseuqBdi8i/dw+Uu6W4hqkCon4P9SLUqUh3GYx
35xpK2rPzgjKXNeJxioaGrc+SnOqBnT4hZch3K+fhUXFXdjEGHM66lHJUPqHxgI6caqujq1FvZIB
kytCLzQ+PyxryHJ0Wjrc+w6finWqWTJaOOgRGVmgxHKyRRR6UYELwuELLhXQ7pUkTOGAUB2GFr7A
Gjql8xuq4LXK0Yf3wr9HT+OOrrhQLax9Z1RlVySgQgdjdbPKptkdKlUhDYSP8NBy3QjgUhGxJslD
sMR+QEJxbA7jvK3v9Z+pA62VINgoV0GmNyPnxG06f4uoYm1y6rw4AM3WkBqQtMcFBupcer7XcgEW
fa32HlwwyiCPShtQHjgnkl3MTlcFNkjm5+E0ARjSGG7mKtNFDOUoVq8ZbRtFV9k7ouo7oKO5BryY
DA11STuPLgLiOx6lOvGUQrGhwany7fFYAR0YN5JKyXPGs0psHY7avee0ByFQUEOY51JNuvKT2SbE
5QBytYrB9oveflBDUjHvFAE+X/tBOHEB1RqNP1bF/oMmBBX/fQMVdy3FtPjYv71ldc5lVH3HdEho
awiJACEVqY40xrf8013/pIzkjw1ZLWVSAoSIo4y84wy4Sl8+Tllee5yQfRjGaQSK0KDgZK2a3hVw
z7hD1RDhxE+abzj5kiDR40ebb0hoZ8gSCoRjAP4tdKj1jpVVZvK29A3HMiPppKBVbl1eZIdytzAp
b9QBCasvGT0AeweGSAOo9lDZOaQNDBnICHO3tfb9kGlVfxJDUTwvP6m1j62vXvetnvjuXTKLwFc8
IGiLugzcjpYcyvIh9oFAZx2Civ3YAgcPl8alPkPjquuZpEbm4+et1+x8o9k+sX9xo9j7E371LpWO
pYZpHSx0GsKsab9EHqVsGPvf1ozDsS99i4MCnKq9tXIblBim42epICS6FL2nAuZIl/p4PErznCj+
L2WrunjsPIba0sAXpQ8BjrGItwSQ4aQge6z/fC1qI/k5kfEtZ+bL7Mqh94LSZ5BFWq1SjZp4ZObL
h+8ZqmRreLWzcllL65Ym+dvIEGa2JEEpY4lXfbVJS83nhw1q9vhwXvWkBmXnuY9NaXYXCzZwQC7F
n6EAuZGrqIyJTFXlJ3SVD7VW9ccDK1ulSEkePQ9kx3wf3SbrhzAkXoSoin1vPDk1LAB7qYEm6LiV
DUyg7/4Qrv7qFDgA0noYlnZU7kRqoaYw4DzrcXjUjv0ubg2ijgqQbpku4q4yf/FaOlwPDBIpwn4D
cFNZad2ul9ZNHoHpUrkhI6dFMCMIcXnvb1riIit1jiosNGSPGd7dn2Mnqy5gGWYxBv++67H1Ohcc
P5VMv1OLrnnBYD15AJ+fG8WOVhLVpiFGsRz21qOhAM/ibYnMxMzQdCaErj0YRJnbu+i+Wvw2yYpP
w6HCbCiBeROxAwTGs0UfsdfL++g1RumH+NA4jO8I7BT5DG0SeGCmPi2SKz7nSR2g1U6llVHNCaq0
or6+CMsbhW8WoAVLJjqHROOu2rq8bZjdy7PjrtEsmTWL7h61kHVcOpsPwr3T4cajSgi5A75kga5N
sKeBOUvTIdttPJxpbg8ee4cLIi0rlLmedSYlRFZgS0G0S/Z83hcAzpK+xlioTWP6HbvnFdW1CJPG
NXH8ziY3moKf8qAkkXWANXSNABJ3abyYEt62Ge7Qt5Aw915sav6eHzVda3iPydodt+he9M+3jdqJ
eefOpC3438AIVruQ/Kf1kje9lLaZMWp+WwEeXygvqBJJ5M2AIBBmrl2RaZgkfNbG6Qt1ivm0mtPX
aqNu2z6hv3SRJDbgPfur9mq5boYDe2BqC5v24wEOWXJ2+ie3JPhVznreyIfeLKYb9DYHYvZNOxMT
5qVaNJ2RswxQde4tKS7BnsXFK5UHFtTohqT/PSoJI76lDbpZ/M2fx4r2vmn4PL9/cYXRpEXC9jbb
3ORji9ZoCS7w7zEvWw0IHSvRkGs1rkb0weNUsseO2/C0irLfjmt0sFyD11QMBzUinztBEoHX4b5P
2YfiNe1aluokQg2Vmdr17eDLL+o20+V3MsSYbwcHGEssOK+XlTV7+uKEuKKQ4Ie+xc+2SW1I5b4h
Ao+AV02145/JzJWe4D6C7zUNvIsP6mbn9i2iOYY3rIy7N0nitOY/0y59XoEVyxNjw/T06OlHVgWJ
sHO3rNOIFgKQZXKocbKdt1J6MnCxCZAQMaCGQ18XKvSkKkwNdfEgQ8k9MjzFYfjSkcwPWa1yesQ/
CtiTAd9jjxv0+yEOLgJLq+BPKMKnOaSNGn0o5U82C0bXizqfC+XEFvs9tuLpyc6cbApsGHDhE4vg
8vZDKvgEHjLrZmyXKLw0S9TqQUssA74MPMaZzY2CBO5ufLtu4ePib9xys3yajrikfvZRorZlsbZI
sG2KT4nJ8vNlWbTtf7rrXtlN8X11erLflGfBATXdTWWLEh3TFx7pGrMiMnnMImzPf+fUkLNCjouF
lb+YpzpyhCyE5jb5jAvV3uC9cDFavxxBR0AkdyynaGRwroJZOtpCfXTbrEaz1NAtvT6VPrDnklgb
R/4PbGul1vDzDC6bPzunchd1oq8KgQM+7RA6sCabu4YOEXKbfl5L71WkSTa/AhAg/Zhpi3tpniLz
Vp1pb6GUJ980QVBW/5YIoIYLTBDTOjGWQBmsZBP2tO7D4fGgkSyq2Zn0bJ3+3Dz9DWXWxcuVfoEb
86s8BhiuS6IeUENYVa/qPhUsMNVla3c060T/Zvv9Jfy7WbFCtdhsuVxmO8zNyBPUK4w+Tf2Uy1hG
8B+fBbCH4ScUxUpspum/WN9ESRark+IW/7qjRd4rrg2ipjnM5O31IOsKujf9izIrWOV1/1oZ0GNY
WTgvF8lfhPdGPn8+W24IwQ7Xzn5REWLOIi7Y8y1xHPUcQ87pUDj6ABKIRz3V/hbfUzn+L4mhW1KF
OZ+fjDcXE0lnIaYnzLllrsIkrT27GGdZxwRFfZB+cHkrLQIiUHU4pNbpAYuCpIRElwBXG1hheb7a
7UYml3LVgVZnmYJceQcNH6h5nadG0LSisgcscDKA2W5vLAXRzakka1rk6HNIh5ihNoUfp16HX60q
y3ZUccY95JuwLStV7dcAsDIZpTwuKwoLq3HQj9qPnFZO2WrxJVIAxzqFMFSWCtwUxyRJA02Erc6u
9kIiK41MJmNmoTaF+OUDuGpp4XFOB2YD3o020MLcT0fedlf3q/5n/PdgAiNDGn8ugz559jEG1DUg
gAtsd5Vjb3DEW0qqYek9wFwSw0cQAVfows3cVm+m9REn/RgcnuuxG4F6MwtNEMvYgROKVx/KN95X
XBhJonVaFELvNgCxEPOgJEPQBiKdJCVEqpfz05LSLNkR6tiWYNOrertqaFM7z5lU0VS8kmOZilYb
FPwWC49KeB8svdUTE1A3nZyRIGBmtqgmRzKosXZoGUSdn3u+FbBzEKSsa4LMadkaaqDjBwnwE2od
39/8BUunmMoSG7EHFdisVQFIOYf3l7bwbLuhRX1o3EgTvi2pddpYhkBA3tDlU1r4u4J97KSztpex
pv3bRSvoYHzGYMnMPJHoKWpf0f57hZLnyawxWAoM3Qqo89EcIHehMSlv8lS5vIO/FptKMgUXjWPt
inJKyk+9g+m894PzVtiFLEfAbh3ySZarspJ/pEQ1J1psrc1zNA07pQCEC9ZdgrKoK4PvuHhWvYbd
/uAod/xRj/wiHN749+RKw62NiGcm12msKpiWVDcuYM1RdEHZqs2OA0HDHUdlrQRZ2W574syeWb3O
74SNj3QG4ly0r+bam1CjlC3FXlwV5ca1QkS+GVCoOVB658J3fDgK966vk7z7nrmmr1Jgq0b2seEk
9PAh2F2qQ8FYOfMJbqccj/3la1acpqB3WQ1zlQXXIt0v6qdGZK7RfbhF1yQyFuEA0gW2lBnhV8sG
XAX23X+ZmqvOclPKRZuijnFFOEnvn24Y7xeFROMlziLx7s8jyqn6Ip9e2vMAOsY2lM0b/fBSddTB
B3Hxel0oAyY9P4EXcauju7eVFUhK3/JDymdaiRjy1jxqFclSbTx66zgUqYRHyW6y02hIQjvG+apx
YUlJ38wpU28GN2Djz8Fg7/L7mHQUiO1E+5P+0eNt7mAtiBtGmX6ubF3irX6bVe767b7mL7GlcJT1
GiqAuI99iHi0T8f/LaknQgzut1eptzFU8S4X3JBJoYiHYOtU/IiNOGieUiEpsXOE2RmxZMKUyxz7
RpVfIkaP/g5mGIJJP0WVIq8g0az/S1u5Cnl6M+c8ICwPYICru0hw1Q1s14ap7r7C7M7k7mwsc9pi
i7XpO71UvdIjiClSoUX6/SJ5ekH5v6Teif2VQrIDk/+2AkObK5UJTH0JaYg/F6o5+khIzY2gb6Q6
rLP4u0ktck/VGc9LQUwmsp6Npr3zdkV9BCIREe3lexunmnCOe9owb2r8ohuBAZr9iFYWxDYlfWdB
Xdx4Xj+pl/4FjY477q7wjWxovOh/zTgAD/0mQazhi21m9gRktc29K+HyAxdTwIWhjH4hqLqy4poK
lqhpyPmQwjowt0TZkgANFQ3kpdYXfqFr+c6rn56RGZGg3HLXYzPvLO0j0T6vmVkip+3pnSQKMrNP
cqG9ilyKuCANrJ31AfptynWAXRXE33+jwzb94v/+5KPWNQn3lf2r88s8qraLY5Mp3ch/D3wQUpXj
VzGWTxd/CVgvPXgqrr4Ujs5rkusAVQ3Jl22M/kTlxz0rn7LrS01WTkl3wg7AKPQt1DaZbTeWtBAW
Pr2QLcoTXhuATrUqh7NbU3jK6qcqB3SSBo9TLMICLo5NvAbHzeM9Nn01ovO0a7dJ+Y4XBmTPjhUY
Uw7VybDNRlkJP6L4z9/Ko5KFx50A+cwcDu6ofjde1NFIOMWAolHRnqKIlGEJS+Wkhs5+AcdDctbl
6IOjPMAJmnj+792hXgFP2tzyhjGqeFqCQkikHdylM2zScyPKdQgT81b7V21Em6UXHtOTsIVYyn+S
y/3OoHemLZgGrsJFNviIOxbhVSeWt/Lj2kdx60t4RpmJk++UIJwjhTySkNixOVHchgT3eUjCApSz
Wg+Ejfv7HLppaPuzOV2PT6Ihhhr1fEWRjVzTbfY2yM1eRuaO00+flD6AuMGg0TSxfiBgl59A6YLl
E4S50BRLWYhl8+Py70dJW91Jyz/C2ExEba7jHHH6xQB+/4Lr/qLXPx5nJlxAgngSToTB6stWE820
aJcYZu5c15iQM2HTx0PQPTPXEmNDf5ZcZ2PbWf06v6uNXXwT/NFYXKsjZ5YZzZXbKT1Cgr4BFgYa
91kvzQneqsixM0HT408X9TCRwkZSHLMivf2PzDqN8X3MQl9nssjuevEi8sEbzxdbGi3vjp5YAqP9
XIfLSpHcWZEm1upNh7C5eT/t5gMpPD+1iFhDPR0vFxA1250/ZdrUC9Mea/gzP7fUedLOlppMVV9J
Bmc8dHj0wUeKmeIv+xJfE6WSZxjS8OHbHMOGawMHD4DxH5i/v1sQ8aCk22yVTtxvObe8/bmTXEEB
Wre2V+Q2svC9zLUF0srq6gSDFDm+s7q7WcHjbbcBhv7QEoVh3gODlcg1LDdJTmQfHdAL7oR13IIT
TjRRCjyZHcYnL1JAgYlOIxmfa4LOXsrvOOmRB5XlJ+43ERkfpK6rXJ0qEo0piEH3BZiyCR3JCbMr
zomT7XwzdPOE7TSTG6EJGLBTSPIZnI6ZqWS+GSux4x+632+Bt0hACfnAYQe/m4FTtdcSglGh6dFM
RbbxwcjPqjnL+uTbAdAyVaHAgqeMpLlhetr8jYOD1RXFNNnQHtU0w2DOrS45Ecgt/9+gI85vYhQx
M5ZixtP0/1RKF4hVkkUJ3fW/UvW9dTSwOpl4029kvkxaxEefZ4KyB0u27sikqGmNMU1RshulwpWW
4aaNC2o37UF+CSYVNft1Zt8iFjZw60/Lg79L75Z7EhKoOeh6Dgwd1xe2FlYC0+PqreO/Zo34z64K
TeulEKaY+gUI+M689dG3y6PefWNgGcuLgfF0Wt7IeXBku3yzW7dBQKFYFS+rRyHn1BtcyJF9A/ns
ODHB6qbWsLCRCHFf3KkH0sZHsv4Eyg0RPcLp8YP2heNKrSTiplcIcLEbFWpQGZu2wWBz8EdCF+3J
XUfvY5eAoj5Dx1uz+FWuDp0VFuUPAOq/zkBtQ4usDXEUSp9fqql5wmaxLz0Uumoxt/Lften7lQxA
xzuPpm/7utw7fHy6z9bCSv07OHHKCUWuHYMi8680ymYABEiueJIPHxqS9PWytSxj5Dbg2LZisujt
XI6bpD73SAehbZQ7bkaIm8JYOkxGBAcU0YMfbEAXtvB7myIFLktLIHyYzv8Fk2TJo94h2/iYwrIf
6NeFoBNfLeh0XnQZvAO7jMe4pW2yMydUfuYrlCppMGCwOAeeI2hXiUbkjCc0QW6e92e51eJFfLHH
EnPKSmf7pJ4u1Ti1ZJODKcuN12+At5w9yXFVpfbMh0kW7ygkvG4JYuiwfU67gcBVzwIMcmQv1xZ4
erhZtgzhMtSvDLJ7rPo1n7UWfqkwcHRpdGvTYxWAMWwVehfdp44+fl0FfBe7+naXjqjWIIqG9Z/x
7LX42hJQsvpPyK9GIynpAJ7pjbW8GcYv8NU8skyFaxwW+MjC4nQrRktRX1a0uy1yWGCgC3l12jZe
CSls+PymLUfLKcQ4xHvn+fGuqP193cCRDAwx/BLQgk3J63XG13CDQ9sRCo8Ajs5XquDHDgEktsyH
z7iTET4XdxPwUrJA9IqDYJRL1HyEoCBTx+nEEj99qmqT7L4AiSKSgzD9h5l/NRebJc6b63Q2o0hq
v8AxKTziU2veAeMeGJ0MNL4nIZRq6p1Xyp+AIHhgQBC6FXbB66SjzETp6yBdDHSK9JpYKoSGQFwK
ajay3dWm1WXBHHj+f8oBYWiAoJz4FQSk/DmnlrdPqYg14+IvYdg2YaPy20bnDYTQwX/wsM2mSSel
5sSwDWHlbIZZa3hLfxj2w5TzRsOwirRIt5VE4nx3Au9Tv4f4o3AYsnE7SZANMfqW1Fxv2LsKNTwb
N52LLfp2K8WyTsfPUCmrQfkoE2mNbD4SRSJVvLfmeEYnsCLHBHwwt83WibhnmQ9D+EY0b7zdZ8AR
3jTJ+8k7cFc3VMeg2cFIsjNpQ+2nc2hLDox+tYjRCngTPMGup7JCraCpOEiLoKvKIwRTv1i0PycM
yeudJthY8e5TokpSoQAUU5EjK0AaqUWJ9BZPr2OKB157fwOB74tmesr3weZWjypVOYiAL5PZ631z
YTF9mS5FBM5gyg4j7wRo1jTwDCLIXoiGyHslNxdM29e4v3RsCJmZ0fY5jPZ5J6XVyfvCQnLdH3ib
rQ71P2u9Bp68GpiY0LBhWqaKF9QSdjm6sTDtUSriGM1mjX9PFFFen4LsV/Jsr9QDYYmHAwi5ZUqQ
YLvP3IoHxDw4/TIojLoc4JuTFvPpn7cEOl83xSrhY1DnXmE8vqkZs+Vh19lw3awPZB0iT9QRiBqZ
C+jAIoZxMLd1dcnWSV2N/XQlIj9r129RLPg8ojOyBnGtyMMzmLIUmLEnIHzS5pMUCEnHE4S5bEf2
yp1UvbjE/DadGc+++wKSKx9eYTeRBJmPuOfpKex09V2qG4WvsdqDXblIPNNskikXYBaVO2MgUBlQ
G54/vO/9WJjd2TpuO/k6CmXvtxDZ/XjAoe4BgypDtPFqv+9P+MQg5s+1vKOaSvi0vEVh/jwqTh2H
IRRXQMFUgRnkb/H8Q8jpz3xr7fSl5MwxzzOihSgL1g9eVmdDRax/DhmasjkJCXMd7lOb1RUseWDT
j++/BLFQu8mAYqcNf8GOpQydnXTZZD+oZRGmTFsYtxIqdsXE89uNPpKTPzZxyMLASApPJoXTuKTU
3uNLh40jC4gwscKStUSWov53Qm13Zy83ZXnyKt6zDRABiPfTXZQDxpuwLyh/tzv0rIQs5i1OqUSq
DuPP77Q04LUcqgA4V9LXVUAvnweJR2V9yYjwSAsFqn2yUZevUsMm9GpgZ9ZXwli8/+WROr/b8F7q
61YcYGEX00Z4EigMUfSfd9/jAuPGy6MmE63/mU7eE+UgeVmi9kEBmFqrkvndmnmkIfY9lncl4E2s
rXS+8vjSB6n87ez5sz1LCW95p5HNoVtDnxhW5Zz6BfSDu+J4wz/if+5d8RG463ElLdkTw5pVxDfp
3pMzlFMiFTcwxFTMgvUQUHEJd6eidBrzEXgnnUKSMdTKAfc7WxHyVQLxbjpJSdd810DNHWsrlDT4
GSdAK6h5qyl1uPTlWRDYQP+l0hUezIZT0uavIRZ3QAnUfUgWM2SP+yV0nqEEcjYY32EYJiUyRHde
bAYBQ2ttG5qPK1ZWuOqkufjo9EXKvaCmKYTVBkCywC+j4dU7g6svbyqgADUBDbf1XVdAYS4VZRPc
fWNM8RhIWUHiXPqpvoZUmBpSseBHFNWU7OHij1WeSw82IeB5r3Dc8MhCl38ffDy0jLui2SS2rNiL
CaacA0e5eW5Sa9q8L41FODzCRyYERZuhCTjcBzF3oouz/Qe1K2wiWuxTAIIBtgFAdeX0rAMZLpC6
x8h1TGLQRdDeCZPEOk3zTjA2e49HhPNI7N+oGjjNsVPRpX5V/1NQTaE0UIUwnMzZhhBjubzmg1nO
eTpugwmI3HNzG9mW7ekV8VTe/W6HvfUqvo5AsDEnDYEMgNTNMXzQPyOA3MJ2uiCr/O/2x5D4EW8h
kKIDMbwYhJO8DZJS9cO0CrmSm6DPhFuoB5H8OIX4JApzyaqIRJeWawLT6RWM/OtRY6NRFieuJdMX
nb4Ih/3ElsWknHboq1sWSCZ/r7c5cz7A8Mpre+8cEx/BkY+PEzg84mZalQ/VJsPmrSzyIsoKeiwJ
cW5xUtexqBN7HBeYkaLHMktVsRS4LkXi2Nor4KCsVtt5VCqO4DhHq+30vnh7WRveEmNKx2/hTXdL
Ls79A/ENv/RGjPfewDmBVQ+G8wk7cQrAt1c1PqjljrQQ7pIIMRRvz7DBB+x3RLT8IGHoRQfrpCKS
b87XGlqOPpJs1ZK4vgKZPyhafjYyQmhQE4tjoSlYOOkYRUhYjP7iTBCvQ7DhXtEK7CE2bLfyk30H
QsV1lKYb5ewk7oNo8l2rhkXVlO5CohMO9RhrEpRPvY8CWaNRrqXgwRUZTWDTvxLcAHhK8HjnsapW
RcCTFcTjZEI+QY2rcwN3BQgbiXqVi9EO5j6TBGhb0SWjll57WaMmjhT2lVnsxZOmYG3AtGNj7Tx4
9pfpf0wd44jjclZlVlqUudWW1enQ28eGApodiesmNzwS1rMwdHbU0+gTfyKIzhPe4bkzEFuEE2fn
yEdgztdXQj+bmt3iEGZUfxJ4bbN6AkCyNausHMhlNCP/EGetg1g1vt7v5foLUUUuIKofGSlKyxUG
pVClosWNY+nex4m68taOzYGKprNZT9D0CAjz2VGJ005dFUV0XTSHlfE+/rA/xbB4db4lxfmkzc2J
Xq0ejcG4R+NMG+INe7UyQ6r68dBKLUSgl1jVZ0jWNB0VKd9HHnms9SbTaFMkpdhvESWiI63wTcJe
J0B4SoZf8RalNpgSIKNi40jjvo9HwfBRbQMMdNTT6rAFaLwy6iiFD/3zS9e2qlF2k6xRait6E5Et
9OY7w5kNsMdQPXab/4PIGtnyZoBTuDBeZYme+72KaX4Cyh8vnmHP20IQ5ejGruHbWUibmZA7ZjK/
CtfHFBvfzRcABtX1YKbyzMZKKkIQbI96w5M4zicE/yQAxVWKf/riWSVCyn+7IHPPgBku1xf8Shk0
Xe9O02SaOlooWWlVMuw/5uQz5k5hreDoTciNbYOYMDemeI5PWARGGnKuAVXlggadYd43Dwne6UDK
/fFx9WeJE9J24HjXrnhvMfYj5QA49p/2/K0V/du1igMtMumZF1YtGOezKN1HfFLL5zNBDMIgNF2Y
kXHxN5awABXM29P5jx3GjuACv2mm5y5TJaI0avfoF0VStrHD9hiMI7277Ma368ETlpTwP/VKGMMw
xf3jfj5O+JFxPK+E7N3WExMQ3Ufll08161J6Jp3qFvZuxLn0Ragsi5PcTMtTVKWvF2+kFkVUEHGi
kEU7hJk9Tne7fpUhOBxMHNCnJQ6Hr1dXGuLy+22RFXQoYsviF5pkZmhFycdcbZTFuJNkwM2/IWKS
uEMh8a/t0kpUUIaKWQzSG/mpDPXtbRC9XM2M6GTyyoY4DqygoLJvY5rGuTSlw/bWIwrHD9/57RAq
BMG04pqBojhqX0K8CKL4WnsVF9Nk3qdpe5PQrQDde/EXoHfAlK2MWgFaZiv412qIdfScfTs9IF4w
AU0vfhpck4IJ773ibZ4THzI6LKSb/oedEyidRFQzalfZnwdXBv5nnwUcnS/Rk1kvjuABy81xo4TS
ms+cJHsq9A2y3kSLpxSQ69tF3vVI8fqp2zuI7aGvGJKg15TJj+kGJQk8+lOtk2+nZ3j5FbCHH9nH
P7gOZhv0r0G8mGRMDbDRQJpnZ7CBSqInwqETHVNhmX3354DLDvLLHxJ/7f5ybssHAPRcmduKFYDo
zPDhsQokF3tPv1+taf1rkyL0m7u+hUdJDdKzCS2ZA5rg7XvrNzlY55yK9MoNMEDHran8ErpeX954
yfYINpOB/kls2JKw+y4amak62yCzMecHzBAj19yi5lVtFX03Z/Svf2m71to6TfBjvObwuLXluO81
hnXur2eA3WrPdpKAM3gpNz/parIYtPxan/7iOCZnpN6aGnVSIne4bDzVWW4bhPcGc4kRV28YWNdp
xnZw0V2lZbwHLYhaRsV4174VN/VCcEk4e9dv5wy5s/6YTcVBwvp67lYNGEjOiB7arRB0Iw9wznHu
wa/PNRv951FdTRgAh4fH1OhG60HmWQ4/VIv52UWNqdhoiKglgqEdu35C5N2NLF2mvyqwzrzZ4QF3
9o95uSnA7Ek7GihNfQWgrfYn9XrSUR2EZzPjFgsu9cIi3mxFlczxty5/pzzyocTlOuEzgmYt1nLl
tE0xiyXFCscP6IoSRVevkhzFwCpkbNQffFfckkXyC3aWfzVt/OPihtAv5iixex9Dz4q1BSYvvEa9
4y7403z/0fpMyxS/GGTGZJhBBRWXGWufv/1sT/ZEnjBlbcRL5Q3CW+kKpftWj0Pa6yWoUMYBktHb
wrFomBYLyTkQHouZc8WRqVXb/vjFijI+EvPz23WnqNscTDrRtv0QJyrwX6yWteBq/s3xqT6zlUvl
wHPwsOJvaarNq/oybOjesNLTSEhQpbMSMqyKMto+xrPvc9JnGLyOKGlXscdg/51YwTjrJWr+3Oa2
LwGSNjnLrqtd/4KCGfcTtStxtTBgYNip25glIU24WXS6B9vyIa2VKCIqNhZbFxoknK/Bs1WOUH1A
AmHmK54RRDz2R2SXQHY7cCJzapQt50o6HV6lIBlSewXgLB5jsz7uWieD+l6cSdBTfjxzIs/PoQcr
ysMRQG0U4qOwrsL8qksnKNfBvn/IgibHjqCqn3Z3Zys+NRjuuP2hR7EZn2dxUb+CUA0bHD67oYsz
krGXlJ4lJVhcX6IiMoJDC+02R/Vsoy78a5Whn8TEGcAXoS81p/2nsp52eBkKdTWTmxYvs9h6Wxgg
Ga7gNJzK7Gk9vsp3wgUR1e7g5OIG2zvYu8zHX3tkxIYf9qG9cVDE9eIORNl8Bf6/roWtctBzP34V
iH+R7Lmr5pggYsEyNXrxBYVj0gUyI26UGSScaT73g5GbIhPe4bAjf5UgSa2ua2cTL1n6cRWExCao
CeaqCG5RUKrR2RmVwaYn7brga3D4CfnChOPIwu7NH82f0dPizT3T7PowtKpEBCaRbDlP2Y5D71Zw
GQQ6HaB3+38I5RNZWwsJ/xuuG4DO9fQMms5deQkN5OvCIZpLD+BgkP7YtD06qAyQgCzBig7b23By
q7HXmYh/EPuEPBTQOI10CXQkTjJQGD3cVhUFMDENyZz3YK3HaUvhWpdddHhBFk0MYpeb6jF6tG1s
1SY9auMmzEuImxyEQTraOyiOEPU0BmIR6OuNQiuKp3fowQ9po6VmGkcdAxg8cvCF1L+6oZlf75x0
+Znzc/zvu/uTW9+8Sa9uazUSmuumxKe4Ivx7ASlTX0/13OZiLjsE33I0aYLUwouNZ2ljidVw/f06
8i85fImU2CkAz49B4menTDSmUgDIzlxqf1EtSnj2V95Upk3wl8zKos2vK4rKmgrBh0wk6/2s0xyD
2bEKvqE08YjTqeWU8b/3cI4/B0pmQj77ugZSK57G6ReuQ5GHYDl7V/8iidAQ5CVimiHtz31vGjlC
d15Pja7kCmv6vAd1FS84WK/DznrVloscS0Lc89HqcH3H+TaP76PXSrchZ6vnKukato96Ezl6fuIR
3Au8MtQY/k3oeJoD2mRaybjbatysXx6Wecq68MAYhCiMERtn/T0TdXLIErdgAe4zBuusYzpp3WLM
T/78OhNqiG1TZPakB4MbWKlxUS9fj0rfp9xddy5y4L/zvINHpkZa/ndQ4hEj3mLA3HsMMWsewYhM
lQ9hK/ej6BvVCpcJF+zz0M2K5V7CoGb376Z0T42HHs1ddnuzYsj4kBl5nmmXxbKclTUJM6Fi7xuk
0XB6UsckrRvQXmVY3QPst/WfyGOLaN1KW7Zjzu+cmbkeDvUtzigfWuUNYdc/0ScEdugIr0X8hAM0
B1n1BOL/T5OsbAzTsOCn4D2GipXe/0PK+z7HVH7x13misrLlrriyzYfOl0uQbr4fTfTp6nepKQmk
gWeTdknxdNqwycEdjcS+D0fbXVYh3fRBVnG0rOUELkPA6YU/emNqIom1x6/AFs+5m9CXSfvLV8pP
RQhi4txeFPmfB41eGB462FaeaInfHI7+fgIbzCxr45UQSm6GFn1w35OflGJ/La5w82BCJSMo+Kei
zl1yHWaaiyEc6qfw3TnCwT3YL/tNeGQb5/LTDm/Gg3lJr48OOuO1M66emtk725Jp7BqtF0ZmB/cb
Nhh3/YFIbVitGMd717TmnydYrdd+ugVDy2jSInsSC3KyxSDPBbWbAbzj8jJJU913NgfZgSdlkF7W
pWwV9vZCNlP6WSxgCd6D1lIc3+5meNtbaRV77pgbK7FXTj+w1RBd9u7RIy03nSaaan6Cq0+38vrA
LbXcgGRGtO2n16u7I/jBzae79XmSFe0eS8E3ecHEBwerLzUchR3UngeH7eyP+6eMBXMR5spM35xa
kNSYpuTSaRfPCq8AZmOYyBUU+1J0pLN3DHD1zTt8bB8oBNqE1KuNaUZ9frZ87CBL03KEBezSNBEZ
rAdVShi785CdgfdhBZPw9fRYJBLtokxj5xRKyBbHg7f6AvulHYNyl09bZr/+ANyq537Z3x8WHdyY
SbVfuso9ZRVfLSeMAPzYEUAqDx7EZP3d5Xr+7/96YxbC/5ZFLTijG5LGmUHRMgn3g37kW0oMAmmr
HdoKzLV3Z+bntw0NwhLGzvWrf2h0VzfgCeiLnUrW+/HVoaB2SeXAP1ZG1dFt1NIVyXGcIxUO4mOD
XgDnoHoCKKYsSA3FeiYJ9+hFmylgejXthG/5Q/D36ZarutYrqYQrzD8rz1rpeMPi/RntIONZI5Zs
C+28xXBTPwocBeg8xlo3QlHLjgCVYYB4BhSSmsc6t3ROANfaRk3o3g2Nuj78OJXWk/uElfmKyP+9
jNiLScbTBU6gMPa03CdrRstYol10fE8ZwLIEjEhioSVTtRpJHRFqfl9rXp21VRKDvZl+1UK8y1MK
Bg+lKopqr5P7dBzH6XdP+DsFSahzjSbkxnr0Pkow6MMksCct/eYuChbyeplVJlhoyG69jLmx9fBq
AUudzZn6sVpiqEaHFk5wmRpL+0HGD4uEgK/MYjQwE2mApj1uF+ROhRqbpKSrAquIUQNz8PNTv6GU
Pk3jiFZtxI8nqH5nK90RpOCm972a1fw2o1+jaj2ySsL/uISjAppgJ7cL7c5DLFuzyieifmd4Sw0M
nIp+OHH8R1ZXiBXZC4RwTWIEKrmy0SuHuz1/wxwGJgv6HcW4uK44ShxWoG4xwEDXCEU2wFbGnC39
BuZLO/Rf19Y3NFokAyWD0oS9qoyyX16m+dUlb+/wXNOrJAEfBdTj82NGItNWm8mDnxEKhXI8Gzsm
M9IWkxfg8lWnntuk+qG+Gistg1KtTvqv0P55Ls83HqUqBRZDXZUS5ddiBlvsF2Sli4x6rEtlv2EB
KFNPA8osD0VOHb1fUfXrItw5qGUSRcFG+djZcMiu4pSh6UJbBSPNmGoUpWE4fbp4NY906F2gA0WR
ZZY06QpeCjX73UYymfgm61lqw+3AGMk3/JuTv9yGT/YWwVRgXdUjvgB4cP2JaeStWt0sM2en3m8z
J1H9oO0sfk2Go+TONofU3cT1KjZYSC8XExDDa9QQjcooHJQn3V4lzReNRVRSAbqyGpKdSVzz776Z
a9AS5ogpT+pgAjEy/xRyedy+KFY6/+rGfZF6gqASOWRn5vF92AQlxOYTZOx9fdNUmNiaY8i5osdh
ijn/J7R7Tdn1qHLWegls97gAzX1weU6cbmIrr1M+d0cZq3KIlI0surNvCwocSizHuxMPovoFfNz7
g0rd00DJBoRmTf7rXWhSPHqW2JnV0KLQxzYu0d13m6+vpMAGYWsJG1sK+MlCLT4ndv7JGzC0WGVp
1DzmecLHzx7rgtBPq185cI5QPK+HAN1JItk0EhYDNeBy0iSwd8H+9NnqiA8t2JdfC+RnGWNgW+to
eRCwvNwSaXMXIQzBfRfBr83YJGCNf0OjcMQ9YoMVDTG7ItWAsj5fRP7jLo+kGj9OoZQJcNu7KLjG
CQ2yNir9M6H621s1jGqSfWWFvHt8HeFGwcrnr9T1pq5ruoA2ETUqPHSPODBzdRZ/7UYVqdJvYAm4
kFGY2v8ODeN3u6budOOPt+ZlEhXfPAKfrRJvA3ZhGpoJMkSHViZyvxWc3yfGuLyOqLXq6cCT0kdM
RjfKaZq6BYPqpSFXXihouimGubXmBoeWlJtwdnbaNA/4yhZtH0X3Wmmi4KNpbng/WU53kRTlZcZD
e/nt/aF6Dn40hW6nhXcP7EtS8ghRFyc9l5sgRVy4CwfYwQmN5ZikkztoTP0h55t1wlYTdlMCahiR
9GPtvum/Pee3hU4i54Io/7lxDJieq9lGR74+nMeAFdrkhFADo0kNuFZjrFbvAnrXliZFbUSWgfUz
3uTjvxvyFcyfLLDvYBbGM0WMVgzJwhMdYaya7eIk/bM9xMFr1YY/q8MkKmyKe6t+wXUkTJhl9IyK
ZZV3C0ZbO31x8HXZHNmsFs2k0p3Qz0BfWLaOYDDmuvn9ubqwCh5JxkSopk14f9tJAfP9mTyHjrTC
u7SnoSE8UdYsSPjMl4hSRMgJSBJAawie23DSHBVvBjCCJhHCfrwcpg5j8V0p+cxGT6HwwiodkqxD
So5yEpZE1t9GOQEAB2EqqQpMeriRqXj5P0JJoOMSQCC26YoBJ5z10W5/e4TmHCmGumpLWZZXtz3R
Ni043t/cQFftjFZA8UAEkso5oLCagGpQruDTfXLPSAmRHxSx0Zq7Grn64zL8sBABJPktuiDUDK1Q
WTikD+Q9XOGV002uH9CpJjDsoWNrMOJ5oyOpeOxsMqLHzHme8T+3VFzLMeleS6gqXjBdc+QdmSEw
2y3Xr0VpZDH2PpGFqsiLXVgVatwsvrk/7pS0fXurReH8D7XVqstCEEobgtdkrRPcoHVtkKQWaQDQ
8XCfJO3wBb5fXYEsiwXzt660VZAztLowdVhi0e1+lSvJJmg/fyYu54RNG8EXVYn9ZBcr7bhFMD7c
uuY5od6N4mzogQXl6GviI2e28Iq3G9AQVzmiDM2xKS7ubnVRMm8Fp3k3GYQUNsE1051S0gwEx1rO
IuIEvn7urWJYiw/F7PtpQE3jd5iU/Tar0WI1z7sNXlc6WHLm8hzFy8AmVeCpwXRJwGU9CJtq6ek1
vowKfm3u+8VibE+8NVOC9651rcxCwikTVgO/s408+Rj6iu5dyjAuRTebnx0lYIx8tdvssb3xR340
iZkWOPwAF67pe03v46efXTBgqfY2wmHCVWiv/n3HiiCicL4+Wj4acijvUcfZF9LK8KJ+RERO6qsc
O7/QHtjUGfhMq/aBuBJFubhI7X7BExMMYCYC4AL7zoHhc6gEcukt14fbSwZM4aTjl4gsuKrFZprQ
uxqWoPnxvDQqXC6xKQRhDGPyRYAPTC+erGCBHpUW3cBILgUzvOdJM/pgbi8NqH+nQ3RO43IX+fFA
gs1eR4f0qI1XIkVCfjuAlTtewBBOk4zthRGt/UKoFWX+/aRevNOh/1voGxh5rLBm7FcWaGdjUqiS
lVa1spBqM/a/sFFuNVdcGh88POT6XwmD2+75936EfGNRHQGP8INv75a2beCZtEkXmuM1Of6Y0zl4
4kJVWXzi8cM3K/kU5oDvYA36DpUhblzi18utPEZ0mnbaNkH9ttHUTujwe/rlaxYQul5Cq6nj4fAV
ptMGMKKpH+PXr2b1/5HeJDxz1V50P2p0n99FwZeI7RFNgoDpRGRkzch/0Oh+lOikyv13Lqsuoe3H
C8CIK149kEmdPbvMZxqivMrtsfwBjenqSTkzhXJsyJO5u7fW5jRuQTG7JjmumwCyyo/3DgwHvD0q
KVUIn4052P7zw8dIWg/BTrYJQbZKhhK2sUxZd9uNltt/TfloZ0OunrTcw/fCvcZm5JLYFd19uwAf
kUo0tFNO7wEXUcHnszxt1VvuKFu98pkwAd+FTDgxWfXK8SJ9c69q9WroFYnhcITSG6bENkQtGmGq
Ec5kBEwCWbL6Jg+PYuEGfc1obP680+1pARtdxpX15b8/Z/Bu23tb1zDGxpaqxPMPB5V9/gkMFy2W
PRvpC/gDpE55ed5Z97CaHubaJCR1ia8nqGuk1NoDpVCRFhFXw003j0vvCMvSI3EUp8PRb2PvK7Av
WMACo1irIJiikeOKOrpgxRxJuexdmKgCJ0Vcm/tmQqvIqFXAGwq4yVS37lgtkFqmFFwlSBhkKW6T
xHEB0wIco7etD+hT8yszlmf+OL5mDX28FeHLZNbB2QhVYy+mm4YI9S3N2G7EHV/ibE2PegUTYybd
C+gPBacezPVOLNZ5TfHF1HcFRMLTXYyqSnRIQ0XyHvyPktcKnrtbhCyYtF5k4Bw95DnRtUGlwpNJ
wV/cTzUUogwI2VR8uD13Glo97plq+Qkf0e4f4mJpAobmXAW1iWk7UZZe56ClXHhcj5RhmatMaZdw
qX3IBrkS9+qwX0p5Tod/UJ0KKBYjF7R1fpbBlFRXZsFxmTuKgMhnQbumKYYOBzbEueOnkO6DE/Wb
DMIHB1inRHnLagBMXUsC/caoThjq0gE3yLGDQaToFbXDCevT3qGavVOSxVJqK5aspyFCS7Bw3cJY
RuxPbE7MN5pyoKrQwAiMqbHMSIfUMYg7w+dWeuaDnfI+6GFommPvpluy2DHbDgV74r5qrLU9JGxn
bYE3ulhXVF7V/j+mLO/IVRF0Dwyw/MljuVywz2tZuscXpm4H/tm7dEVdOR5OXwKC7UbNO3g3eYUr
LIdSp66IyXyODi/pdqKNamGebljf9MUrsjIW05OtVJW/WTMvjQQxu1uGuNeJnBZvr7gpi4d3YJzL
aWTe0xTynRMVYoXu8Ggc1ljOzu5YHBTBxc7nrZI43LzkipqQsiVOAV5JlISmKL5BVWeDAixGrPnZ
J+uIi0u6RcsVBEWbwGKDiqUkLbYR9XHRERnSGnsbgPyfNrP3cqxsT6fEIG2d07jLPgjjOttZKmP4
m1o1IkbKbVava8Rp5NfhV+KdCLhb0DZVjVArjPCHpHSm4MmABnh0BNoeJr4+bWDNtRiPWeGpsNP0
7PCcxITCVw2OdRAJHWgv52vhO1Gd+9L5WMVObfdczfx5AyNhvnoXPphpHdOJl+LnVECRDTfAGg9r
Ydn6XUh6vZgcBVy7iyJSreBVKhGgGxF3UKgleuiaUEBQwk79mV9HVQvW2OIYytjcO0bVQKrwp8we
QkD6b26zH+53wNxDt6E+Gim/wZ44HOBTd1rzYn+HIDq0mGtD9xK3bUiO3k5l9sWF0cxiU8UWwi8K
zPxJO4idCovpr3ZxeIT9usY8AoUeaRph85Wf+93KnF3ukekxwcZ+7lolLW5IzEaTzxRLLDZ2ilVH
AqT4/UEQqzQdn5hdNBNYzCVW3T9LJ0a96ZKlAYQml0w99dIFOPPXx7Oy3NcBZK7KcGbaurn9CXSV
+rFMHJsVF1UBzCuauLON9ZLOm3Gm5ffZeG0quSlDdKyBGElre+27eH05CVyqjEowkibx/gpKb8oQ
a4OPJI9n3zzHEMc4CH85TEcV1jM8icNrMtV+hX57GXdcCLiJp6eVSfiqSBEz/E9peYlcGgs5cb2H
Iyzm+aUNOi2m/F2bCJKyVZNB6Xgv+BNJNOl21BWUb0sQOLwNwCfOhHQr6/txtJ0AukKWhL/q+5YT
yQ36uBIBaRxCJWCD8ykncTLDA9iyXYXOEO3q+sbNDixk7duHcYxFDK05kWijj2r8jHfqhK5BDg/N
WeztRPyn58VUzmni1crJAww461f4ieMA/36q1zDK2CBl/GuzaiExXG+tOZxlxa4wNvjLppkivt7y
queDO5hsJsyW1CvvPPcz+EfK1HTc6niRT3vGjMqN7yI3df7+vLnsYAztlFM44R5xG8UP3B6OZBdx
b6AtR+TL1izc2DoOP5aShMOQ9eFVBzjhJHnGXsg8NBClRG5WxKO9hGIqHP5nQ8IRilV1qE0yMhPu
qoQf5BdDzDkjZ3tFvLqU4R9puC+g0S1ZwZwbcNyyQ8mpMlUyjzICZAEzkYzyFcXKWD9WTQErqfth
dQNxUuZTnmgcSxZdIMBU7VreJ91yK3icqo7FehnBNZg4gloYyXkn2+OdBs4p1q1coWe8DHa1Y7dr
lsKqpcHWiDe5/n89F3+GbSbKNRlI7R9Ngp+DOBS5UzdGFbN6giD4puoxGVQJYJ/gK9jyIJ0KO9ZE
yil4PDZR1ue55CwM1L64+Zpss0izBtP24R44q3DR3AHepAc3Zw4KhiggaP67SJ2DdHe0W9x3C8st
s7C1GMu6avdX8P947LVZqItlZyqfEud2R3lXPkuMnHk8b6zzRPjZ47eqYPCuQzj6LfPfRClCwua3
oH7rRtRnquJs3JdYKoT7pX0U2toJy5Q50UyTIvbA3cNFv3l8Nb2x1qXJ37j1lQBDZLGL5Ujb//ii
Vf43dlKPBkXCfNthf2jP1tCGQlBqebH9fRFfnqF6U+XwLnlTaEyZ9M1QMnJt30VCpvcekKEEzGez
7nWdY3zDTh8SpLoCXP3MIzHH2JCDW1dzjH6kRF66wzxvILblcN7PZ5scth25V+QW8QwFlQHselA8
gTUpjp5NHTRPFd4d6YbomfY/YIoYWryPABsNZKOF7GAPOaysCsW91rWXeaP3ILWiSq4jmUCa2Bnx
aEcf9NBxQIK3Kr/Di7Hl/0WQaflHA9s506ZjpRvT4do9jty/O2v7POvljdXoJ+3xiyc4+014THos
T8F5/qAwMyKMEFOsBi8i7k/xdoONdqctDsBMfZSkjH+ocFVp/xbnwX3Rk9q2BrWbEV30frgM47wR
PbsJoTlvSqCUwX0Q9wjnGbjJ3HbBYgi9UahCR2BgEsZua25zCUEB8nogQW5Szm6fg38PoZCIHptJ
tj34OFUDFC+qs4K8TVDms0Tu7oHTsm4+IQ57mnXrqkr+PCuWd+WaskbYwAhytgg+wAhe+l6JMfNi
Vh2KmHilanwDw/3CpIHimFPOCXzOQvFfnEFJhA369QoDBNeTMYaPV55NpeRgLIshnyO2jXpoZgls
2vsR9rCoT4mfRFH9SSnjobTIqU4ksKH/CNYOU46lePZdf/sxH52pd/Cnhluw5irEBe58a3N5IwoM
CcKzm8sjYRTsytXk6JUahomLHNkSHlb5gY5Sf5Iikd7uVTKzFD3WSc3cWdN2/4ZPIJ/hyllLiIBI
N63X8P8bPeUWyOZLpH72cz8f7BiorWiO1a4ElZVxYDnJAY2wKjqevpoFViTNRslejdVEhxKCn5w1
VCgLRDOWS1xjF+BqbhFPhvYeHGG1Z08K8dA1ISOp7Tsfo+cDfFWHXkr6xhTQHNXJe5wJsoGkczfv
6mku5HWTjXIi8CvPMcGHfO2BUdjIs7BYqdQTnEueWn1wAmG5vJ8IxGFoV7R5S95Zzwx1vQX39lpD
Olh1N0TvWUVHIeTOzCw9/xJoGWdTy5Ut7LD/di4cfzfSxjZGb08O2psKG3pFzm+VzBoMHApilN5j
E8nmFpW0lwEANH2xgr5UwtRSwP6RPEc6jl/XKmaRlWG3AshJcjEmHjBQWiK1AWxyOYZro2eet70q
bdyuAcJVQkRb1NYRxN6iboxQsL4dSEHz6MlXJBzaN4G2nAtOhWid7N4nFAwqV5R1aJF1Bg8fz3+T
TWdwKVqdU+Nb3gxmQAIEOSjgBuKfLRuyYO9btSkS4mSjsuXde7TFau+gOY7ZOuMxbO4tmw+U523H
2/aBuD3KQ5x2nWhHxgZYJQIht8zw5RiPsa/tS7ssyzbGUmp1IePR0gzgVqNmEd9QI6X7p7RUOoUt
9GYQVqbq8TdKWHAL9UXLAz3cU6MK6ue82c/YPdwKsn7nTwOu/xmTGWw2Hqi3ZxuFImck/QUMp8Sl
/kLtULfeUYev8z7AxaTnrYlYa9OZSpuWPTY8YDtTNpSu9z3fqwNfMO/DkKcJIgGOFYj+4TF913Qe
mtJBNLwQmud+GZWgj+SkR4CrH/PCP02aOrz9jz7Uap19J74s9M8buhOuMVhQC7Cxhm8MENoqTqy5
BHl5lw/jMwhK5BwOqv4LOAz7K61XUfIaePT7sTmBKknl8cZLvrokcFGUEpVpV3ORzOrY/AMcDghv
bto2UEJbaZ9uLsNyHci8NdRX6XKn2Wd4qmz/DpUDoqLX9bnPRs7o1+ksfG9+TH1iSYwlja2PPZZI
qvUqXHZQO8sYeLlhVpkYhLideJUfZnGvrWfIMJ6eHNysxZU606GPctOVfxrRGcs0Yz72nqTbats3
t/aGUAfqtilK5mgtiQx5C5B9T1FDhRgmU/rcbZnr1obXXASYDvvcL/AqPw3gefd1R8sJuN/MKtGV
2GAK3LFd9G7HRk0jrR4oNP74Eo2KiBxdGVon62qfuSt/r8i9EjMA2jvmRY1gudJXEwywk+F19/xJ
noHP64n+FjKp2vNu/0y4JMQRwq5dSnr9Wx/don9lUFhyJx14vfoHkLMTEipCAPR+68zRiWrZ+mRh
dR5uiEPibQK9BxgY0Dah8byzxXad+cByrhEGQ7aiBtm3VkqOACqZPRx6b1Pjzr/H4QGC/NYOaU/S
PQy75mYXkkM+MJZvb72rNN37QmGwL6hLEwymGhyfb7jCb2w7uwtUU1vKBJv1OUmxmhEc8/6gwxga
co3aYIhL1cg5FnQRfl8UfFOf8YqF0I3HD1DgGdSCLJcgyW4tP1e3cebtGCUGH2dhuJlo41oephJ9
hZXtzA1BgL/kf6zdQ0AQbFVITgehcSGfWEcl1Mcdm6BJT3pvMtz5i85W8kVh6bQud58PP67J747G
gx5h04KrP7vLf4uS3hF6mNsbYsZSMQ9KYdB6czbU1pY/piLmbwz9q0LJPu6eY/oCYpaf95PyvD6f
kija2A5EA+6W9U3IyoBL1CIl8nh8zrkuQgUXjUD2M5I9X+eCQ/lONbe1kxXAavPJalgBWNswuTpR
O8/glaUUoXRDXDRiModjE+j6deqVFBlTFq+qWxnEowatMszaWUmKfenf0BSqBllCtyHLGwnBUBeV
rmpLcQs6sY2G+xhF7mQgwCdbGiS94qT3HT4Wm35FzKdcJxT1WiydvgMPyzLqvpqidpnjiPaTRJ0n
jCFzhCTJSlFdTpnxOskbNb0Z95ctxi1cDMkHnBaAMbEA4d3OtpmvChG+h47CvjAFNbF7sg7vq73k
7iUOqj1VCNY+5DOOnndNWSNXXMuGT+mCOLD0Kj8sJj0xiI0OT/c6i690K+NNuwWSZxxb6Sey0T78
Tb39gdG0Pwf/yIQT9XxKLH+jpsNhMTpN5PDbtaIAwvDRoceH/JcmmFZ99ctjbkF+Yz3QqzJznSMv
mrdyUdGYrlTTXSXJw/DlIWeAG47rVvFZUM6Nsr6HPccROhWAH0ZQNQzvXv1WLecvMHfCZ8TlWGeJ
IEGMPpfXIABRBuHYdnsBC/azvWBcdXsjXYh4QMeJO7wzGsv97QS+ZxhYXykYjK8jtvmvoVIMVHzv
VHmnG3NUwg0Az1O6Id4A1MZnG3fm0zTHE+kvBgCLfUiHtiJEDAd/kDpg5SI9feGxzDTimxAP/FMZ
I47493Fi7fVc90B30pVk/Y7O33ue7ecWoGPVL7Rys0skNv0wolVblndDIHVV+Uwv+wlHGeuwIc4c
GmD5wbPghduZV2nXGI+vlLKx4B9Zk54bkndpHZlh29tbQpl4LLmbXglZaI6nXfq4swUmj3/Qxzau
Rt9DZttePiDrqAc+ZhYdmfT0k+ib8POlIcI0C6zOlb6VA44MlyFac8YqfXdb4+jNd/PphU/X81LO
pQ6uxyNCcv7J6Jv21ONwXuMFiC4QKvfz3+kdyo9Tns0txPwQFEzGTKn+oW4a0RcTqKJHlIGFabp1
u9CyNj9rq/+0xpfpkvmQvzUN4MTr7tQe4xUrh94KnFSMuXMwXWozt8db7gFs7QtywG/+1LV2kJ2o
XCSSd+oQI+JLzJrxDOph022RPI9YrJqm2LrtFA9RWYU9sAQn7M55WPA+r/Z087ypbrT1B8h6kWkI
y5NOq528ugGJAT07XsaT4khuMVdFq7Iu1KJsKAVKITDnyexyNt46BPzY3ibjlOWWVq+rTJMDg2TE
VWwpEqkiPuajteWlcRIViUr+4QnaIEUx8fY76Lpph9mbp2qUBfjI7bIwsXsG2bcYMt1IoQKDakl2
3GaUWrJuBDDGVXmW064BLwG35ooxVN/JMD/EP+8vWHvVL0sj7aVvj0P7eYnzsjIweP+eNfi1REoX
LSI8HevGHZnUswzSYnTR1rXU2TqjuUKGuEl+wmwq6HdaLfAAI13ssLXAgd1Dqnpahp7atPUS7QH3
OtygpCwDPXx1v3Sq01KeESGA8FD5d4++Hj2SIQSP3lORjsuuWXDCbGlS0lxg5rnxz5P8heZ209M0
zJCheYcKuEc4ko823jIri5DhkVvwbJYmHq2vaeEWG1BQsO9zLLbj3Dvu2QDq6i69zCTtOV+BG4YQ
kYwUvlffgWDpqeBIoneBDq9q4HPkAPsnUWcz1lBJyaqnV9/M1xPYHpQQMUub8s2wtVQrDKbT9yqO
b/dnDOnlBgI/ogacuJQRGi5U6hg3JRNnfMZtmpl5es0aceuwpLUq1wrSMOK4Mq9jJ/RWvpMfA7I0
y5RMeZgzKx2SxFquuIyW0g7zGIRH8J86vuHX6pcT2yIMkcrZ8R1mK6MP3Q/JZ0oBRFOJ+yXQS43c
rEx5ChOJwGAQ241gdGV1hoLQjRd+vaK+j0y4XlqQdRYz5A7aj3bvqRJI/xKkgWVrYQzttEfxS6SV
jJq+L5h/LPak6AcaRETQcRiOX3OgJP0P6+w7MLJ603OZ/M/IF+ACKMoqo14ofBb+FXjyrMrqGsPH
/p9XUEtZgqme7XWV9b3/GlKyCBdvqg35MhAUhzcqJbKQGKjmHa8hpiGZqkEUmsuMrcStNICz9VXt
PugTT5Tn0d7AN+2fo5XC707dIh6ZPocLgrFO328J++QIKj2QjHj3sEi/B7qEIUzIx44M3aGiNn3s
hlBdXpvfaSvRlmAlqOj8/waHPv4QD2pO9j+87JlYZpwIKR20I9pf/a5zYZhxnTC1bdnWtyYgHLjj
SeDHO0JKmeOvkio7q68qqd4kLdCXAb0vp8Yyt2BaQksi3ed81MkuRWRYAkMba6/5Sm77jAzTwiz7
41svLvl1kb/ceHL4vUwKSTmoIrfnJwJy4s7pnBV0dhZMsrwoKFAzOs96IOghUUaMModFc7Abdnvm
IOrjFOnC18nTEuq8XrNuikGbmzo415TiMWBAjYNkyq6PyIUiiwEuHeq7WHP1nlUv30mS6LzAqROX
ibv6EW0SozPD1/LtM1DfoYrnMKSaE0CgeVBMrkLAE4SKrX+7ux263P/kvm28k6vnKMPsAl69x8zZ
5m2i6UIUuuBIa+cdum8pNr3KaBYRAgGIRgal1u2e4sZZw+USJPwutAJJu7DdXK8nmSc9JdTozmpp
sRYan4F1y/SUU//qOvuTPKcvP2SgWAOTxqMu6LJ/51GiZrTO9QzcbSdfzfxuaYvp3AfyXrdodK1y
Dh7GxC1LX7mAeYKb3p9jenvRDdiGK8AMdchDLgXhjfUozeMHv0ZL6dHEZD8ITT68oOmNiKkd0MUa
CNDHLXTQ72S560JSEJyBdgwOLAUnGbWwzJ4p8ePf1WUU3cO8GCBCiTOnGtdz7VhmF35Xsy4OfjO0
ryV0X3usZI5SafOYUdmsqOnpJrUpFow05kdzPlprxh3lgZEciRXAAVh/dkpPw/DhtuKruzmwOeQ/
zXcl5ocexm/1aErBLcigd3SsBUtDexATG1VUZv/Bu15t7d/e5InGynD/qqJiUtSV8LMh2oNaCnbm
Ok38NkknGiIRC7Lyr3lb5G7YeCxBcLaCQWvBpOq3dypjzw7rydbuPt/DKXZG751f6EmwKjYzMO9v
+JIj/x7QSacxFSoVeGoNZsyrHx8nTVKe16GD6sVoUfw7VLgu68W+IwTHL4m8Q7qYYUeCFmFj0Pyd
a5yu5rXlP52M9fu1j03Zx8ZVWjO1/57wDkOcljvA5en/hAV7vY020sDzKg9rL7Nh1ITrEjRBLNyX
Hniw+1zVHlEgMYr5b1CCpEHeS3l5Y9ZyW0kpzmlOQiIeZVQnz6EpgbsLG3+yWXv2tF0zlunRbov9
ggdxsax4lVD3dGtfUFbEY0EoQGIT/4VDWr1VgCOJvostw5pz9SfWt2B2bw0CZaX4R3LiPcvY1dvZ
mO5R/fAF0IlOy5o9jX8C9dG4PmHHKiSeXoWoE7AQUA8amjVUYd5WrdhrOAhwq8/FiiAlluEqWBZ7
+gVhsT0eUn+egsHJK7T0mU7L29dlBcx8o9coY6RD26jF6HcxKYQEFsV7Cg9IzyR58E8d6m+aQAVV
2ZglPtr+LBg9oDtAQkbLKl7DnQt2sm+TGSDUrjE8bl3Cxf6pn8P7om9Sp7Eldykj4HlM6eXbLAtY
Z8WiOQOIHcxGTecEuPNPnKzapNsgOPlqvTwnaAF0YLUVCLwLqAJ30wweW0gFra57OecHIuEOAH6s
LaCJDXFHJ2lPDLRG61benYuWN4qnc/Q9BmFSQvZIwfragq6dcp0Y8V5pksVG0yvmBTCqs7jvvj8x
s3jUw8EzLoS1PyLCptSMWU1/aHWLQF6uQ2FXY/YboiuWMtbbALr1KEByvXzOsMi5OpDKEYWegBH1
pxedNDK/NYKOYrzsKRoo8O1TGaN1xYp4DdwREFm7i8A4b/5S3ogyXzKD0je+gPSHLhEn4mn2x0Tx
6dfHBIbA9mxkcaU8OZ3LUoYpKAinwIjMgF7x36884vjrZtm2uqk502Mhu8GSFNtwaKp9lJ+lpc0n
NmOFsgtir6fPQVKgDp+YAI1qNR4mW59fedDmX25fY3YwrO2XIFMHk7WLjiZkJBk2LZJGYEeNZ5nP
i2LQ2gHNPiSBmunb/l6kF0nC0hPSOTv9OrMtBYONWKjWt83knYHKa9FqK+4x6Nzjp7/sIOz/IVTN
XnUfWyPiNpH5Np/UiVYnsxxdplIj5/eO4Vsz2/kU3mDY96skX8pF+G0FX1zcT5bmqRfjU/SW0+U7
HvWUQPzVt2kXqJaQxHrkFd27x1fnavKEGpqbVpzLC+kNmEwd3riMYAT+cn3TWrQCcnGDrdaLrpm9
Uy+QTGPSSMttSO7ePFc1lQylqzjNyaUunEJ8Ya2uWC84zfxpL7EM8M1h/u1kf0I+oV5WNJ5JKaKO
Ve2DBY3rk1B0uEHa+h426/swRBAHE6o6YQtGvhyuduqLEjenZy2Xq1D8SCDHapk7JsQ90JPfVfzx
eX6taHbz6tZ4mIIN1SI2vGGqAZaVGGJP+V5SOegf8cQRgS0bN70gUAwqcTfJnHf8rkMlH5lM0kgx
C9pq/NMNjYQTXVywiCI9uYI+pkKC4HYRcR1owGHuw4nUBT2aZbNgXqq4aLd7tPGZ71PZmNoDt1OX
oSl+Imrw99AdsoYi/+PMfjpQF18hxL+I+RXIZwy2BifAdXaZZS0s2nnvPa4+UeDBawPGNvWldQlw
pFhzOxV3dTg9fvareMaCFf2z0QUNbyVokwBS+D+EjCgAfWpjBG50hdkBLmjcIPYJfPUwO3DIyTFI
aqkBTg7TyH2idp4mABbEzSTyMGk34ja8quzTnHwJEe/3P0xB+9SIRpKE2Vw3H/DFtMpKRpXQQ3gF
CZ5PCRzBZ1bacPF0Bv0937BNH2/ZFKArHfwhoBhF/ghsNSF6TUqidOZpzeqfoggrYh5bV8mxauVr
4+ZXmK36zgoTAOdfkTXxNSPf9RZ9c6zCcEs3CMTo1TTRdbXgtKSkMzIB9qpGkPiW7o/ydi/b7igT
ycXcp6+A5/puz62MBzaTpOfuf2Ba4ADBL67JRFL6O5Rrpug2qAnIhDREyxKyz7T9Z3vGlSeONGVE
mvlXg8FPaIz9jLItE8oKTepOVLT96KwlNJhcdh7kBRwW5aWm+I0/A/w5Dt0cYI/X9ROJk+wQ5asG
IK5DDUbvn4E5O1lHSLn6H4TUCl4xtcfi/vLv6cY8+TOwp8DYMHkzMlC6C2n6m8JHfq8Iw2sYi2So
D5Ibz46p+2tlsZWH1xy9RrXfTF64ySFBxFQBp+LMNZtVjVs/h+8gBX8ncnteVrTPa4wfSpMi3o6t
xfCcDt1o5xMM4dfDXu0kFUeKRp7SEPcpGwUwwgHaN8C4DIoQ6oE/mtc7RlHGvOr/l6x272WAR1RX
C/aCCB9wb6ZSgIRzyd5UsLuzHY0L3EdUyTMzvNhl4nEHiBBUqHEtOWKM5Tkn9gJvaFTUGzrARhMS
3Zy/aUVpU3uEA6NKBA035t/iL2K+OO6k+TsUDxKCjDEWt3zq17ONdu3COkd/HUshfUNv+k8jQDsi
fsrE+yMDwCs36BbZuWvC5ixnwODZBWEa4dJVCAALAJcv4mIRZoTRoxyYdZtjtv7ipQ5y08xR0CNU
u5igRYUUeuDIZsgvS6dD6xJYKFsAxR/BmXaqZGU/RQ1C6AneIWeDIGtAh+BuSlhfl/fVjaEFnNaV
YxwBvakFQUkosBMX6ydtthloKQUmDgW54qSYBASUJ81n0hENbySYfinE6HJXeJYWKoZMlgbvRlAF
5cLohzaefE4ZGTqet/VKelwlKK5N1TGcjsH/zkBdj5xbeXjQAFWAJV6+OCqfEzpk1X1X/ZQP3LtZ
S6M36XVRMkw3qaZyOvLGUwH9s+X6w3YccG0c+0LBsW0+9DuADbE7WncCirgD7VDc4wxn4V0ih5Hp
YWew/B3p4RxMjqMoG/27mzCapOWuDeR7jKgBf0djaWNPnO5bPuiDeve6Cf+Zs6adCD0Ob0Oggx4r
wHVXEvCYUU6FUVAVr2mTn62J1J2S4BwSc7jZ/dKa3WMY5LcHJuv7Wau55rrHNF8toNxkDMuV2qaF
ZgV4rzjgerHabUP3k0jWyaD+VJZTOGHpxEJG57V9V0w2JmLDKXIINDvhT+dnELY6GeiuoQXVg8tK
Gic9hyakW2ZSo7bcW73nQzYGPJjQZOwYivM6otIa33ym07uZdI95WSzHQn9My6ZbfMSeBRZyXNga
XOtB/Oi3uOF4vhOBhLoP9u+LOhfoN3HQEwxlhB2qvnP6A9ttenOzldaZXuoxQ0C5jaGY/gH1a5/y
FwXXGzKZLu4+Dbxv5yDG1EtLPREtb15UQos9nSuXxg4NZLa89dwaW8Tadn+yntc0iAqLNzzatv+9
lpIIK/JD19NQ3y8GMVTk9a3b9l5AtHQN6QiMAD7pzxN3C3lY8D8RoSsbuWjC1yeIDHpDjXGD+zCI
hqQVOFHIJ3Ig9JWMEE7j7l9ms8bvse7UCn6Wh1jCaRHkdikWyM3uSQOjJba0N6n4ine3S5/yGLOC
/mwxecPMTmzGypzr1ZqFdl90yn3NKSXyTQd0KYBpuvSQ4ajsAIyoZsCVKK068YQQ2sx0YInVwAT/
Sg4u7vxETCOPBFx6fJExSgnExoUOKVyJhox5/9+VrKGXxWRtuKAuuSkkgIBiwqZjOSoE4DDDwbF0
YCpxrWoDrrGtCMYHUAsYseKjq+SN/I69cqrHNRd+ZM1gmUoPzglX9dm4OFRkB/dDvDbMF4MfTjWK
LQVwnYeEqv6CRn+V4p5fv0c8PgnAUMoWZXFNkY4/DR3cF+lQ1uFOIwpwt6kuz/IPrroTYYNxV+QY
WiL0qws9BeneKSVPHG9aKsTedPc3hBhcDO2LiK37+S7eCAVJvshUog1SLX9gHIAhiGOOprVf7Ey4
EN9BBvC5zdp5IE8B9eaMx+aHXWSd7c+xwN3l8/IUnhNKkjgoy1Gz19GeNZEtPppy9wGZtMOY2V9t
lb6UXCdwZ9WtRbJa+HxxjPBoX/h198G2C34/4jLZFFACpoPVu59JxNdXM1kTzUJGJzpuhLgo3Pq9
su4HTfM9x8h/AkTQ1wYnxwX47xRlMShbw1ne/yIsL0N5QtBDHRn3mGNITfKO7m/SYpoJdNubDGNQ
dYUOGYCKDblOePVXDFqgEEvhso7OdXm2EYuOx9Tj1DlusqxE962MVu3d8evQjwUaOy9tPFoL6Ebx
JIfjcPgUD9ODB7XNwk8IhSzOpf4AM344NFvCzR771Y9iED1yfaGAQXlR/zvJSdEQixVzJGnh5AR5
OyK6ZfPkF79HvHWuTqrfuA7SkBLNNWHNNbYVkxIBggiV0Qktr0gZENdu3gAibpPxLDPDZhGbfjeG
fsm2W1MgBserYkTxOJqpS/qd9aCrTsIoV6nUEjmZRO6bD77sOdtY8g5hKPw71pFJhadPER09sMWW
N5T+c5zyG5qz9MO/1vYWzj/J4KGye9RWheLamWZjSpipCxitdVU1GqusiN7wBgZdlh8FNPerw1vx
56aHKe2B1hPBHNkLH2J43ETWSak1e41zzil6fNcCVWT4reQss08t1vafsyuoezXNtbJ+cyrGbtbu
dHLI/Bp1XfQtT85jsTkhPnrMxVgSG3EsRlgf78zHZTAjBfaTkvUVSlEMphad+1HZsvll4W3tttOD
JFqa+JGqRcv7wF7VaZouK5KwfLVTygN7pxptFdHHQC/4Igbirex8mSb1yucLCaxyhfmBx5tXk2Hr
zmDWzjs/YcPhNzYNTkhT9JSm8jp5t3ipppPYZdf8OLUpdBcDxN92I/NYY6qIEDvlfBvyCZ16ap/i
eiK/0aVbReVQbX0WD+JOb29NQfyxcZtuEWC8NO9phbkETnTV8JLj5yAGGwaGqIcGLxmZgLw6LckK
nP8AsviNzcvJAU8HYz+v84w4qCXFYeTc/+/pRhXOHhZG9kSBJtkg6mq4gZeHd7nCu6+E2J8vEoPE
vPszlc/6Zq2NQzXyUm5zJQL/YJPU0esrtj9tTnAWHcmSJ8lPaj46P6awZBvICD917GXJPcJbe9ZX
wBQij5cjVmgjULNf5lu23xZizqlgs7Ele31k2Jvj2uQ21+pl9bzljfPOXt/bT5NOyjHNf2Tnw3yr
y9ggRbXpRcmiaUcE8ILr2GhdxF8YNDuuUM/60c1E5fuLdBoIaZuCMuzrx0JzMbJDQ1bzJaCMowbX
hm8+2L7jDW+uZaBzQGJzTd0cHXKNcSWmWZxWJwKClr5+pju+fXGkqex7wyumhzbrlOpigs+wbL26
EUF8ZtiCJ5zU/sVUPYtOeBdpJ1/KXAo/cwAck+SwzrL4VX6uc24AxsvtvroXDRSTDaLs155QlXrV
/Pb2P3+71OrmqwSrLvEgLggBsrBlKMo5kTt4m6mUUrdTJdclB+y6aZuEtlmhgSuwSS9/CcGjZDZR
roc62nLvEHd0+zqhFFqgEZ6bl2iU3mJ8DMtvPF5ojZ9tp/wejy+rG8N0V04Qg3/tbP6v2oYgmYUd
YAwln874t3gMQotIU567lKCEZZEN+vtJdIUwaGHL31DKeSbBlP7XYVcwlEaJ9n1s5jpcBWUtcD7U
3AoXbNHiacfEgAMRyWFqVhKZRJOTkzOUEr8htEB2ag1HUBft5bzBQePWBOMWc+HyJocK6SZ8toiE
nt1tFkxMq3cfldR92PB2gsjqsiVBsjcX871mm13DZrbfDhbCgLmQQ/w2fj9l1i67znmjkz09LYkb
I7OFIaHY4ClE9aX8gZVvVvcxz4laHGGxEcc3dggN1flFek5TyI951yTAzY/GXDcd1zfH5nq3p3w0
RkWMuyFmzZbBIo/rn4UKilwLUJElqrkYlHwZ4gxz+HXUm1CRn+QbUo4qQm5m8W6gsAN69hei7/W0
djSlLtnmAmTCcG2qTNVZevB2cwHRV0obQuaIVzlTRxtiZ572GIaG5otYf0h0rLbNgDjjTRtxJRuE
sg2UZgy1S0Sc924vZQgk5AiwOJLmkPXntHN4gchezf53hlfAAmCMKWqbGYUU03UXwL7phToEewdL
Ylv6Ll4xr/1ihfH8g2xeR6iwbuUQ6kzuoxtR9lqulAwh7P2+CDL6olkuR4ty4L9IaPT9AT0sikcZ
W73n6MLjnkLNsd5AKNBvLc/ZRpHFxqYbmipJN0Esyuwh39luNepyeURMG8ke8z7s4jErIoSp/wza
wacdPC/wLIHtkNMmTtR/u2PElWz9wUDQLshShgW6zMvAEpLty/rXPjNDyoP5AK/NsONlqyhrgShW
8dyl0iE+ZHe4IPMzwekwR/ENBnuAmPVF+Dyh+LqOcXX/XKGOFNYp04BzIbKuj4CYzKQu3uYRmisR
FvfvQ49fgddHhIXKRp37xNkYzqbuj2wINSI47xzppsP67VsRU4EB4Uk/CVSxBrSvd3Y/hYF1P+BY
+yKI23NdWd2qD1IywX69aCxLLCNObacFURYr5pPUAYeREFlHfXVKmk0HeAl43Ug/OTy/23d13GHj
dxB4ubZYhw0QAHF3ys2VCE3D9HGn9zXWA9U5y4p7isYSmXgeUZndkhIcvsIdCGJlArFT4HPGcswK
Ed6TSXpmlWnmO0cU+o8K9vKMxE3k046gtazrm8Se/t19ZjJCPcA7y//7ofWqS/uwg65qqAvTszK9
MR4whsOCejZTRIGMlMD1/Iz+JQEHhbHkPi+IDUkckKqkoN3cXPkRD7DH/S25VA6h2k2CohoECuOt
FcU5WrS/Ak1HduZIIhsiuLfy0dS+dsZ6MWnOnapE/9KjVcjjUowGfvRBwSNIX8niKfY5Kdhz29k+
YLiNWb+YftMfsKAOEigJCNxOFA33VRE19jcTT1AdhLmQoYxjRPP2v2OJIyhZqY3ek9a5T5/Einj/
h1K7MniJ93fEz48B8LyBI3HWGsDMdy6vk1V/F0IXIJ/uDANJia/3nL/sUYaO8c5iHARbxXcbXqeO
JS2psnpDbz3wVNMZjCZQVXRNbL89KYpKGQ/iVlHg36EM+Ox2Ow0S2Q2xVNNQsDI4LtI68jg9YA1Y
u89ePliRLVmO5jgHw9Bjhs/BLyJBESwfZ4RP5tMU5YIqD4fHi/YIeTqo5DXt5NZj5KH1Afr/0f0y
7Om9nL9L1Xb9oGhSISU8FGkoHwO8rJ+fW677KqEMSnX2tmifTWh385fj+t6T3wx9PsORgkGu8Fwg
2LRQk9RMKYXRk7Z095tx9nPU5QZGenDjoxrmxTP6TH63lecHTnIaGHdKR26Wmn+kUD8oO84vWJ2M
Tg1tBxIh4JL4ngQYN0MdqGsR6HfryMUcs4rQsxSPZhowIlYcHyN86//Ex7xglfCAOGVZb1utXMd4
GORdsAPeFEymSdv0kZ7el9gA2qPW6KL/tTuvRUbSfPjYGzwjMDzyGp7oPq1699gquVahpv9hLNSl
Mgw6i85waefiIh0u0hVY1XhG1PMikXVb/LOV4CLR0cOf0t0EnuMWbSV42UM//FxLd0Map3duJPS8
8B8Xbw62kG3gsYqK3ziVXru/z9OB9Fy2GHQG4d0QaW0z507CLJHwrVQoXZSBGHVW1CKryt6vYaKK
PxuJr4jUgU3kFsX0s7Env5DuCG8xvj3Yit9992cz673njPIKlRt4zO33kohtw9ZaXQrhexpGLwyN
q3OAce2KeqO99Ct4Hvvu2LBAM+nabhujtuw1wI42/5qyupStSwJKYiaTlbBO0F03j960pdijCskW
mFENsCsPLAHDCj/XwpohYpzcwPF2iqwaJ0xx7yGdqMx84oIItQlVkqsJ62CcvCKltPQnEuxJCxcR
cSmC26Pm9OwnDMJaAi2XPYhn1P2MJYfLMVEELSdiF830LGB0ENH3theE8jjAS/UcDVRySILDkxEx
DxtEFL9/IU6cG3ywKdhvrHZSdTiKC2y7jwXQGHryCaT+hwOLzsT8cP/cyMRlR/Q4bbsve4zSzQHz
64yV0LTkExqlSOOW1nTIad7Wxj4DM2MsmiF1RVOyERuTSYbTsUmAbr6nsVss1ipo+6R6DW04GyJK
IMBv0bLMAwl/nbhh3+8WBUHpcwcPzdWGr6umPWGBeEQXPnYoeE51Ybrpwi1gKl1OX/NKf6RVNy2X
6LzaDk6V7zte0tjDDI2kY7I4lyE9o1534pSR+DHksszdCaYfxH78mrRe4xBDoQMxHSwK/GTeCiRU
UbP1SLCk2Ut+g6McowWZJGWxlW2X+zH71IJYCI5Uhuch2VYvG9dJczqoqcfM40nOHEx+Wm+s0PbU
YHUfL5gtQelQ7ssagrJSOD/DYHxE3+Ux+3Z8lJkEEfaoMSfmxVFX0Awgs0XAxVSJKb9BQ8rMKpyp
XJ4sOQaVTD3reoB1cuXE8OnldT7ypVl9Lyc8hYlHtsmHG6Z9zIm4+OLzlGNEQ9eBBd3+J+bTmLTW
OPhO80l/szUqwuYV2SlZ+YtCxfzl21v1wv1/2pOlF7cPj6ejn42w08mqxt9P0JwU8qFwW8z9ylJ+
FhxonMDP6aKkxfJPpQk/cGqC9Bof6h5P9bqDHTiWsLs8ZXsl3r2KVVIIs0Ep6TOdyb0rHKzmM958
g/yJiuY0R8T5+TpQ16upUGXLBQo6vIbq0g+TgdmTQcKV9clpkMjTfHI3NYomhZr7pYumZkrOCeV8
y1oVpMOEjPcVSGMCAc272qsNTwGgDquA2ShbGjo0mnCO2F5wBIHfCwSP+v9V9REKdU9wIBYJYORX
Te2tWTxJ0Eu32Abie0dsb5yd0393BM18TBIQ0RHvM5RHTPTkOND+XWL2V4WUjUKgU/IIhUFc0+ZG
5SXoFTSsFwL4FNPiUlOG2yWymY0EwPwrE7MmpFYPvlQ9/x2FMvNoThssoGWRl3qT/YEaTcRPB0eo
V43ShrBatuCDyjqeaVHkpmolXeMoMQZRqcanFIKKxh7DcW63IkDEsI1XM8Bro0GfOqbtAH935d1t
qGilA2ONFhsZreguKdwKqpL/4P9ge22YPpn2tGLzNh7wKCn7WjEJBdjYtgOC15c9GUMVYXD19FXP
68ZOjWGATgdVe6je4fmZlUHmES9rme10G7jZjvSnxKbja9rdRYEz1eeig0XA6GNS7AjH59JoGyt1
K+FJd0ANxpnrs+bAkNEuCfJhJmcZHT5tKcIHWzNx5ZrNe8pjifvR4+qR/z8UvQVN8HKmVFx7Tjfz
REywm5oCANogj12+qT3hyRd9sggTwNvQ6B+s9P1WiTHFPns5HuumqanXAmtkT/ylG76zzNlKkNP+
+XjS+C6C0MfnzJCXIioNloh18OB/T6hWs5qbLxT9RJAfoyF10MF3GJ0K3BOXLAiFWX8M3+bQLzsk
dPAtvOEMujfiQbaRCmDjrtBYgzuJsHZUN98h93HcJgdgGwDcKBzJKeG2mp/56RLp2kSid82ihHaL
hLJ+X9/rdACoJ79/LLarN4RtT0XwiQCVs8iZIqIcFGtJiXk/VAtOGRg/aY8BExYzxxZw/fSSQFYk
Fnnug3SFOOsswaR/lwFTGID3VneP2hrfU+FQB4H0cNmge7Zxf5amZL3dDre1coHI9sdA3eIaYqjV
nyRM9zQNlph4szQebEjv2SLBpeLYV74Pn0JNQdjyHn9V2QYr+aRazPwb4if4AcjM4B5M0O1hzaj+
DPW9/uEpowTaZchYP6gf6VMjyy95unKpNucVt2BdF6Jgr3PhW38DjcbOhTWkOHWrW41Q9koGMLDj
s77Mi0u3cLFiMvu2CPEUk+z19T79ZpeFNyeEbmy/spvhREylHa8VtEqD+8IN01hXjWsrSAmz+iQQ
jV3+xhuhkpBUL/CfxCvVLnfKghjAxthbTkS7W/8uPmUi7YtOVQRz6XSa7T6GKPIi1biND0OTmL03
GzNUdquyOPvxdsKXWeL7yaerkGVoZy3cP6i57GVvDPXLaFWTt8OitAXgN2h8tXmRxHogeKPopPwU
EvN7hyi4Kvlwywkbqcvf9Oeav4o6+OkP5Y3lO93a61rYz/dRSvY1GWZWeQJ53kE7r7bIHxvCHgHM
voLpkBT84OMAqUhjWf9tNLKyxX0w/cUFSpzSZhLeT08oWTv8/VZwnhCXXvwtxbWmHmsCU6L8sBor
Fa143Zqmp+LkGfMopSQzMK7wWZmoCoM/hlewTAwVdCE24mCL7XW6Gw/UlCJk5kNghrvuZ5OLJS2H
VFbgcBi222W+fQluS5Tp/7fJH7Abm7dqbzMUlNlzFQr1Sy4kuXsCwyXex2S+d5ZCaQ5VfWvQ03Rl
LKwKLc/GNq0A5xwUxu9QR2WrrTf17jTCUwsk4tbl5hWtXRcHqzAHMb5f3KPmhQH+7c7U6YyUcvr5
7Ybmnjkp7aU5LcKX+DXT+222dl+0hGHVfy1M+PMh93Wrk5P9Uekd5eoFGqAUZOSg7KlF7xgVyK4Q
qXSPNY8jm40EbaNFJSyJt5O3EGQ6JgFeQS63ANcFN3sGv0V/YT5uJupKhqtLs+5hyQWRQjfO3SAA
WmZAdWLnMIc4LZ62aW3U1qGaQJvwuBDTO8vk0C6JdHsiZHwnpAHTeHblxmVD41R8hJrER0auOrIt
o548e970zhIFco/vb6lrtmCzntEwhI0XHoHkb67FnKBILG+NjXGm3s0vbfRt3ulYphUVAsO0EZUZ
evoE50SSCdaMC3UXWX84zW4lCBcXFkBhViM1GovNTKUHxO6v0Fvj9D5soHJsKY0NfxxqaGqA4vwA
7olN4G8F00ztqdGYsHVQa/Bc5kPE9FY4d4XGy/12asP78jK66wz3BuV2EvDFyH45B7AMvjwOI0rz
hXAOc6X1kiODo29CRyItMUvdJLE7VQM7FF1bCkJSu/mkPB0kBYFaDfz72JIEI9ZKotP+Djg2/TjA
Os6zK22MuMjzu/i0shu11GngzW99cignVzlWLWY86yV+xKNoDHJ/evKtGoDg844uJylOSlJfOXe4
gG/bgyHvbR2FATWUFakvq9BDlrNI6b2+znLBxEk7CPWDJ7+qW0vPP5hq49FxU+/DNzOqLkCu9sJZ
bpELZMT4SPadgm11KGgNQ0ajudYZtG52RK/eECuGvIWkWn5rgBIcSBS91g++9sAePdMw/cIDqDP4
yCS0qsgyJcD9WBjJxp9bmGeXia7U3sVcvc9YIUeGg+4CblBFGrbqV10Qs4jLLLZfE80nMPipKOI8
abgdiylxiPu9SKLzTeoun0LRGGOQ1ZszLeYQ8+gmgiIzVgIgNqOipCPokmmJ/dg/1rhhUj2nMKQO
zQkR/z/txuYxAY348l5/12KV7YVPzfWHjkfhWLltYiHhEJAqsE5yblKj1I6/NE+/OcE8jk7kqACf
vKv+zt51hEv5Rudco7479s55r1Cd96FyTbAJ5A5ctsJXtib2nAHTnH7FYwuFROXOcZmcO/tBj1Oe
J0DLU9mTeOpHZuGmZ6aMATjsh8sQ4TmlQJcrdFNYoVWE/Aq1DxV7cJQeVAWbQQvmSoBbdnR1VWYS
VmFpJYY2QJquXRVfb5gkUiz4ZW0+1IOpJu/HxOuARznyW8FA2kVEyV/Ez1Yp11MwP1S4C55FgC51
d+TTLqq1TzQ34nEBwdEKrS9h9qwkrgaPyCoAMvW3cP8lo1oXTDPS0pUIz3jeTtfHDGohGr7iI1Lp
fkEeuKx/MrLvhVm5Qt3kz13VI7PN3pbHO5oRvXFwR3zDD+xVMDQTi0Z1VOaYSYMUPsVjUaXIGBPb
9lOit1biJwgaCuc33tB2Kwo4Th64AL5MjFYykoHMRS8mEwU7AMXtPdrDPdE+5M3VPgqxdYER5Zn2
fm2cllSaznyoucDphKPMc8A2s5q2L0gXjkmg0ltGM9OI737nGBIzmi1Hfg+wcbWq/8DI+GWWOTAk
NV0+XzJK4HayXemWoHz3bb+KK9DnvSQABFuxS1r6iXEGIwWNBZjbXwkIxftdWVyRF+WUciH1lyEF
xdaXRy84ugGGjDRKqqeu/IrskgHFvuC4/e5DKq6Fgxuc11K9VF/MhwaB73xtTzuGHWbREhSAfoyV
twLfPrX9i8nU0L57DTnWZUJVqXyGxldouGDb75hY4B1lcq3DpZIwVhYjCzRkbsR1ciKnOYuQV0sL
fhgqEw2pwAW+EjdS/3Eag9apfNfa7YyJ0cspATZwhy5I/nWYMfHdxGfnOjDPq/CQEszHs5wpGTA1
DQpMa/a30M9dfcJYjNCca1KwoNGHKVHKDSdf/ts4KlRitucWJBV8kFAEJ8hBkDLsfrQ9x1XWWcCv
fk4B8SLFl2bGNPYh4t+NNkceA9M7DfR9tKm/grvaDqk8oVkjeQz7Xa88XqA33VNICtgb+A04y4/+
01DP/XbUqAintyBwA0TgL/63LSGpwwQoqXenUTkRVcoww2SoaeR0dgTGDHf2HPRTaXygCP4/8k3m
GD0jJoZycO//tRNvjfeMvOEzzct2criWAtZM+HPmFdyR+iaS9mbAmu8JbqPEJzngDvQFh/qSIQ8D
C6wmiYyNwrO9xc4aweUx5YoL4zBW86Vaq+9GgpBKZSQYuZ38bEyJWFVh8B2dA2INpwwdJTEaiOxA
jzJMWwZ5GNmPZgSos4XM6Qqf4Mze8LxGyGWRc67Zy6vZyFo63HP5Y5x5kuUwxPKVFkab3KlHXUr+
WvimQISOmQMplMDtrXONjqlhzTqMm+u8z9Hu1EyK/1uEf7L/pjmGXdcnTwoTiGaZuDcGGevMP86H
NYLaOzW4+fo6+pv0IuXm6ULl2l4XA4PMQZkVTAm1/1uQR6aydonyi3FotIaejgC4CHFDWfhu/VNC
XTva2YX1IwPCwCpezr7n0nhdqtOfR9LkVxQBKpJHTJOmLbmDYbFf8b5/kvbygyuNhMIKdYjN2h14
HHkjHhMG2YVih7dhdc+4nNSw9dABspRjgWWMkhtOauYzbH0xkmGzDOJrg1FMREGW5kpxWJq+zHpz
RZ+GRcKrF2OL14LVZaTjKAriZFyTwX1Io+s6Ri/6E0D+PqH83zModowKVHAN44Cc65fq4tAl7uSl
YYruc2sWnl7F6gWSGABpIr2fXDndfi2LjIDuHIpRTXOFPvWxeqC0URddwbL02LDKi6PtUjaTeRlG
9ab1ykYhAywYPML1wctE8oK/QdrZEQRv0TPHXxIAymLZL3vYmIRBUiRZhERR4nBh84+VTX+hODZH
621Tylojm0Je3IqrVKP8HvpCn+5f813poZMF4TIl3dBJ6KeGqTIfsNxppZjRPQ2PP6qV65+1TDRD
9iuMhgNQzMWh+S2ZxAoMyl+tchhmcjruuId5J0DI2SXfjbQzfr+ZefR5woFUBnlUM1YfrZnRbn1f
lK7Si4dO1MHAmqV4w3roNuIo8Lrzg8+7hOFaenyB87/ug+3A8MrWV+Uk09cJgqI9Bxt2t1GCIC1J
SF3qVz2ZKW4tHHlAAROaCEiCPeJCqk+EWviMYNoqGo+U7wrVMCY3XUrZw1/0eqV5l8UHX0MYQQSW
bAoaPUm6BtlIGrbk6c3tWtb9RmpJZ5FgAqZYx+O4Qj70ZQcu19ANUmtWDiR44m29HKBzPe+5h4T4
vQAnMsmsRlHNxvZwYzSOYJA8eJHRDgLjrohV7o3/IRGuf11pwNavhhHjEfOSESfNMJokyed80Jie
tUB5q+xOjitj+j1bt30LfZGv9f57M1p6lypxBKvAGTbHDa4RsXxlxGZV/GqLltEEGnmhTiC1M3iJ
D3rkt3nzWogJGnEQwpJUGKx1jFLwIOVxrSavKrPoFtIbGl1PunCoyvv2OdmoTwnf5xihvo1Cegrx
mPN05/v0ohePQeXhZVeCYvEsxURqaI1Jzl3LOSa1ktD5HeA4NbMdp6YBxzVpQ6AreHqLUYNpTkW9
xIrUpwtPBVcu+4YyylnQw+kISnd+dz0KyBnx9amWIce+oR5oXPUmHtpLd0qn5zwX1m+syb41DeWs
paryyFPs8usx3EPtAMLGSGbI+YIidSeOYztQOUsoNWmXAOzhdHNN6F71UIo/pBBjmdWa9KSPvoRT
GwLytjFeaIud1s4J/TXafEoNIUUtyneGqTysC+8rcd91EuBMpcYmly2MutYo5RCAQMO3F+5BGtY9
jy7WrOEBDF4fTQqNyakYE605/XKD9NASlAbANxPHrBXQY4FblDsohsYQAL9xm2Iexm0IUA3rGbPU
hiX3S8m8VwkwWg9+vOUiBszzdXtb1tHYq2Fnm2V2aNb6e+bmTuQ261kShLqnJVZcv5bmkmgAtZE8
4zrmKK84/qbUaluj3pQQbtp0e1KlK8AnxKDDRBdEEzL9eZq9XVmbtAXTIBMxwLEV+HV2WQRy0bGU
gV6/OVDBCmkI7TXuStoMBqflmzK6z2zej+ggfqW24ZPh4fpbSGXhrZ+31jd3hE6ZuwHbx85I1I1I
lcok5URlHUTbldj/f26bv0sw9vd43ab0kFc5ep5/+yerFmNka6n3XaUp0NPVDBX+Ujp/3AyJ1TuZ
gJlg0X+dLyd/J2Rd63tH9krr8YmCjrjm2LsoGuaLXTbS6eeU7AY6VxOa7sdF0twCi1/DQ2gujEEQ
YfPDJ7uH0rG6nAUH6XVYl1WMXaFMs2LsvWfJepYylq2vGtiRhRWK89CC3JDze9fKojUt4W6q7CIN
z3pmBz2rgqkgHd97fTgKXPORLwHHqi0EJrYt9BclpXJNgfyO3Hpi1UZfcPViz21/7Qlj43s0ReGE
XhIzpSFWO5TPihwt73kQycYCzfs3B4aNoO4ooHirNlrYJSZn6kRMiQJKdW4XlRCkKvkJEwdl7PtD
iPTgg550Ut0WRNbHaRH5wW8zojVmM8P/Q+5qGSVr4quesedCDiSskrgdHgL1qdolwe4yjBWjs0iQ
cdtFeEuR07rfHtoBi/nokD4w/Z3HYpmIZWqXjy+OOu5zEY6L9pJfvh9k8wn4wfMDJHPNGOrXPhXi
sAPbgV5nLs0M9s4tvV6XGSEQBZlCSUHs/PhSnpypiLTjiRVxHh/8akh2rXCKcAAoZ9TGgIb0vSNR
P2eFaYTdOP9CQeVbRAB7+DtDEW8aABg//HPl4Lc1WwKQKkVXL4SB29Z0+b6PtOKEIHYRKOJ+i6Po
rnRBudYZ84MVXo0AeHQo7MfFwXBUTInAxOLk1skULXeGn/KKAItvp085m1C3rXsxdvitLZqw33MI
LA/XOoG0LpT0zJkTmVzCEhB5aAierNMxiw4Wl3L8KhVZk2bgUvAdjSoM53PTHJAs40GmwYIZzVfv
zcgJtV+Q3ElHg6BEm8KwAfG/OAANrxyF587ky1YYaWIP2r0/1OwPN7XICP5tXlks0zDEno0zWbqr
O8vp2WNDlrTh7mRri4HlNk7OE1lf5hlO+ry/Qi/LbxZQaJR1SG3hgCcTAD4MaBkzQBqHVIjkOOaY
OQhOit2DYmlI78VSDP0p9jBidEju6vQRdmKCpc5POXgtL120vh+N5qVXCfk29vvqoipPlyGCaBGD
uOvngRByhtKIbrZr+/fg9tB+nQo8sKxqNzDSdVOPkSpayAzpp0jLPX1oI0E1poQhiYx/AL+hspxm
YopP8xTv8Nf4E1E6LptKlZleSKt2qcqwh8BB9ub1txLHzy2+JYc0qaaSNzCB5ae7XMyMsilROX0/
Ggq5A2PXZ1GJEuXZ+JE9T1yOc/+uoz14rMbV5BIwKEOtirR3fb94enz2io80WeqcJ1fFZM8KUrLn
dHWCI+aoLnouLGEwS20+IgUM3MSzrQRQt1vDFW+/UTVG8NihMnAY6dmlIieNzmCSxxjLXqVZjk91
Ek48UN6CNqPBWqc4k1F0/js64hewMn5WEUNG7cylrRFbkmIfmSyH9ZTGmS6nD/YMwtlJoycGhBnN
ibaOo25UaNUVQGePlcfeW1n6SkgWlAXFK+l9y5WPvfip1dHmoZPxPLXLiAPMugI3LLPIQNZgAoSr
Me8oXTQRuSx0AKMVGosSuyvg7WDPKb7E34r8U3isy6y+9vlmXBIfQsv8a4AhdidFmFJDhCXQLa4A
PG2Lr2KnVOvEJEDOdkDlIXjFx7ERwua7ykIvHN2qlOAbiQ30f06t+MXMeBK/KFQmrta3JIvwP2JZ
4NiAdKZDYg4p2ms0PMhA61bJxQ107KhCcz3SSDLvSdtM5EBg8GAR/btKZWW7YA8NanQH6yowDfmf
qkiWFI8RszxRZp6irugA/PaYRDRhn/vnacrnFrtTU8FEJxXHFw1Yk2mqoUK/1/KxSkCs9bOaFfwC
G6QMHoBzTzmGLOaDi+taCoB0C1tcb62RfPIUS0XpC4B2trgUmULGhkdAnUIuX8Pgul6qDQYziwwY
TrgrtrZFHQ0IzJL/qLIHGVf2H6Ow3QrLGtb/9l617Cvzo0IUWZ3OiOw3VLO8mlakFF4dVLdyGXqP
mjhywFzvuEG/RMq++n2ngywcm07lD+B/X8IA7AWtbtx8EEP5+0PoNGEM0teWnGCLyMlxpah0blMs
pIw2wncsS1yujhdFGEbOWE8PrqxVjOJ11f8BknWoIIt+nYseH7vGJAsJota7OEPmMdJIB7Jd0zQg
zsaV8u/1XDVEj91g7giR9X+eAa0opjapM7tYcrMyyHH77SxpYCZ26eW8i1eKT95/vfD4oXZuLlHf
YvtroDNLyEIkR+aNymbAhkY0csci7Qk2aNVAX6+Spm5STNNyuZFoQzNta3QQ54jSaxJZB1BDhwKB
r0oHECKa9RfGf5X4o2u1lx8bfQPRNP9X/rQ6iYaJTLbcV0mC8+Gmtnt7FD0QCppFXnGWdI1fZdga
OdRLdZtnZmC36iJaEBZf2nHCaCd/Ev2UPGdfouNsM9tdmHxt7N/aAlUzPYOKNm4gYOpzoU0VZXgO
foKTLMzzyTxpO8JKcvAg+Mxr/j4sGMujAnCxsdAUQ1YWZ8pnPS31PI1PWm6NHR6PtO1iwil7UzoD
W0GNGa7ZpUH+KYndPTiKMYSStNB4Bu0i8axrv5kYgNRIGfkbJwT1bsyZf/sd0QdIM4njX7ru7+Ua
LZRBsefx1qRKDy9bCLoa2A8gxuZTzcRzph827pRHrR+0KpV00KdPTaJt2LUmOxmes2CajTA9gqDr
r6wLFO+zrzeU51VFR8EnBSBJz9asRut40lBpBTXH9qgo0wy7QYaVdX1uWY/v47AmGbrZgnarseel
1DSco3ThMJeD0O8c2i8+O2uviATHINtUaTwy5Wvz7CZQ3Im7D2KkJnC6apocSoUycstL5S8KkyOb
N0OaKk7P7onyS5VWlWqti6n3W+b4BgYoy8rJcCFR1VirB9wjCA/7/moOXt1ixVgKzQv0BuWOx96i
MUnEDek0VTM9GurcMG2kc3KpV+9dHWzgeZ8jNGcZlToFnd8a12ef7Q/B1rREl1IZop/M+VzLlU/n
8KseEySTC4jNAMsam3vIDCMsczvmRdBhMDi1ruOwAmqf8Qe7Km+SOLg6dObh6nZgHCB8/yMC0pkn
3AFT4JL29KLOmS+sQjrUsgeOBvVJFw7Aw15GFfm6IY2Gzf4OuPI91hyNxnO4V5uSyWmg4bgAhoYV
Na5KGP5BFEax4zB+w9RRFPQHfFPU4g4XTfOkdDDF0eBxSywA6GfOmWwYLuBbZWr3MMX2Bbp4ymCO
EVzeDN6dGzfZsP/gYKcRylQqRDLAxt5M6yDHoX6egWvKMVrrL3sP0HRhw/KAGbKklX6uhu2QLkS6
QvuulpriWXdJpkKoUFeY9DLc3OgjFih7Hr3TiJvyLaGPOi37HXTyPuKhMVj7rPmjGNIfoiYcaIw+
raz6agjoY2qBjNXEICoTgozAHMOGfu99r5TD3zCcQil8suRMLO4UE7ShuFwLKe9OBFj1YOP+X3Ov
708Hf/AEf49+51CWxh3td4hOHxQDP3Ogi5FC7vbYWvum+qJ3jRzoYbMrkZuJBYOWJOWsbLwdpzqO
Ma/s8Yj+n8gMzHxrXTtNaTJ1LB8KZIEnSjjkiSk5aqkaVKAPeQ7W76/QUSXcdBW9AAk/cpLvL2To
DjIULTFVlv4MN2za6VssPI8Lz3S9H/YolTrB/yGgDEYLiKgHZL7HSTYsRbrMqsj+8jJ34vSRrZED
KB001+txBQEXY7AD8qZphPSZCQXVM9erd4gtRXKJFtojYWiatRW+rcg7qThMnXf6q8g3kDdPfu32
I00xkDa0Jo4taUFFeYacgJKsbRobnIoOZqzobiIz8Qhr8h6balDUy+S3wH1J9EaAJLhtLJpP4IRi
1BwgXsXVPbCwjTS/mLWy76wpP9GyQ3e+mLudAF+PgyEiuEGr9Sf4en0koEodBBTAdBvamgNxOJgz
DaDH3VvWxDBJSKNKZOipfpZ1/PXLvGCLGlJvuSw6K6BJOggkTsJ0VQIiDadqo0qaTSov7Ig4vcSh
ZeX0anCgSJaZRqK9yr4QnLxH6nSMzVZAeRyefGF85noQaLBtfiDqTWBl90rANT7Ne1Wy2kfbugLN
8ShyL3skPJaTGC4JufeMy7MK7TUbwkFY28Q29VX2ZM+mSKLfsRlPZj3eMFOj17nJ+GT7HJwK2Zuc
c+WYDwZlNEjBv0bW/G/Npq3o4DPAaUaiuExIIfJ7WYJuFa3UKxxRmBRId/WhLmeDEPAD3R98kUgn
aixUivjw9r6Tc0oN0cV0CTfNjkH6qtkejTmQEr3xHHgO4E2TkV/kTx4t5woTXFKkxitakef80HT8
er7idp3fJWGzYUSn6KC5qw0A1mLebLxTRhqpTTZxjFsw6ll1ryhxPQM2OGtJZOGzWbS+GIBt+/cX
wflT/Frg8Ba+c/KmzplB4PTduQ2emdmvi/qMO2Kj3twCJQd15EZNUHm/dVnFUs1G9mLGNWmnZJTU
dIsqCQVD12wQCwJZocZlh1oFXSW2r3OLu9ezeT5iO/0URRnKaw5QyZluS/4NJTfAjFTeorcvwFwn
QYjMKBDefFkOjSRcLp9KotCshzaI0i8ru78jlEJf3X+mJxBSYmr1krFUs04ma1gt+E0NfSUBnIla
FFC4DItF2mzTjOOsx4YXcjx4MGWrKn6aHsNO3ADiKv1hYxPZO2lQdaHT7Bmd8n5bwm3xiwHKZFSI
szIvbOQCyL1PaylwASou1gCdlbJEUnmteMhcIk65CmCUNmF9pPmxazeu43EdRzzZiPz72R92d7py
m7PsdZm+HP26ksl9k5a+e9FFvELLp9N8ClejKriBVUeVf87tx/mes/7fA2joI2nt57nSkud0WE9A
vCKsGvPjwxNxv8mjHBYaPWKvS8Ho05fuXvMyKTu3vBSE/QuzruveqrtTpk1kykEbnHMpHeSGEOKM
E9KQqBeb5NO0d6d+hl8qouHpDJDR41MpzUcv0DEr3vlR1Kscgh2umi/SPA/9x/zLaqOHEyZlakHR
sE2NUDQaTk7FmLaqo7odbmlnqjynwKmF9lMKHCLGq7nwWRjr8kMpAx/mxnCCApYl59mtWxUFRDkH
WOgDJ+ImW+YAAoX0b4elCdBZTMyO/hAs0A51bwt0CkGEtZnY4acO76MF6q8DMOoOHmBptox3d4Em
Qb3QjjNR6yAhqHrtmgMgfYUItFq9NoLTpvgRZMkfWvPvhwqFZ6pQCwUWSj8tH9zmpca6fYrhl9La
45EqXqVbYFIqnczJu3TkTj+RK72yoLZdE/4LvKIV11UDv/Mja9FY29OKAJeddvgJ95BCHbgvhHrP
Xs6ULnL5u9I0ZFVAWAJDeoJLxmZUckJ5OV8HaQHRlfi8WADvGNFo0d2D5762hQMBD/qZKnlGrv/G
gtZLeMflWpRsyRMlj+I6mDqfs1OSaV8ns19SLECGo0gvZrvSpt0wMtaEJXcn00VT2o0oSbS4YqWP
ItyaYybmeSrzQYm/dAZ8LQpVRRsWvJuIsCC2Vb5sNg7PCc09Lofhg0ss1H5TvTXwGAXPEqlpQqA7
VybIyQbbwMaxgpB1n3TnTvqiE5NjC+hsgr631SNLkzsOgwycO7ta9uWI8bxt5tiMfprr8Bm/rr5x
CHmdNfgAbQcohNX2dySwxYgK0mklTU7sfAZGAviJvt4JLgCZfoYRBRsFI4g60wOyyv9WaOlibXVp
d0cSc9x9CnBva7KwasX+TNf4Np9aVZ0YPfFoM5UJr5V3gFxvpUB2iP23dYTfSahrV/7hEXCqYHDF
gUdeFTJfN1AdzRsdg6/coJzeKZ2rliayP9DZK2Ik7wgmhFoWcNyQy4rDjSMYMuuVyIgTvQC2Ufdc
zTXLCkoiSNlz2l3OwhBWW/I90KkGuvi72wsziBJC3QF8qPFOJ+uDANcMcnogQwJ/S2kxxVRrXLi/
a1JHUwfi62qxwNYkBzVXBW+NekzslEGq/O1B4URjqYM4mFzffKQTHR/YSQkbOlDhRtN5mNn+Xb1l
7TTrxDsWUad0jr0apStLjLPV0r1KTWesy2VcIEfMohDC8UDit//2P4hvocTTKW8ivZCjVAVRud1C
YUPtR0jP4ZJ9hUAoQaQFS5GqZniiO08yKeE/h0YKuHmclqL6P+w1PH3b5m+og0A3cpvoCxRzTBi8
n6e2u1lsYg9xmpj2kBdsXtltX+mYAqQ3LaTLfP/4meJ55/6n9AeH4aE3UxOUQvngnLLbBWnAXnIv
sq13Yq2bXreu+GgVJUs4C0g7D7nzMbUjnQ9ipqi+lcdhimGMbRZFZRZzl9KLmJmbGpMj8r6r+JFt
bVRdwzPAp9JKW0G6cgMLWrg8MGa/WVEe8H7zOJfkllM8v5PHtJ5o4STIoat1gtjUA984rzQunivU
1OpEfLMLgsAmZ/VMuno+JtPIVadBDcyDpgRTyLdXPVtloHyKrleaE30f9MdYiJPXpXMw7HDm7Y4o
ja6XFfG7FZ0Y2X4cIAfv28xWdvEMR4iZEQbKXBsG7QltXY9i0KkxQl5RlOiDFXMJtgITMqu2P/p0
Q1Vb82rqc0+wxmjPDiZMojdNe/hUQsWnmhnXGbP1G4pMEox90J3V8SE8AsYAwA4eaegA9LsgXM9K
CT1bWnEPKnFUZvrkD4DLaxg6wpvZOONZe659uAo2xlmrCL3PuFnDgjBPIDn5/ad4LexD3XuZkjka
YoKvTNDrKcNPZcsaVRoIJKhImA1F2oQXzlbvU4OYoAv3jfTO8ek/IvUo6HCI/qASzxsXLAEjlIHy
4ejm+a9gj78GkKuC3ns/VJfEsS8reOvpHsI+dvCkK5nBGAkvRToIJ4WsmWgqGZn4/sJlFj1jtVVz
Mgz23st0fQBCt39UF8nvYupgitKE77RE5gkQ5kxKJC0R2fmSh0GVfoHxgJvFHhcFe9eVkAYrdZPQ
tQJkrNAO7AaOgCBByIys6Qp7n1FTocV5gNWaZ2P1i4vG9muRtlTZToUJbtKPf4MWoGs/1DMNL5Mu
NHoSwrquvksA66ALeQTjVTVY6FuDHKcCg0D4lHqdzIjkcK/rqq2Wv8O3EgxY+JIO2+TdbYvM+3uc
N9FllWYARyVnTwj8GJbjohRvsEuwkrq09mHerCrw4DTuVVubOJApQCI5VynwE+DGvwaJ/0uChQNE
AxN+sE5Iyp0wtHUSH8cLPTaqSaX0Xgu/D7VfjiXW1kqXKU16yka51quL020RgF7cmdQ6Qa7waPpt
u2LkCuUq7mRXU2gbJlIiiOhD0R/9mHwNjEDezXwv8eaXzvOCgxvFhjY5UvWa0qxkyJiu0WKGhtfv
0JaHKpSwwGew8qrK2o41vzZCpbgtqshSWeJS6oVW9G8+m72xfEYfMQlZ9KR/88sypI4qXCPQy9so
Dq4IDgm+jeT65POg8acccCO2iIHFXP9Xx6AuGiNHbzCI5SqbdYO6b4E9i1TRecDhOmNRoIkFDaYg
EqtwaRIEmFPysaT97dwycKj7X3uyW7VQjUShCoazL3MxWl2O3wek7JBaZgLI2c7zOp9q0EuO5kov
O66ex0D1kP0pFfcywWZuGMfvtRuk9bAi3+8zlJ/37626ukDYql1Jo4aRGVYlwS5YpU99XsvETEl+
OOpv/Zc4/JstRsX/DtUu5jrfjxRNhHBQHomI0DCMEEMq4w+YPzY7eCkvumrz5Z2YlXiiBiyD0Flh
JaiIsB/iuG0bx8+Q76Y3ELtK4i/7YI+uhMw00gbjxuU1f3dD+kgJPJcqggrq3pm8qYbtH6cpssob
XoXi3GQtav97AzCWXq1/IWzZjFNGzUne64m0x2anQtF2DgGnzL7wdBurQfCECwzOux7zNLhcqZFJ
mtHszhr+pmMy8R07JP8pB2FCNk0PFUEra5AO6jHxnauX341vy3rqV/8a5lf0Z2hdgz1rIl2s3Etp
aKB4Uu2i4Zo4+LYR1WtvGGW3c5ecbDe6kITdeAYR5Kirs5s1bDqAq58LJC7DcVy7Bii7se7qfj32
d4MUgCigJeMNJJDLpohPWAqU/RrYZOB81KxKccXcfv0i7vnaUA1TrPH4tzC2bp9urBIQsFB2anVy
MpIQegMnajSI7zUnU22SKudCYtLgJwF5DAyaj9j0BGiVZ+YLoivC1+VQkznPT2wfpEmeNPqEFBfZ
GWZgryB5SeSQOOv9auHnh0mfULUJxFjfLiui2FF5k2luDO0y+kztDdMcqOvDr1sOrYr8qBauZb2h
qoW04XZpbUVjhD58ViBvUW72RqqBedvlhYxSI/+CiJzK7X55JHPnGsSOYa+stsmtjA7le/gpufu6
gSeZ21dzlwX59INlQU8zTWI5FWNN3oib6IcuLo8K5C4DSozOxsnEaJi7WE7BJO87nyvl4uetgPAK
Q61QUvKfxN3a//ubnJafB0wkB4nkVtJlz+C/SpKzmxz6nM6121oUy0dMtdfnPfHshRa/dWnYBsRv
q1cJBzUfqMKExZdmkLubBtpyXpEty7NKaqGvWG7TrqgcrwBhMueIkxWiK4OiSkTGc5D4xShRLfPM
vaBW/tSvAHA6fdeovk0gA1h2OlE5CJsMhxNgExAaFNdy13Voqx4U/zskW/w9qgo313W9kuXg/wZ3
LNP5Tv49Zet4Rz6WtI+kK5ZkLHw4Hvon+cMKDfM5nZoBat2vJIxaXal7G1enGWv8IJCxJ9gWLL5o
Szf9mpsLCnPfrzrluYxypywjpZhbcwUt+MZz6AIt+OZZQ6A3FXlaMEulOsUz4zjW7EgvW+SVkxSz
VpZwpmp5Ct7mn4QgshI/3isQRE3Mdh0i9akO0aVmn36QNgmMXuaa/Omxujard67rGwmor6780FaH
YBmJtrZ75o38m+nHHKVWNutvKNk69YrxP/ztax8HduTbQIbK1ttc6o7/P6lTMnSsbkKSpbrERHPC
fyVgqP0m9LgcB1ATXjsz/9I5E1tUVVA74us6O59wnc32XfbHvj/jkphPBmmGQ9p4lq2QVfsqROFX
Zrq1m1zfx5+5uRVA1uLVXBlqZIeiNA2+S9TvxJ/RcG39UFraEupvUWulyKChZQJu9aafvFvwqfCD
5cYD0dgPsXkW2yuuEH43Y7ZwhnuesDWLKW/l9isCjxQ1gK47PNYRH6nYKFgk5sNaNjDf/fFNNwz5
2SZ+ipKoaDsncE8b9/ijQHGHTs85rP+km8t7E9g52QMuvwZrpQlazfhz4Ls/ElQimYHAu3Incgby
IHSPmzM9RdR3xN9SXB/VfLExN0/SrUf9s2nHYO94+BrneRw2JSB1xPgAK0izmh0RAQAJ8+Z44+SV
OySIrqWhZ1tIRREtyTOikYBcRcjcJFh5kYqZXdJTuc0izd652BZ6s4ihUmobZyNd4nJBCrt6JsW4
wCkiR14ovHrDesBChi8QTE96z5n8hkM9u2cGQD1BZ0oQNQ9UYsG+aLDgEYm1N7qxevl4eIkEsKYG
h4AKE097iVYkcWZljPxz2pU8FG2+S3qU6tlmHLJammiFkWAlUUDfjU74DemzzMlV27KSk0Ql/CJW
KrJ071Mxrh35QBZ72PNxox3ohu1OjEtDbPNtyfXMxRYBo7jIeMvduuhi71TtamhvmS1sPIpcFJAO
uBwDQf8Ttb1EnY2nVL6/I6y+pWUab41kHlGwtXvF5moteCBUl/cE46ziTVHukSHF18DTnJcvnAwu
3eRPfvKm1fs4DsPMmeZt3f9qDmyU35aD5jK3IGZm9/CspiBFbpOZZDG5D2cafetemSl7y6Hob0HV
hWDjwN1Rk5BolSMyba17HBjrkGFwJvpvAAaC2f6pn4evOsSJJy5z2FLt1sHp0muu1OR1XdSuFuvX
cEMNw/9v2TBiuMmmvHm9u7YHm1Ejr2rU89X6Ez3Vw/CX5Rg+RhEeOFLojI/LqyaTmZuWcouwvn3F
X8p6PAbCRnQUjuJE4VIdPYBCkD/zNHtmnk1QmRZ051Z5HUXXV/9J5AMQU+/suvKna8oFKKWU4wiy
KjDluGeEcnX0WJS198aJK4iMTmUhrg2EiDD6fHetNlWrtePrzKWALExVQcCMrdKY9jOkYo+HW/NB
LJZqdgQX7XlygjD5pgsR7b9ZVlbka0PU+nbYrXQHV5tZuPyiM3KgAc32IRiEotJ3yMlSGVQzHJX8
zGivuLEdaqEZXrghKW5i6CUoWR/cr1yRDnAMnViw48Bx7wDEz4hhy1tFuLlKlF3lKYaJ7JmYn2lA
eq6jpL86EoDj6E4PGe/YuGbrYoGcTPy/Kw/FQJ4udYaYODlbM3yPCTOcKESt0hLTCeLyl42QB2jj
RiMLKDLJNAWwsAU+6RPaCcgUz7JhC90Z3VAi7Vt74EKjfEjlmGvGtpGdoAkEKJIOwCObpk7JfQDX
T1RagG2yA2MdZx8uZXiJiNQRZKaiD1pLyJPEUCgZ1hjsAcq+v6Gdqo1RKtKjwCNRsnbcEiqXe59m
WI9eSUVJ1BedraxlwWoi7fzMoNCqjaGyIDdzgIZkd2PZiJS/sNndNDk+jgoq3dvCYoT8Vec79E+k
JnD1pB2RK6ckmOgEkDxNtzs2i1dOVlqudlHHv1xf+F614wiRyqLXKs0CEA75H0PcS1g/eYDl7bgZ
K3iLEKd7D6dmbHtjGfWn9IwshJLZl9yb2hOzg+hcDstXHwSuRT87YPfcfO2jkSBFCJt7GJ787oI/
2yDph21UBMVVqwDRMpxxuOvNzC7owU27jyCxT9VkeZK0jtzd80Dv/4tKmj2ofxq32cm7R/5lmK/I
y7oQs8oVp7i5V5KgDbF02XS6c+1EExKP68ddxj4xNvz5A9z1qt74YmbZmhU+0t05+/HpvZGqRLQT
bJzaftNlHm67xRvmOQ84f0e/YZ1SNkQCqF00dlj1TnYUxlA5jZGXSn1LPHdWvD4g9Dp/rAsnRV1E
ZyqZ36HB/zfc3pUzTbPCNaewZPt7G3Fw4UbXtNjfwgTmuBVLQ0GHF+Q8vyS0v7O61JBTPUpKaHln
b5yBWHgDR7h+BM3sBmzoWKUgJJPQGXScjIB7NH2cslNVsZCafW1rgQF6Tk4StGbeU9ZeqzgpeX2a
Sk/58nQJxafr3H9zTW7DfP40M6s/sbeDlzPrC7xqNARgnyTo8QwHPjFQ59xhl4hMKgA/fBAemb4z
FJzmanf+GkMY+Nisrf5SJJ4CXMh/TYPHUHe/uAuf0I+wAiwrFs6v7a2I1CwJW+R3RWST+WNwaXSA
yVOiMv6fKcbXYyoGGrvmsn04E3m8lzXA0Sf4Gv0WhRK4+8qyZH6reufcso5Fd+roukkavrrDKKBh
9Z6y798G6BzRhkP2tqmJIpbRg5goF43md/H4Huqt3QGVecWL75dM9nt9jz6uxr94bZEkoVwvfTHa
QiUcyeG6cKyqKamBawQ1Fs3Uj0Y3zlEjvTpf+bne9Jh6ygY4VoJg16FjdRO8zsoiWLPZh+c+vmIg
q5M/guLGq9gRYjohxc//ekG86oE/4evK6fkf30ZG1M4F1ZJztLTRoHGFW5+td/WCl9uVH3lyKp2e
/XhxEgG7+xqaFGbIOW2wUw8yuYJ8gjhlENmNOgtKRWate3LqVWNKRrlpmP/yGrgpAeLK78DKsrdG
fA+p8H5UHOSgymb7Zu21/af7x0JW7n0R9/VfJD0oRbPWSTa3Ky1dfPNH+hi4usVeVq3mVXGlbegR
P81BeVlSDqnTlU5eUItxVK9ugn1iXsfuHDKFTwKSeC93dGxZYhxt6ZMDlwu3H/3OtCgMBN9lUON3
U/Lnl+MN5vkhUsdj9KPkuVlC4QedvOEYb7L+R/6d96/LBXhE208MVg/izKzU9HAVrSdZn7+Q7OX6
dkSgBtB6Q+RRjtKgTmhkjalLwLFklb48MWO18sfE6wOVxTvWjJ8rDytYGA7nkR9eXWKt13iAhsF0
LKg646j+Rt10cSFXWySwZif14qZEHmDi/JvTE5//5URQfz9zsMxhXYlsU6iBM7ki+zZz2dwkcPZO
Lp+dQFTxcee8+wbjoTIzCSk7CUTuXCmcJMQei4eOSJ0s9gnma/2zGzzRFCChxxv30Quj5sSI6WoU
d9etLMbESYaILroj5f62dhqfxrh6OeHzmPzN7M7q0Ro9Cb/+7AqhYGoXOgCntmB6YOzxUOENXZnr
m0BNVPXFDpNZVopOJ1seWg/Z6qwdVmhGPrHMnwPKkoNi7TTopXuAvmVX6ymKly1VrcXZgcqoWHJW
l2s6+lHFDKLsyYExKnjXunMHivCSBCCU4l/e4FImZWLf+Dg0IebsqmG8z6JGj3Y5/qPpPAMvnSCL
U22rDRUVoqlLSNIWLu0B8HKzEr0rcadlz68yNdAtXq6zF3ZJHWTN6fLTlgJakojaH8FduN21oTRQ
Y0YH5Attokt9bJA4U3CBrpcaMYLu9IyqmKwzKeymhMi1UvpiJwwSTlso0LePbUglzC0MxrEweIQE
GNrDhGsx18VWp3iTpGtRelL7ali7prVp+iaa8pnnKmBXt25QEiiLpKhct9dWauOcIggll+dSClfI
ZXffc8Z7rPuh8efm+8dga40vF50T3NNqMYnTdeglMyP0NKmlgVE+K2u9+RGC2v0/9QmxHFjD9rXL
5C/LA6dl1G8J6VjunuxLRFxnl5VYoTYcgFyCvwKOqXD804FQIWc2Hwk3rQubL7eS7RpA6nhd6mmy
r4Pto3YUObn73ZJDb+tDTM9UzhOivJ0qkR3UigpaEWqnl1v+4x7rdG2xhk99NWocYoNYJFxIw8c7
YNO5l2l+952XwNc1fAqb9/i8c+UEDdZQg1qqP5azh1o21Wf8pB0rX8nO1m55ChhHhItI6oew8bg2
2NTmwOICC1OZYlGJkCuxyQyS2Q1ZCUcHZCPYcTw1GQD/vkodaI3TsHL+E5xTHJsatGDHrx9CEYiH
i6hJM7aQP0jEgBD23IGOAR4RsL50iBjXPjd9f7q3jIfzZ6Nf2wxNY1nZH/d48FwNxvBBakEoZjjF
FMIUo1iBAht+qzAhKipU4ghcwYVzLE0dsy1nSCH5BGM/PhEaOPMiciQeCs3sR9N3z2jjKM1R/gLj
YKXEh3jQe8V1DvWY94dkW2axuQcXu1HGRL763OoVCQTh8ioCp0BoNs7f1muDqPjU7hwGyZivAMzj
1fwC0QGIPqWs6o2s3NUoN1FtbIXvMKtdTeSqAXSWIHuTc+G8TQaJppxIoYmdUjHkms8iWy9QZMEy
L3sHn6ck8lVJFAmtPfIA7pg6qSj9PLIG8Ezm+um1FgFT2FntfTHdXDcqR2HRHc98W4O1iyN0zj3V
BEy3SUxPX6e709TlkSEOoqjArSvXRUaRq0ekMvFwuw/OXDnsnMMF+dAHu8imU3RIO/9e4Bg1w57t
0HRjZSPp7VWqmrhYn5WLN3PIqK/qPf91u7sojUVzEkN0vHt16EjofJWutqN52nWlvMc+6EwMADTm
+47zKO/tamh09BrkmuDt2GyXUI1HNskKaIokOpkDuoeAYJK/QUCgO3+Kvmck/ZUY757yzAzm3kWC
b8e4PUnGvFWTgPA8gLBFUv7ewm2ETiK8gMNOuV9DxYLfbs/QKaY6aIUgkghFTJMKBDlyODeLnf/X
MxpfqWR99ToIAbc8oS+B895ZIi0/FCCzadGaINdhS/0poIF8KH13p/LNmHd76Tsi0S6DJg3liTO1
gmqV82AFhM7dn1PDwozZz9e+j7YyHwXqZrPNQfyyaT0IshFfJftiT7Ynm6cfBH0kFuk30SaMOakf
iYSNIBaRG2UvH9yEQIne3Ia4RJAhK+93eNLP7wIHdwnZOvDPS31TBsNTgNXe5g42zSIEGlMylRRg
nFo3IMwBGvqhqsdOeyJdPrPYi1VApfvOtl9Se8Gr0Rh/ZGnWbS1cWhYw61YMRUjKDTLfAFMB1OrR
1tyRKnW/Bd2M5hAXjVE6CwklqSD1g2J7HumobkQ7IeM3y1RXXxVS+LPhmiY3tZ7KRG5pDhtiY0zh
YD/hsK+OayBibSNd+4uSGZe/l5j4plHEhSZp3g1usWn3k6F+LnZTkpbgWOF//hDNik3CRJ5G9JZl
XAccEtk28Bpo05jHMvwHqHa3Vrx8tUgPPXP4sRzYBqSXP2RMWjWtAHspAX4DDPGfBVg+wubu/JsX
33bjSTmsbXUmG4aQkU6Z/FpnFyP3ZxJYoIleQkpcBiN2Oq9B8ZSlf60ukHjuqXL3iCh0pRis9K3a
og4qTo5pG7LEsvJR0JZ15oZswK0uJAvLIRd5oqdhgMXR40GkdG7GLwkimUmCxy7o8FUHz/86osbK
lieBQrYgvzAd7SPAHkWb9sS3enFFhRW9n2VO112SbBe6xxhDLztokihivgx1ofGbzRoRVW4WjIdy
nkdjQaqe7uLOllJ7/mTfFXyiK0IK5l2YK4/zz4gHPMTDUVYb/HLFG5FL60GlPz23ZUD7alZihgdT
QYajS6ggVOB8BurdsdMyda9UeD35Z8RSj8Z90XMYKAOoGn3jzZjh2xslCuZu6xWwpzVwpkwc2nru
uAFoEosOuwr6AWhEES6inr8YNzWmWwFUnASGK8qzglXaklTnWwbvAeFoOHxjDW39FOTmIxjaqsS9
LnVWZieIq7Zm9Ylrysyj3ikR9pGFn1vyjZJMShYtfvpW1j1kYuqPHOnaOLy+4cyYqQr0iH5WjBNZ
9+lv8WdyfSVykoYZhhX9Q/GKZfkwEcAN6M/KFQ2sLfDh2EV6rY+LMHPAM1ym9yR4mBES20Zaz5qX
vTnf92g7h+B6fkgme3ddYB+UZ+ZkJUeR4n2AuqdJv5h15ZHQdYF8oKlMQ/mKYzmY6z06ORhwi0lU
NZCbD+gRoFKpqzEqo1Ruxyn3G/bC35/WgbBQTMLGCckcRjqpAMsQtmxhyIV9zuqbNaXfX558jJul
PEXJvKoEfxGr/XFJ6RegLv+Tu89msChr8zvpfGekvUj4lpW8QWfuAi13UQI7kqE52AKqGk33l1wE
6PDEeH6EiwxU8aM3oPcTqNwGlPnVtsZxRWTr0ZCuiDbCXskvv+myodLRpMht54/Tc0DXmpANADEl
/r4BKBNo+xXgFHsDj61B09bH19CNPG+ci5yLIynvgzTmuZ90X0PYTUsXD8PsG4AjpAPEO+RjhFL0
k/uvg8OzwWrzVuWlpduTL6v+9hMO9kbKx63Odjt1MH8gk5uwfMgq263jhRls7XiWjMnhIyGntKnz
j5mTZHEoCnGC6vOk46STrzSpwDfTd2qjC/LMPTfxHXGWQC8wlCc32+NPuI60ecfXLCaACkiB+HZE
EloWueY9oPWLDYQgtegcwHu9WaRHEU8Op4DFcItGxWqSjglEcZUQBCZ+FqR0iBwJrdkQTLAefa4S
e0obGGlI7xoeuWLLlReEmC5AxH9SSpO0KinJ2CTZhSw+/h7etPVqZzSs/f9kN7PnU0jbvDYWPvAz
Lw3NMHmXSROQ2AP3/TmP2rx+n0O8cPxqibrKlzX1eULk3C6EMw7szl47W9+6VmtyaAVGZBRRcbAt
Iylt8HQmtSS30NAIr/Fh3i+IPiojPpcwVfaLTQycPWYmAq4KCL9ZwDPHRV2XvaIkNPHokPcR19WQ
+K8BE3A03X4JE7YrowapZJ2YRKZo+tfqTZF2MQUYNonkdaabdL7Uj5XAZvWAEQkpf1+xZFDE/euy
RgaH22xOar/pNan0zPZ7L58gKWyTCItw38ew5sxSYBRo+AsPK/tC0bsrZYyMmUbmCumotU+ZiDfp
lLlluwvuD9Jpl0i2WPRfHNP93PCs/6gJviOy3QrhvkqFqfm46wt7UKA9nbsIWnCf+um+RjcJbdTP
RSHdPW2x597qE/uHRbtyGQCDoSfH80q9amc0MPiIL3wmrvcwi70l8x75WG1UdPhq/TD+1vWSsp/v
lE9vHLPrrcwDjeL68T1mBoNFaza74FRxxkeSDrMWvK3cLGMJoo3VUt13DEZ4P1BYHVFTRXQ5zPVA
DyxQMAr8KG07B6OfCp58XFo50+m/06K2LpDL0nvyYrUPDQRrgvxtNbkNB1S9qXCEPzeoVJ8xSXAl
zAwIcsgHjeYCenVEy3iXjXcCswobBHqz9QvmFncBBb1biV7DZpeq4R33pb7XzVe9fxWd3Gfe/z5Z
bJCY0N6YTt7BJ/9eif+CS448nzyv69NBhPHe4FM83fVZHjXbgVh6r+FVj1hEgXw9S0Lp3lmQaec5
/L+MOAgCYjQ2bsl7PKmY1s+UFFzjK3ug12OnpDAf/d8NcCpkRmSvjj7qftXvSMhNWQDzAklFHj0m
xgnWVdj/sgiCj74KhY2EIghNkKwN8p+JdhhNBNYHAmonq7ACqSvPBsPVSPkzSMdrqr8x2BDESaYe
4xbTygAa9IWWzhS8F1HTr77qNabBnatdfnHqdGEepBLePjdmLWd+6p0aA/zyXlA2u7zzKZUbzSE9
uhIGzKKJhSpyFMJx6khtRAwFDoXhBEUpcuc1wgrESCiWx5hInMO5iKbe7IimhO+p+4EFHjqAc9pO
MJB9ubeQ5SgsSUXWdgoaSr/4u4CkiVlMgbGXFIkWTuK8awNj8saBstkYCb+hIxjdI6DuOeckjiKN
fH5LiSNsrtShN61rGemmIsYdm9Kizf31rMrajlYl2ICYJx0NrffwPJphlpL4K9nyVsiOSgyIXGd+
oSmtUnuwwYCiYHurV/IheFd8eWY7W20lU9ZgmqtIkUkT18F+cNKglWGqIhB6O23ZXolSBqsvrXF3
H+fYl4v3GAHbDd8Eqtr5mIqQKM5wOBVr8Bt1emzSDLElbjN8hfPOO7UdA3PocVeh47JudY6d7iXh
ebKf2Taz3tUXUeTaChfu/4j204rKoOMZEee24mLJ6LZpU/nURbsIMAmrEuwBddEdnDX4aL92HnVv
fJt5RjBQ1RRw5SFh4o0HSWVQnlA01TJ9KYfTpdQbZfj8qEDg6lKriUVWksDk1fXhscwb5J9K0CjI
QTTVVuy4joi7raXAQ9KE0dPh9yChfFALzfCN9/B9ODI7gb3ySHBgDH/h1MrqcvGhYfy8USb6LWgf
4Y7IvLxSfr/5jlFq4oLvS6uJa/fDDokyePwAIYobooslTt4q8ygbdFvJB35Z0n23TNUxT+/9baX9
BLHRCLW+e5QaBaUBIavoXIOKZF51uAVa4hhKmjOV7CKRZf5pQoJga1JGSyC4eDvokJcFXLQf2Y00
Lgtd4a1sNj/8IHTiAUzhymj0ua5di9SywqFF6D86/NNHIBW5A1CMr3wpjRFRV6GqHDFPZcvkDcys
BEN/546lSoAzaeI4tAiAMUXfIQ/x8ouND3lJKMQ10k1pBuZMIr6BJkcG53b14JhcQMV1vTyVolpe
xKSz04hokDnmy7fptDkqrclZTOgTBe73+3foh4c+KdpvctgZPTcgrgrJLqdHwSgrw8h4ifRqgyg0
z4hVY6HZfXII+f7dj1wX6uTBtucdtjSDpAC6aAh4ih/Ace7S+cnpirOBZ6zrKGghRe6M+e9PdDN6
WjENRGv7mpnDsMWdCr5gPUWbKZWaMawGcGLN8rquRe+VKM/qKspjKcbpCVAgr0I+cs3YF9kVX7Sh
rNuWa0RlHNY6hRSRBDElmjFZTL0kZEj6iDX7ttPwKP/iiFEQ872E9divtJmhBF3tYUNZr2hJdCeS
wJTy/lcNMlbbYgchVH9f/e8QHSAilTNdWd9SLklhSlJNXbkLQRhGnl5PMtO7XS8+V/G1QE5r9dH7
QScdEnAXBw+8SjsqGe/UKrodIn04HsrxWh6mabApszL3HNEXMXPbFKBPlavj0rZgT/JMJIwcmLB9
4wA7r7UyFugmNaRKfrPDGnrF7jY9Y/YiuGmqzsy4SxUd4XCiJsr2/+iSWgz6Ki1P/kpu+Oq8/hnA
tvD2JHbTabjyrUK5OB4jvYfruKR0jxBy1fQQvXjIqDLEzYpEDxx0oj/BgWO4z7Zlop0zdg8Z5q64
aRvP7pKZcM8SSViTfWHGUZsuSIpYmHmp1pzt/pQD8Jy0wdeP7N47vEJvuzsiuEQGAUCUUVPrL+If
mK5tpSCv6QwsnysaiwX7Sip+Z1iEZVKlq7ZxjE2+Y/b5yzwp/8NUh5SNyf+0k1ZfGI/3zq7Ds2/e
z/H4uomo8bcyxE8goIsJoqcTL98iNLYyHwpUt8fY8qSy2szmn2Kh1YrrRhpY2F0SW4VdZwJ1SQy4
NSm/5/U57nSQRNao6Z8v6lazil1xBlX4wKwYB+PHV5hhQMOy1UxcEYt1m0MRa01xYgX9aELFp0go
RHvs2wSvXlCelUYW0OCjZ//c35Be7f5vquX8pP0ZUlkcdEk45X6Kq4b0RcWdKvahPY7oRK9ayIHI
kcIku5+W0MV5BK0QQZQbhs1p63ga+NFyAx7tF6uFb1GzEsJbj0mYP9QwpG0H8Q9wTa3m/T76VGvz
gwSC0ts/L0f65AUGpP9wY4Pa60YhNHmnwRXUAY1QdYvTyvpqrC1zvc38sGMJ5h+4NUMk7V9YOivb
cZj0ttNF1nIK1phdVp33l9eCbGNnEJnPwhoxWoFKWGrH4/1AhHLGCDZtuPVq5n+RcTdIAQXVpXof
GIbJM5MC8AhBbg2Gtz6WKO1TuesOxUuLPlQ4+98kcLj9gv5i7Nk63Lp3/iQAhU+J2j6GNrZY/gEK
fDVzxpvr8fkXYicSZmZFX9pSkMDmOCoUvDP4beSNc4XLUxV81Ove0JnGB+2W3d6XRhWGUKFJYesj
Mvq/yZJXPCPwT+31DxXzoqO9J49SE8vqhs4Y99jlnRm0ULoL7dbemYQPFEJRzqpAghEfZyNkdfv5
S1EUcI890kRknWOmmGF5ikQZE6SdomiJimPiwQXs37NQfFU9Td3O6rti4MYgVwvxlyl/vrFEeJp0
eBeSgjeUJ81EhCATSzJfv+GrhmpcrYQWIcNyJBBnm2bp8Isi8QPnh3rvHiaSL8USD1+7SLvEZbbq
b09uLZx11LNQIkS/UPxgA8KR2dacgUvVEeXXUkFO36BIJTQNk71CWmIHMf7iRAvEojMUaYshz9Op
R7x6titedbKO/tGspH6pb/5CUq0s7H6DXBJ6vXMBM9Qy2ZQr8DgFOxSMhwciLVax5EbjLvGAncQ7
0Il6CLJBunRG2ZrUhU83J5fRFcQBO12c/z9nCo/Dg84KSIOdFxnmgWYFSG/QjLRl+/gErejlITIT
F9aoynFn+bIWe+7GSmUud6Wuv14u2orfIwdrwIb7u3cJfCFFFTQIZOAqi99pfgOODFwVVdSU+42u
6WYzIshdHMk9SiDSmg71RE506KLndkEzN6qPN8+BrMTQNGVLoup3Uq/q1Tr8/RamcTclcTyyBhXg
mYor2VmiwFp2wEPYtPnLdjPefczM5OHk6/eug+5Zlc59MPmqwvBNrGaMnEWF0TtCx0OSL9ZVVKiT
/Xl+r2yShwwFXvQgp30/1519nANS3Q4tsefoxgKfDz7uBA0B5cd1507E/jETF8mi8b32H2z4MvLQ
8QJxd8qtJ56By+tYhqvZdgyiOLgPqyORQP/Wf+Eqd9u0DQnqI7kaoRVCXXiK3Y07X4A3O9Kdyww/
X4JBQ0gvTL1Hs5EXJXKnQqItcu+WIW9o3stwz59aWA8JQnDK6Sd1TS8qmmwg98Ou6lFqOVpB8z8+
hnF7Mhh5hcioAbz9lK20kJ4es2+RlgTELKzpibnsnV3hLNtBxM9WHWgNgrKjsTsbJijkafwOFXhz
Lje9Lv0tsXWf0fWj8mj4SRHralokZwbmOAoB3ECaKCP99qD1TsAUgKrZmzJUXEEcyZNwEWbL8Alr
jzxcq7//QZAJAD/J19gAYpQuhJ5/hc6UuZXicljxAZwNN42TOjBhjAkJlHuttRMExKu/rbimbrXX
0juK06fDOwqpJxm9PS0WdYFsRb/9JksMFXsF7jpVIpKedFE8gQGB0fFGG5kFqFucnc4ajKJHel8+
PUqpeKxI40ShrMVYwmrAsgVtVd316ZBZJl/ePb9JB9HwDRa+02/dVw1a4IchkIyQ2ZgV7siBK7CN
mQV9GTZurYzOwP9TYDxLl3G0xn+mKwtwklPSEQXFZkGmlI5R4tdXrwlJ++uWt14ft4bjONo1hOTD
2P3UGugExToiQT/5v7TqWW/ggi8Ij7PmfgfBQFQWEe6xG3kO9Dz7aAh4U1V78GcBiuucJ9NfTpv5
dGRBXb00eAfrRFg2gnl6hedSkTIT8kmXK1DUgtsF6isgitYb8A6e+elQq3tOtXYNPlihaX7VDrjV
h5d9tceXLX1sLZhbF0ZyaVS+e26m3aIvT2IrdsdzPXF1RSbixJOBTByyRzl1BUqmpBZ8/ASNm6PQ
YwHUnPYXR7VZqkXV8M6JLEhGjDAt2mroxuPULJZf9CIQPzrLPF1+ByLiuouB0CVwn3/ILmY4RCkD
I3RYcSliO2XUKczaj7d4+q5bX9BQasmTFQ+vQncW4+9745ZGGTVbxANnJcWj9ox+koBpv9+wbQSV
+/vVxV5NWLhJxHCasfMnCEEVetnJtS/VE/FqDuYqF8k+ZvWymg/L6yoXCE6sIbcBcD9Ofvly9WeX
evsuiBmA3MHOCZWq3Y32Updnrllej4rrEeO/g+wGVISe1Gh3phToZiQNbuuWNv14T3UJjHliD5+c
9t0qzCRmjYhZTJM/ZpMZ37D1lHLbybPcvVzh7pBhorbK6OnPxzACvRDSI/LCP5jQcbK9S4Zq9zh5
YQrUDD01sNg1t1nD9DYuJsYHb3UFRmuG/47RUXIdwdUEHIh+9z586VPWoEH/lAMERERFWCPfjVYA
zkGYecyHD0gJUBCZEgr+eHFwu9KY8aXsfXUgFCuhx+mi36tMR4ocYpSOIjsQx3gZY9EB3kOmayaf
GrRpnfDFvsKKTISmtMhhAoxRHCmjt268q4GSbMKc0D0OakmV91toorSztlE45X5JGMa0fZSivQ0D
zsY2PHdK6k+lkC8iDtMU2uEOx2R1kk+TYq3wy1EjLHsgnad5c7RK3TxZuyb0PQUMC9smZSIMdL7g
SMuxD2TFU2b5pH0Wf0scIpilnz9Xa40GSiBR+yuJgU9cn82hWYu8RIMuAtVfBJoiIO3GIJ5c7PtZ
YWX8bLcLztKMSOz/kFpDd47NA05HOKh62/3YchmwjzX/pVNUrKxmTdJJASj1eYwcWqPMs4aSDrOJ
AAHIxPtawECexXgEc8ZbAsyTRDr4r15Fae6QkAzHPGMvhGzuIp1l/FPJpi0VLTrgiSDoFAZ2NQt0
35JloY7lQrf/u+B5KBnG0i+gbbe7SFydWb7iRRbBcHwDhfr5Ci+nis3NrjtodEYJFhHfQA6oflLm
jQPHbezXJeyOntBdfDY/DtHUOMR1q5+5TqHmVcNXCnPE7bHWvBnHkZ28MBbvthAPYGmhQewuVvl/
ZeTCSa+Rgb0vX0GmeuRRtYk5b1z/tHQmCpoyYnUbzkEqQwwzEnEWj6WVYOR7zQpYm2nkH9CG50wu
JikeAZRdbn9RxDSyZo80xdkSjlcT/s1rkh21m4XrHRHP+bj7ICcWTPylG6lNRM3pPnOgbA/9T3zO
7NMt8NZDJEE76PkKScHR8uvNrwxnZRsjqxQdvF9HF5kpNbsNx384Phjs3Mg73fRirn1kGXisqE4g
2RVb9KpsDu0EGf9tuN9EKOovy80SkJrqxSQahiZaHZJnha6eiGaTM0BQNFrpp00Hg/5Ol6DUpwtA
B1FsQHV+DjREGenWiLrs4SjZiSPpHr4cVcP12FN/EHgkm3bRviSck3oT0l2kBFYInwMCrhuAsKZg
6om5UPH46t9DLdTbbFVwR8wTFjVWcNsit5eaRXt9JrK0aCtc+1132rhU2keUO4tQR1ixpKRkIr2L
7m5PNYUeHafGPy2ATK+oBI4pPaMGy8tYo9XXORuep3VVw2hD+B5Z0EPw+G+pqXAgpnPX6yzONslC
l2iOOySKA42PWANY+fj3Z9ZyIDdcxUV+DrqvsMN1zvWvcjYagjYbtO8cyYHLVBJiXBacWfyWzCeW
cT4pSG5XRSo0Au7nV9qaLIrnobD+VotItLC8w0P6Qlr6u/1wRbDfemwVQRkfyCTiH233w1TNGYiO
d8Gs3fOMV5g+0/nVxiCHI8eUw36Vfr10TJwVy7q8EZWShRBr4d9ZrDQiU/NMpzx86ZRpxf6vtnpa
oE6gZ3w7d5+0gwwi3QjFy089fQjMJjR6leMfMIwUuTK2U9/a3NHhqVt8ztEs3JkNglOkZGTWg7g/
1j4PtMbopIrFez/9GNAv6v3WY6Cs/frzuJFyTJ6GHsUt9oOkOx8n/LcJcDJCDOn4NLrLhSoF74Uc
PbUNp1Qyx2fvgNGydjPbTZnHLCc4GlEOCndFdkQAnuFoedSdXqbuRNpa+aSF0j19z0CYRp6R+4YF
0Fp1qr+dwPl1//xsyJeMN/06rzEQZD8/rN1RyzVUrmDvfs+OR9ySJU1AXiZ2H9eUFnfQQJs8A5sv
GhvsqyrBsytnHj3fKdepO36+YgrNdCqMjiDxseSBNEcYBozHhzbtdvvGhXH+se3yymElrj8jqV1K
KTnzkTjzcrPFhcCSYFMYYIqQIWjqgZEY4CzIALdv2cAIOE1xaVSxe8UNba4zJGX5Q8g9fhupYx2w
v76UuDQglqLWzcn2pH291a5kUiRmX7KDOnRdKE0PWFFVSsLoHdVlWbbmiZmUXxfOcq8KHUKV7q61
fGHMyUPWfEzjCM3wKUdLRQF892bLpWe2+BfSUvBKMXC2GLg0XBtSQHOn3YHEYz6qt+0aIj2obkXf
oAcwVpBc8yUOl5tOaPDn4dqOGDOQhcWYkHupOUTSVOdaFKE27N3k1BfhVEo9Y7onlZ79XOVrjSNi
jjmEh5wgyC7R/NcAakH8sUYCs9RUzynlQKMbN/34mR3swTxsyj8DDGkoYmAXf4c8nNcUxTu72w7E
WY1ceAHbfhiX7rBsi/zK5wkMIp5kiyV5k4Cm3aysCGBiKw5r9E5xxLSMt2V+ht5xjbDI9Pyn838n
bRowXhJI2b/AjzfsfKGy9Xe8hVvCZSpjhylyy8+d8w3z0FLep0D1/kfZGVDSlTb7psjmI7PKP1sG
9+8Aydgvak3hBTRAtOqDk1oef9QeUXGEyf2df7s7EUl4PtpftXngEtpxi9omRB9pvG4xaFEmo2ac
X7ctfTPK7CNT1y16DL/yW+ZQmNESwlmepXsQ6PKQYTDzCcCruUlELQ6jJP/pGA2ymD63uoWpQwsA
dOa1wi7keev4eDA13DGmHUbsoUwcAbzNDVrsSER6+5326I67AbhrEQH9xslUyWJ+vrGxPit5zmXD
IZNGEH9P+oH7pHtw0LHXVlOHAR5WfiC09hu+Z/NRa5VAAe/FfzDPJ5LJnqpVdDHs15NJzW6HwoiF
Yl4k+5qAl3RQ49QJG5KydkNjb7GK3ANORRytacmZj1JLa8+mBTm7Y60ic6w/LS1S+bxXWPmHoFMT
xbK5DtPCX4fC3reVCBE6MZwnag1kjsdsHrQuaWTa6gQjNTY3Jd8ZOVjJNReVHx1l5NkgwhX/L1R9
bWVfb923tZE6NX6DYmRpwgX8Y3ga3ES624acpJ8bQm9qL1dG6AlE1tOpfu2MLC1H8OcIc6/hPauF
N/ZuSflev+TCRe9CUFKQt4JelL/qc4O1IfSRk2SIykXOKQjPpD4e2cc2ibrAWSROH3/PCExVEjib
K63yDaDVsfDIRL2jUzurNhc6wHvj36gQMApihIyRW4w7t/PlRa3l3wNWip/BXYVQtbfe1MumpviE
e0qwJ81oDHiuOEBJoEjXGrN9J0kv7YFYiIP9K8m0ATc0/XjPa4VuIjyI/NdfJDXdu2gRnitCZs70
pjq9lgPhiCTIIR845Ey3cO5wuI/+gqDaySkkNYoMy61Zi9cse3huOlXi6t4Q3T22EWvx25f9UkV3
BQJ7/RCOUufP3bsDRW11HUm3QSbgYVS5VpKKNzU9ARZ/ZqazbGBGSbE/G2V6f5zzxoDkDmvvvIgI
ounYrqwznYlU2c0pdcxxh4PeG+gSFhmx90J2Dje1xEztHdikZ+y4Uvlxbu17GfQWx9gyq5K4XZD5
Ew4+9KXnI3PbVrxhTjlg8Y/bbBxaWnUPpD/MIU/7Yd+l+kmzTHNKmKcVJrEBmjhV84que/0567Ax
1U3yb98xcirhgRyJSGljpSohN2+2cStG/FVP1ctQRv0kmPbCMaxbViFkd5gkPzN8tazPaSoQD0VT
vVYAI2KJPBYU7c0gsd4r4GtxH6sZvMy044pEedMjKY2+1ahKrhaf46DJYVYu9WrOBm/H/6L05wTt
t3ON9hKcIj1F96Qz3QLxnAqcae7+6kKj3JwGCkfNjwD1yvfqlmZOKWquxbfUL2woL5Cu5Om98lpW
EBE5/2+mgddW14oCuRNg9zBsDfU1fK0HBpKHXQDBN7XAh4ZxDc2V7cyBPqeKnH33tZoH3WhiK31Z
aKF7kUU0kqBGMBxmzRdFTggdLuxDiQPeSl8H7rpMD4JPVy95MBjpZ+oV1kwWP+jw2FP01eFG2sG7
eTFFS37TTRmYLBm354byvJ6nFxBlQgrgFgXtNTbCCh7xWLYHCrzM4nuQckgvFQMQv2nix7/fUdi3
pB1tOobFttaRwEk0cCuJKiWD7UQBP7otzQFEoWgQe9itP6JQgVl4yyGEkOWP2jcBpz7kqZmeFqO5
PHaZY7DfllcCdDuyYPmT8VPfLUPGXAgLlMItC6TSa+WOe1wGXmSTIgUMQ36PKd1PcMrIMMVUjeCL
+fApQwSCR98yiBVM8w3fQ/VE6WlgTvcs2swulpBguVOWR6CSUD7XZERY5uYUfmsU/NrNdBuDui4o
xPbLdFosUgWCIHgs5007ybMselvO/yi07PfXDTIC2r+4aDnahxRnmlBKBp+K6uAe1wX3Fg8ipxcK
2yKj0mgYwc90wD106gO+THe96WIqOCRZabDfU9LSFTItnTOLzcM6BUijBSS3LJln+zZt7arEkUEa
tqi/kZR8B4KYJyhW+tX/RWnqfChLJbMgdIyYwRWEhhE8DbOAWV01SBcMKKkGOEkxz0VhFS6ihNap
B/PTXBAFRDuuYEJtonAWrVI74dcleVGpa3UxsGFqmHhH0NGjkBH178WK4m1+JcNTa2y268oLAwYr
5v+7fG11KkUdfv3fjAaZkrFDGeSh50aB9FWwLRaukI0pAM751UrWjtjwKgpmxOaN1VBFVZh8wryo
CKNvR4hfAi0XEf4n8rALk4DxD2g4GRy3vuCx0oHjhahl+K4TgjoNXzckI729HxouyPXA8/4d0qlS
CpWCz4GS6uu4CwCxsFx5SLRjoXomVCvTki2KkFl+BdpOMiq7S9PMs4dxM5cDfzuvQi9+OVLs2ju9
0FHlU7G7dlTkXO8eX9IVfK7l/PFwgG59yuiMAMWWA7Zj57xGkVjKFJvA87QcORGOLxXzxeNkZ/v5
7YlCBKscVZ+nvOH9ohEQFAEJYzBXH5R2+aFMJgaBlH/JKVFQLtw8ONQ7/pf9+ViYeB15v8b6a10c
8u56ewh4kihctMkghPBWEve9YsFiz0OlosjjG3eL/kqg83DINL6m07gV7vh/7JFmLVQ5D0zbVVgl
21xRgmNqcGhsU4y1uKYgF7Sn21LIFBo1zykRSv+aH9bRav5a/2xhi++t6mkS+JeFBxce82+OXuBR
ljzqTFJDSfVaHff+k5oTiwyhi7Kb/w2DgOZiWRsaND2EXXjidd5+CPj3rFcsc6eUnX4aXS6rExn4
23utN6PaXR8yRNgNxI0sliLaYnNoHlrtBx8TbJo+0o5JNNs9QtvuSA4zaYCjKUjFyLBaz3qJvw4+
p8jV4Ljuzi9XWWH/83sSauYntEkmcErJxiX0EN47MSSZAM57IGrsoCh+tVOLnSs/nJx9GTU7nAkk
2fLWPxFtY58uwo4AiVHdca6Ik6SLvfsdJU+oLn2zO83C+3d5RLPW9cy31gLuI/+9F3I9/KbjxqMn
WoMxPA1gP8rLrRFjJOQufvHi+kimkAtgiEosHeoSCUnH6+VOCOrrGu+Pp9Ka1wvJszjAGZHe6ovV
U3CAH5XOmJCy+Hgbc8FS/kB1Up3HbsWKZQWlEc0ntnMogbvf+OM/tVF/C/92xMDvk1rDrPtJ4Mrv
7rmL3l5tdWlzVno5yHsgNzBZ3o3T2bdoW1NpnSDGEG3NDHa5MW5O2V8YeAFn3+zNMYJcYaCWCy65
XxJ23EgUUlXNOI6wD/bMLoMeyetPbLllMmsetxFsR3IdZh9vVdj/m0utbM/4xvuSS9WUaZ9LKSkV
Lf4iPUru07SxVxVY9PSVK9+U5BRvuFCHiv7fxUasDs2y/qfETz7sKJttF/GraW58Y7nT31YBNnYP
GoA6qH4G75wEG7bg4kGxMkiVhkdn3KCMEQ5MeGcAJArad2bS98k/NsuX9aC6L0R4m2ZdEGERknQ5
Uo1x2wzmoxx32khH9JNh7OUsNeaB5xhDmZsLIRcjpUZPnvBWPvgv96u4L+EsitwOX1hXJGIrZoxF
BeEOXmiNhCgjT35WQ0PDGtUwwMQ1aVBg8WeFNRmHRp2ARdT0yESxShk7hdhwoZMBplTH4nq9M//r
3MzC9TpSZL9H/Aq5XTyGele2VP4xckF6lK80L+2ipPh3yz0/ccdRQ8M06u37G6Ztv/oURGdmTDxy
CIz7BmgXBveV5wpGTuH634TyjPxax/Q9Mg4eBWXqktj83uKBgR7yOBxvSRKkNmFMAhbdweH+c5fq
Kw3SHbW1ETfrPaW88X9cBj+qrqY6jAT42jKeLWxYTH04UP0GHUiG8xffJ0EAxE7DGyIE88ld9FQ5
9uex2UuksxJZiOaxnQ9GPH8JcziUrVmCxpAiVPpWvgn48yivQTWLbO6AGz+9rluVr6sNKUvAZMfT
7vY1pFXWKnrJ82sJ0uTrcMpDR/o0I59Ca8e7km40JRvHNi4HR8hh6ja4rGworOjQ6LiOXxZ+F1vz
mFrnwdJYhsNLecUelzacuuIqjBVQrxnizC00d2UFyZh2oGJdB9421JE69zUkl+L4otGFM+Y79ZJp
ocOtnbElBryVXaTckrgi0QPepIBPXXAWDedsO5mh+53U5DAwi8BiU+XBOX34pbLQU12uuu2aafrG
c29ek95n3DoOxGDd7zKB46IyZwA3YtsBXX9A0BS6hFMziO7Swf+k7HC4KBsJ/I7uOm/bhGO/3Dgi
2BniKV5RQsVfoU7TkgYpXmQ7OGajS0v/xpOdiiK/4jDCECCO06+7IvpMAgdpsWVlw5p+H4f6X6m3
fXNpx5alGe8H5SXEQKOhsM6zamxNvTbqPjhMbvASfrhfWzW8WF8gWNPZMfg7fMtlIYf+DfO0IUJJ
61BPJ1Fz13eRmMG3DXR5ujAzrU4cKPk/6LTX0XmxOqNfbfliuRQI2GlfeD/Nf2urEkV5jsEKbCZK
PQrWIWR82rAFqYaTzRMXXEes+RQJ7/AqJswvhfgkcQi97yYvh8ltyOW4KMk0v15+qDq1D1+Z5HWn
Wt000CrZMOmoeUPPdum4QjCbY0qsPYRc38vRJ9SBtFbe58wUWJ73YL2l8/Sj1ghECuucC0d57fUr
7Azf10vv1CjCbqe3qepo0R847h5ScMZWtbOw5m6c87kGugJnhnvYtZ2KcaEod9EFkfu6s+IX00pX
03W+L1sfDyTyEtqFQ++DkeMyYYJa64zbSXF38UiJCacfuHuGLSC5j+Uaz3eIRoILB5SGfpQElvtt
4Xef9BLwmVLLstb2Rq1JfIvH28lwolJlxy3qlksWXoI9P8AVqcjJjor8jNIL4Uf5HRZrKmCOXGju
7bvqr5WGjftBEX01tkCF2ZNlz0aWdpz7O4QJTnr1KnY8tC4NEgFmqpaDGqU+ObMQ804XgJR7IQgR
4q4ZCLJbYHQkTbTWVmPxq4Zr0YqR0aRYa9nGErycjiNvwGp4XIrImvkpuDKSJba9cWcL2L+rKHtu
n5u0V49gdHm7czFvhJM2zTWvzBHh+uPrSH6znApKOqi3IFRLBaZaPt6zqyfrF4H7hAMdtrXifgoZ
PCFORBm1jHfb420OUMUDT5e91eIg8g5nLqKIFteU21jGvODGkAh6Vzq4jrwOBdgrXT1P5Pp57nPI
u9MJHHHarmcVXFkkLUYs5loahRdup1GgG0uzdHB9oE7hYq+ucSX0EYLmMG5j5v2gXbiH33QJs3Xb
uMZqkM+HkmbpcRcn0dKEM2uRNxtuXhxyc9GeucATaDUspvbqPptA44lTdSUP3+mWVz2Kk1hpTeV/
yubBtRKa5xFfG61uQtPCoCwREwmOJF8gTp8q0JlvpwMQu+qYWTsfzOm9SsOSfHDbwjbj7IxRZozT
5yZzfrHAURBcSDDMo53t0j9a5qVrRmzQM/K0EwaLMNpyWMu1S2UmoM40RbZXi+duYawtNVf+Fb6L
12ZwnJo8lDbvJn00BgJgCOlkLWchEBczqM6YLKtO3uvmHeC+GKeCUaJcPqjA4X7D5//zi4LWMIJf
0NWHteR8kTsOe7OTHhZxnp6jaeK/mWHd9dpGJCiItWjM09BE+hLaHwcmqPESsbo1ABwgOiKSkhBd
N6EdvoQmB8G9Kq8zWs7DjAjlaD4ZJXpgZhKv7u3/BYBAUG7ACE65w6XKy4jxtjs8y7OytkkbgF6d
0BCzZ7acjJaP4WJxDBe9T1EyR7eMsUJkusZKucm6wAH0QIQEnsMvOIk8/zpGrfISjAxvYxQE31JA
h8tR3EfmmzFKbFtDvLuewN5QkAqseSPhHKoK59Z1+q46JNrgaab9FRLIvNcGwxjxW4BCHs9GdPdI
nd3ms1UrCp5i7PaF5E/fYthXrwQLSU7UxShhxxXzfbjuuC9QoalaVH0rJtTG9LKgeK238NJsZsYq
BhZ/oPadgo4fL0oIT5oZB+pl/3X4F4vha1k957ds6W9MLoms9CEboNg+1vuDbgk0ZqjHsGoJ56wG
EjBC+Ag6kUTiW3jjf3DCZQ1WSzA6iK5h+icFUfk+2V4fQB8zmc9llhawngmhv3LllNoJZB7Y4WHL
2AOlhnfzt25S9lHcKN2pVQONzpzDbCGn0XwELRo5Lpm9Do0BGc+QRGgi3G+GojSHgtCAXRgSCarv
CvfylEIi8Tiw2Y1Ga8sWlnN7EZPK6gmvTFTOEMEZnSKrIj2XMUcCQhV5rC+KK6ydpHAh26SacVt+
teQSxWS5xx+V7QZZuLmlbs78akrcslLImkCmasY908kE6q5u3kmgxGhFeCkC2CSa+qasqog8nb68
G/FDf6I+dOKVQEvXudwMGz1GzIyc7QtkhxTqiWirZe7ZR3Pjss1M+CFLlFWzGHtxIcRzTiX73ri6
s1+5P1sM6Yv1Pj4ZnV0dFnd2ehce8YdKkRgq/NwFGb26ANDVveSwR6sQkhJUhsDQVuQ7BLPGcMgh
EzcqmFBHQiilw5UFBs03buPVnx5bz9pSZcIjuKueGJuz84nERuaEVD7esdtCkSdhn9M3JpJ0W/hj
MmbiQ543Gt/cnvX3t35YxKV8+ZIHx7d4DFzFuwtxAh0T7rym0NXfOz8l29236JDK0jQnzpRswyht
MR4w6iKnNcffht93gwP4cFw0RtPXgsdU1B3wnJvlRpeP12CiLTTYBbOcrCdknsqIAdKznDcWduCy
nUb2rpUhtLHjD+/grWIFHCjc1zObVklu08h2Qz72U3Uq6VXSoQ9yPZ5IDBNaiSuqQUkXYXd8bPTq
uyjLc1hh96I9XTddsg2HruAZG8u8cvxqtKrGbwrkVR2N1T5++ouEyH9e4xG9Tpr910hYuN7yr/e0
PwtED0SEPRky4LDn+H8pc4XNGWG9PM/LFm3Nma316nfJ7fTaJIfyN3ofByMuGBymoVrBBIXg1LTS
FeeuEnxzsWd/eFv3n/TQY1IDOQKNpMCGdNVwHflgIwQKUz98HOohTxicLX0etEGB43TgdWlVNerj
y4o2LgUdQcS/C/827PobeajVfQefnleNW1CibV+4LlaYIaFwBXbjfz2BkB/NobzIfEF2KbEmDyXO
8eRm9pQEqeWx2odNOM0xGOtt8RjPw4gck38QKBoiHnhuSVScoo8m3DX4LSWXkzG14LjmqeHg+Bfu
ZhqN8mwYHXDr4LvG5Rww9p3/RNhTIxSSsOC18XYByem7vp7wK84lDvMVeCICt6C8T9u6Mfms4ayz
adIefwzxa8jDGSXhfRWJDQF2ZIUx/5si2gMidNU5S6YUqPPtl8V3LoIXwM7ZhxaX6S/NvE9r/5JE
oOWiUyzRybBbxxK6U+FCoRFOm30DpU7ZX2LydN3oal7uf9Mea2tjRIG/+HpTLF176eBHDSgnmVTm
oDLHuYjiByeSxVsyYSJ9G2MKSDmweBCv+mWjQWNfaFloeNOX3FfColHuSqRk5AQfg7ylWdZytsgn
cYufoM0Vy2CchKwmTDc6ljEGmo/AWeRXQ+r+BK/bk7kaoqbvBvQlPIaBQlVbvpEu0ogCns/GvRn+
70bu1s4zAmRv8m3ZKjgygvpiwqlN7mFRwZGo0Vn7hWqjQQo5ZQX/6CIZ2zDTXvuRQ0n1cPge60rp
pYuU4fQN0WKKssFnEhCZxZO9/ESp65DdH8trAnRiooSg02iojIhLMiaFekoN0hG2WnA3kBi/QhhD
PIpnEfERYt7nlYYj3STvJbMQfWSc9wfO6+GR0UQljWc6ahgAJgSzDNSK7domi9P730oEx4ZXvl1F
XBbCdbkKgyCPTETm0/9ZmJgosO2UWL4IcYaIyx8h3fBK400RirwGPk96+C3NVS+/X/A5YrWZ52mh
NKwSPkGkHoCAHMhXuG1ML8nBYUfmUDIzUq1htglPwcxitGLfUokT5OGPfWeN0tkifyMwJHQvUBbo
01Wud87MV/5wCMlaLDE+mkw070fkA7/sKh+C5/1TJquNIN659HvLJ3SzuNgWZaL9k/cjWvvgfGXk
LWwCN2K6Gt7D1C7xEQ282wrT8W7E6En6ScWNwuHz4W2cR3fFWdvHVsvYxbiWg7SIL5otHQC3zIqT
NwwcvlarFAWnShnesnVCut3oG3Q2t5b9fUXG+ioFckV5RXOzGht/IHzm0mKguwsJAK+hFN6iWUy4
kzq/5Q0jKNOCaShEyo3AvltaDL7pEb4kIjUQzNYzvuTg7qNTTMwZ2hi8aGaELDGJjMnrJXgtJZZd
aoS8XoqCeZdv04e8AR/6TzUuaybIcod9Dyk9m2avduuF3DL/IsyDwIs7NHppyVNiOawHURnt7pKR
OOIsiCt5qf2J84v2Ao1LSqhR2iYRDng2JjnivKv/Lsq6qQ/awUsbFtlN25+UOa2din+FYxjrV0H1
cyQ0o7YXHoPxlgfU7efr0DQkJABlMB1ep1F4keILsNUqpiwqclYyEOHlac4Rl01Q4eCPDNUzqRgl
ku7ZMyRwDWzuDAWUNTOomHAui15wPUPf896s39Y3vMRYKBjL4FIwxj5BROOmlc9QLn4SkJ6HMdw4
WmiKcNUzyQqMm8k2XHwYKgo261A+TslpTnsU960si7hhCX/6iRKhHTQLFh/grgj+u0IaYpwbUvrB
/WX6oBMc6/WqLafaB+HGZUPpjrM+QIkqvQMIsyXLr8PTsulhWvQfgfS1Zq98UkW1GoL62zkQIuhx
gGSxk70DmGtB0RwxCjL2FPjZn/z5LrLU5H/Zn7RGq2NYD/lRbsCETJzChVCNKGVS788RzpvuLLo3
LnYQBk+T46B2n494L5pxvknkg80RakX2yY2GjxNVU2eev+bPv3VclGkjvpalxa1kFhM7OloCd8mO
s+0OchLsK+yo5C1Y9Q+VmVsAwMheLTKAfR9pFlrCrvipU435DUlMOxVn8K3H7fAWQCwFyQG5WTYa
4OQrd2Lm9SgBZ/RH4M/U24+0uVtNh2pgYdCcE66cBrnpjhzgKCXDsgHSIXbtiAG0JTNErnhS+IXd
TiR+jH7Vp1NL4wUowPC2LAtlDyhliNgIgIMkRwn6Vq+E8Uoc4GjbS0wXUBt4XGVH9YbfQXh8sto3
sF9lyoLIfiCCye1e8KjlpznuElo3Kw2swoavfKcdcMp4j1oOWAK1Z+XgVSVbrxLY0h9MZUwmPZ5U
ql7Ckp62cZkA/v8L570hX5TEixPOCh4+Yi5Mg0JNXpKlBZXKEMtOFKHRbPzklJLiQ4n5zzpECdG6
qlLNqZmbEv/D0ExiyDW3N2ZNeWe5+nXMYhc3fjGc0iKXa0hncj5/mkm0SkVJMpQg1D5TP513Srbo
3KB8KH9Q/E90e9gyar2T2HDl72eXSFCvx1ECTjP17ZLkJB1TPFrvptCYxPVd8+6GDshoxzbAVrJ+
a3LZCPCJEV3xdAIDl0W9LtctWwaUgiBRANQnyqhqZWy/6AbTG5I114BClUKnJKaP/OWg+SpY7M6t
/PiBdzdPGgmpfJ80M34Xa5cYdP+FGUzFahOss9jt6t6JKNvFkE2u5mP/RcnwYIGNOxpCrHoTeg14
RZgxh6RTWxfIHFlcusNd4wAUXP+OQuCK2Htsxn/7GdzeBsAdN8wgBUmHwMRO8PcWsivG6yMP/P4W
jmDC/8U/I1GWLrDB8Bg+9MajE05qjiHDOkRLn53FUswf7vQ4lyJhPO3Lkc4jMtvQXnbfUVnFwsa1
5YatL5bRbWpTLU1EmZXAAt8qp2AvQ8TAOZYOUdaJDmahxPdh4aPbRxBdpu6cOHWjInqPzp2a14t+
KsMZb6NNhsFzQT2AtZpCvDAmhX40NU3pXF3NjvnDuUYt68CU68100TgrAIJ7oQ20lYtklnx88lUH
0bkB/5thav3lUPOj9qcFKy+CtDJfHuLBvCR/YjiDU17n1j0Xq8/673W6VonZH0V0gWYhc0+A0iWU
jCZWQ7EznOJlM2HYTcjW3xUQ2E/iX2HOJrmNJyvKSxfhrmKSqty0GvYl/q9AXh/AnL1lXG5A9aq+
8SG9CuraObYd7SGhDS7mhTwcfKORam/0TkfYz9Gna1A8AiaAFHl/sBjx1tE8XJelWrOt8TNPu2SW
f5YaX40pFC2mQC7cK0EhjvGvj2TYYLuHRfmseG+pCHdARPXoo9hHMKoDM6UFCjzHv5fmr8PGv+yS
7MopsidC6AUu4dI3S2JtesEz1ZAZ4QaV6vP7S07uUNlsSQTRZxbuwlqHD/7WZ1FIibPzlJa2rZNI
LNvB5pgztE7zpZCU7H9HuYUR+MS7OVotv1dKXrbibXFGGaPgBjf49tduQS8tlKj+kadYjLGsZz0w
uj6iedq5VIfgHGSCVbtiHU4CZqJTqPvbTjQCCJYXrinCGK35zLTlJ7xe9VVCF6wzd0M6voNt8A65
58KRbGU5La3s3itglIIuDWy5tF5He5sw923nrCjoTFp7Zyek585Zy3cGKiTiAQw95E8Xnq2vs8cu
qkpTDlGArIuVqNa9XFKivkc2+r/xtUDwuVQmEDDlNP/RKYQjc/Vz0w9Zk8dpaDnnYJovG47e6E8b
RHLdRsQD4phgS8YaZbsamho08saW6vl6SYkiunXVJY9vPy5pOx8Y/4mOtcrCmYk0SyP4vrBZi67F
ddKI6niujgf9OLnHfB0syzE76MJEMRfA7aFSBhR7ioyTDE3CGlS88EXTD0eIz609p5UYBcKhnOfK
LZlw2L3zSZGG7tvbKGdT8x7qL44T54tXhlqn3cGFZmErq7K2h1h09lfQeqsVJNUgPLQRr54vOynS
a/an3uBt+7FnQUoyUBHgknOHb9kKk9TK69urIsXoof112EelmzE9tbekjcSudSI2K1l2uSMkp8JA
2ROgqFfVGsqJy06Q1ECGEu47Lq1J6F7u9cH+sdfzZbrVm9MGtiRpGTD9/m69tIMwZmTPZhLouhhJ
WF8sIRLWhjxw07A1V8FrG3+eU7GII1Np0YHdQLddCK6wLOqQ8ULmK+TXusTQ32hrVDPbGUtHbkl1
IXRe+t8L9SUTEOk2ivC45Q16JPfsfZqGYoc/qJ5mZ5DrrDuZMAAFyJ9hJD+FGLd/Y9+SqkJXmZQE
4P6s2H04s43ThNgaGQi3BOyPUoRsEyiaCE+Yk7q88M5Df6nm67RGFW8j+JoYYrZTTOH3/CkPRRGv
qJ0ANq86e0H/+/XRUrBsIK0PFnOgDTIqBM6rNQLDn+qI/Mvp/scguq2YpXhi6RfbGoN5NnyKaKtA
plTjRUWyM7t/4YYyuhLdwT3IMKR4oOhcH8TknXyBQZhbmO/amj5K88zK1rUaB6lTFoZIYIItRP9W
gf+ZuwgioJ8eFv5nowRbsqq70435hbSqPeIUeddpqKG5Vjt0GUrLmh1CO7yV21nepdhbSYjYRdeX
c53LoaeU9QBDVaMfLcUPH/maNxQIo7uMWTBsrItPaF1GC4u8DpKXr1NSbm1iReF8kTWenWaI+WUq
WAzp99p8CdreLol6shCR+6jv5EARouRMtrArW64RusBnGL3BCR+0mawDAKoMxRY9NPtk9Vwob96m
RqjB5/utadM3V8K70LdsAXHZuHlwL7nr9434IJuyNeBwueIDyvXXOqCheEhKFHK3kgS+dlDfrs5p
aRzc1w9w2tFAXuBp7o9eatY9pzhHEh6L5wZVDlgzsR0nB/XDz/KdyjTQlfTmof6Ip2n5toCBQSPo
rdRQD3vSZpUtSoltlZwDyvvehPVzWSXovMSuzVuzD0L3mlEGXsue1SB12ssSdycMUcn6cxhvGvYp
8YKQA7CxBEUFT8evaBON5VaXSijtvHfJuif9v4uqaQ7auJfBaA2N/ZRjUUaRyV6wDVOT7wFUupXY
ekgiGQ9yhDGgW4DTGbnyyedtq/JlExiH3e7QE4vBlOzj/hYaap+70JBVxbmqO4VZpqigHMnXQIQq
4viMHCSDvywoE0BbwsNf4onvZehmG0wPnSAjziVbkRvdHprr0BykCsefJyvwzxmmX3gcGplZWntZ
iD3Qx1QqkC/SoW8k/tSUvc4xhUA+mMU+digHC6AcRLowDTJoNgcSAvhyRaLQk0Xi62T2TZS8OS9f
WHDSQnNp2kHYWwrsVcsje7mJ4kkBBC3f1+A6Dm5AXwSggq8ilAWRjnhQAn+Ri5/u/2yiR8XdhwBJ
L3HoybNF+ihSGoq50yOAYEQroo7dSo64mmkRCYL70ayEkigcS+uT0dzLTcgASNpLv+DtBm7qxzSf
KMZkRcu+rnud/k7toY0cQwOhMWb+QLbiJ7cm52hM34AIlc4uoafVkuAJ6fFKISLdKcagG4RoTTx+
yHu+ooq2JwP+JQb6hIfp0PgJ32Gj38Pisjr/ztb6vHndRFmbEGoTNUaB1dTQYKqxxUCNIFi7SxMT
hmLQcD9TdfCXAYlPnmegvqN7HSOphuTDcIQyIYTB+iIh4D166ZS/PiQswDXZmelW5zZa2E3dMghJ
PF/ve7lNEzEBdyFv9hWop2SB6ULnwLF9rNc39A3/RH6TXI6ZWxLvY3ECWh1kS0viyH4p7PFv6pet
NxoxlGw9wyZrSyn309QVLgylXULK7zst2gOd33TOnJhyPChtGqII445sz6dH//68bMtC88oC5w32
HKRiDMyzTDPN9kQwanmCxl1WC4lxL6uCs8gXsM3CMNrKZlSKn5Imm3aIuY+v/NWuNLYye++1ZCdB
sENiBfbgsJlUmtFiq7FvryxWGd9Y3rKZodRhuppn0BMWiYkFjKSLj2wAL3Nll6si3hcyFQbWCgDT
gyBVcGBlVzIaFOur3R/+dQEa5Ep/acJOXmDEc0YCy3ChMeqRNulwc+16JF1UpYO05R6hanYWSX/5
glS1/ZpL6Y7DmHh/5DjjZqptB5kQtN9sNzuHPP1SklF6ify7EneXOC4zbdR2CqH9Qj7lMJVVEpEg
JVDne8hFbLXjPgA9xP/4K5wfDrcuvfAT7MnHlBzXK1gAbncx/Xmq8P19KAFbiL7gIEMraygsBH5E
ElnHGTv6PHe/usXeLxpaUkXnIJUseE8e+Hy+//hw2fESDOOGUM7+1d+aU5TdahwtGJ+ATfU8lWCA
3+QgGi58y6JXDZPKc8LiX/FmJxB6e+lDF4B5sERp6wa6nRHRRKWx9UZuNqNC1RUqRnFSF7jvNyGN
vDYOBWtXBlQ2y0GESUhCzX/0cBYzw6loXaaf6ezsesUmLO4wZHYA1GJz/I6Ah7jjbaO8Kfs+6fBN
Q/b+PAl2dtpyOOCyim+KZ757DdCZfN0JAYIEZ3u2+KczdrbqUbwt3J4WAIZJfoW6Q04FhchwaZ3b
z2icIWsQYtykqW4POwX0nRth8NEfu2anVYLnc4dqFgPgEqVixT7HrkgLPOSbi8VDb/Q6RCqtw3Bq
ZBboZxl161rehKRyluzTfrr9E48PwB2lOsuUozFXJXIrKdOtk5PiKWHUC66R+phHDjEvGfzNVlEx
2TeWfQPJqWY3yKuMOLAlqMruq57kacr/NlIUhxynaXk2dtjSH+iA90MnB/rOXNe1UJAXBf1fi9Yu
hsXAtbbNjy8kPruzaKOhXrzsqE3iOhUqca558lfOqWqr3cDJqUz1kzgjlQgJFwDitJtwKSzM/Bqw
HLBk6jJU20H93FTXPwGilld8/ZGX7Zs0r+wnej7mHo7kVfIL4Dh04499wBW5I/0IHiUHX0RxQue6
TrpTcJWhs1Elhalf4UfK51/D+klGlkKwRvbzhsoNXqLlu1B0KIN83XVOJ4ikYyaMqHxhtA4u4LFo
X7TmaGqoGNdOFLeumqrnBe8Fit5aYAYNjaAwDBkWssuqq7ZxPuGWXL3boWO/rFMoWK0DRNcfubrC
fwyrLE/uPi0QAg2kUBYtR+K63C06P0CG92eDDGi1nxho2pidiGOxSmWv/5iCW9dQZQnkcKvMELHT
EKKVrVuN889zx76Q5iXRSj2ri2myOuDidFJyaEBP6t94h7fPTTL5IkSsaGy9cJH0tXiNBnM72AS9
VGmf31wKGsbrFD5ApM736h5wjn3sfQZ0QEFjiDN8wTj2owS/IhUaMWIEJRhiTs9mFjpQf8sSotVA
YwSWYmKsT2Syw5k+zLcQIOOInRskDgk/+A1OI/sSwIFufTmEq/8RALz1x7WpuW9hrxwNQjbyiU0I
YfE6gxlofNihHWVOt1RwRp0Z1VRS7LuZSzXpOlEmYr1gyyvfX95hqzY9QORmaG3HbQ2FLchx/wx6
IkYtL3vW7+UMsiQRoQIjQ9ZsnnJEagDEz5tycvqaCFBNoknTWDssXD6YHtRRH74q8qvi3M/RZ5Zx
mZnvxV7Tg/cLkuQlin19wbqj5TgYDVj/LtfO4swD0vEkqVP0e2sG22G0+545G5Qmus/4GI8IRi8C
YzEqqedy9Pq8zctWWQbn1sULS9wps1GFFx8745Ej5RrsnD5Me7PbkpW4avIDlyUQBvmIr6BO69j5
LQ1Uc7NdhW/1InALvMMAJxxCty+Ah/zmZUJ0wSKLroKnZxcGld0+ZLeUH4ZzPOzCZpSSAsN4pyqJ
6l7tjZBYBxNjo9tSCwWvgfpYkJJ7hKKxflgBRun4knFDC7QIwprAxzYvuXEOSbqE5/JJRQm+XzcF
RD9WEd888S7K/cc7YHDb4Pbe1OAa/T46C465+ZNsoGjPTkI+DcAUiboZAc7j46nKYFMUFbkJXz5c
SJ5Ye4GWKvGT5XYc3hyVTSkv0p5o6mub7yYD4aNofNKN0tHxkl6AuivSnodmTLD8IZvvBER40DWS
hfoIp+z0DjLViZfJFIMpZKRtBw/71HSb45xks/jAnztHsKBsJEhNCZpyWkzMR/BN37k0vMrK5VUG
opX0xsCGfJR6CMsXThkmtQDcM5+66Ps1iSkUF+MU5/Kj06HnBV7Hsn35LbOwhkN6W7ODRHdkICk6
FR30dN/FHbFxleVQxS/SgBZ6dA/FjZDvcwGtxq20pF9hWfGnAjbJ9YdIGKNYnKpR6GeLnjxqLkHH
NKgtyyptAPeUEIYJ/xyPtwKG4sEEFIYXetbFWtxq64G9XRjbEk/LW0NglRjkTlgnBjzTMhOkXDxK
sI02Jpke5W4AfiQbtFRHtMIXWAvw8WMSu/0+ZmNsSOpizvJ+V0u4sBIPvEUIxSksRvNlHhICvUdl
vDo6EzP8i7OTTtLcJCR9xTEg9z1lNt2euaVdEZ9k6G/+CrDFze5DiNRHg6BLF9Tbt1DYpCFgo1d2
8BDxSbjhtG5DHUKKySfg6N/Oa0TC7IcaxyxwHOu1OW59YI7kxCDfC8cm8ZrbhsNU44OjHNJqaUx0
LINUODOSMyYPFAvn2Ic00Zj8GE6bTvsyvT5zmsUr56tOfc2c4o0o/pHmCpTjxTs9WxYMA73f5iNA
baeC93T8NifgQAMVahPTN/tZCuNnT/DMcnz47GeYeRYTzGP11ltgBGMLQ82+EMPI9hMK7e6v9QuV
PdgUcpAEGhcaAEMuZDATJ/Jwis0/aJDCvlKylDKt05fshYJx38zbLNrdTF9DVAtL7Fs/R0wnPdyV
DM/Vrp4keJPr1dZUXoeYcIoRZPScHoiCwxC6gWxIQeJqn/DUp/+s47tkYcqoUSDJyFxYqD2KSsRg
ZpML1ad1vNCJM4OaB5M5ezRWjfjKvxZLyHTMQHLNPBEIjTuIZRg7qwdbGwNVDEjt3K6QZMmYciJs
576c6UJ9QTIH6jRmsIZ+n3qTk/DqZANNTamgyIceC8gppEXQQCNlPTcdY7/n8hFVoo+XLJNtLK14
N4XsnsI6t0EfZ8dUrj2gqnLvPaLck+79msOVje3bobf+22aIl4AYwU6OiIaYhhULCE4YRnD5x1nL
v86Mowf9O93MUpZ3pqszlyQtQkUPWb/iQD698C72QsjwL69m3fIlERdwbKNZwg8e1fNS0SOfmHQk
EWXoCxcyarLi82woJpXgR4kSGswkxgzTH5ytt8FAS7QDWZAy1kR5E1e4H7Qe0FWZDoBiVBVT8NU2
S3kbkefZhijxQeSOYRZcdOCQURW7ROwFlOtZnuv94oRRR5PJKRKqi4+3nHdkJwY+2jPmO31+xByl
H7ou3Qv+uye6Msp2GmDeV4fJPMBxVN4G2i58tNY02VPXJTbVw0vanY+n9xcUBy4o/QS+goX45wPe
aJ04XMz3guzlGNzklvC01VjV0PSn+ZdTQp+8BOX/nhIScpjj9/ymHqPsoK7DLmOWj17ClK8o5k0S
PyM5f/7KKHcpVNgHshcAs+1IneeiO8ue1P3+umbLudH1vt9TPoYlvcBIpOQ+Ac2PHT6qadkjqKm+
rKH4ObpNDSjf2g0pqqtL5YiDuPvkMVZSCAFd5arw3AOoRp4eYgKP80EqmGGyM53l4iBZ1lod69Tr
J5YWNlRHK0mHh8DSs8IEnAWMGB2w/z4tlAFiiKnJb1wE5llT/+1VNCWX2GhmrzwZycSDT1IYwAzt
HnY78f7OIo5FUWV1vDdRmd/7/ZwFNvCys3HHC+fywILzBqMWI4pnlpy++ke1XSY/hU5rXCr7LQ1U
1qmJEcDMlQ1XJNCENqypM2Y/fM5x7GI9Ar/sOcifroJOG4IuSNT2X/OYrYMQXniiKDNxrhCGFcpA
2x42zDMZLe/uO2bsRhQxYSjkCnhEpXZfSzMH5WxmnzJy44xwRJhFQo1mQBewHW2XKIROSfDj5+VN
V4S93EesJYm9orUgGmUrSRYmMA4yQe9UC0gqgBdJEQ4jZ5lPbZv/Bp4CJP5/EFYrNVekl3G3FvYE
6Vro1gtNdmwhD82uaKPKX67ajtBE9zpfuD/1bd4n8Jl672HaJmvR/YYedOH+w8L4cNFvg/86SwzY
MKZDy4ifvYNzxALqUOYMy0xJByczeP01olNoyv+nkc/OvIkJ7xxjz13VxxY98CU38SwDJKEJih6V
j0SgouhsjZeDKnOxnMa01M9RI+1umkIEfWMh67V9kW8Q5OZ2HzB/yfO2vdERvKh1eDnS0Gn/QMnv
9eFJDa9JXeN79PsxwaK+wb/a0sGva2OutDMw3aM1gUZ3uukbMvl77G6gRBi4vcW8V4f2gzjL9Kx5
ReNtU2NCJ0FyGa6SlhJQQjr6LtTqE52m0CetEZ2IyUNPSGNKTc1vazJrYXmCzKZDQTgAwnrk7hF6
69cFXwMpF38uSGX4+DU9akt66f/TdwJ/ozNvWVc/Laq20t2xS8GELhTXZ7ztNn2ddqJBFRH/8Qws
U02UGe4Q2IU5WifuyF70RBW/AO8tVOepG/NSykXemFtwBat2urX8DXNx8t9dZP6SnjVF4dVSO7JV
U/uFcN6ADy2ai0XT1YMDcLJJMG0Rlrowfi2hfuVqDLjufDgBEg8EVJLpD9CrJ9DlY31pUbJ0Q28e
f3vJQ6YDliONopZlo7gYDx78hFQTd/zoWkB+mZUERIbdfxSjL76Dl9jjtAcLkyMHlIDg1IIYEY+r
dqm5Jqj8RQ9bYi6b3PGzK1/VDMzvibw8O63VJLW+xHJAvZ4Qr8hn5JELvq9KUwxmeNI3wyNcFGr8
hb2B6gZgwx3M31lHzboHicAwiRNYlmFVyErN1SJyov9OFZ5kVMFkm3qrQqujo8cqxYcl670J04gm
w+5UjB4785U5/4y+XxGBc2c/EsNy5jrAeqH9cjoaVFnJj2YBoHMcdxsPrE7+DmsIPrsOMUUm3VMu
d2VQ6yVbh1G2s3D1TXaIZnQDgPDiJW7hGUxERlVYwC0l+AHamJfMawZfJDM39KAcsZdwgXxx79uX
kfPr8I2r5gWHu66YhRGiBO9cysBvcV0rObS3lfZnoxqSivIfAS/Y+SlhGOpDyOB10sujg5oP1kql
8q+Eh3cHnTgU/D5G4gyx+xADnCH7pYUTbu3bdPogqkZWYJSRQIwfzrvWNNZSfDmZsiN/Wf934nDi
hCgmveKvDcgdHCDw/KJJkr1XTksqz9HhqzuU8Jvjjko9eoeB89xqNC0/nU0UWXsLyuaxAvBFD+wo
0t5Q1CI05/8vrJkFDLET24/tBpX1QaR3lv9uYvmVDK4exYJ8TyI8CLjMBmgK0h25muXZOS20Dowr
d3DR0Zq+Uq/ImthiBWkBfLhj4FpL12cUmQV7tjt2YrgVeiyrtmjbe1xk31rTdDT+UoiVx3iw1Spa
rJ5f33c6dcr108nW6cRHUE7lC/Wn5vOsyBIZXmPnAwB0Z45dYpbHLnwjoXXiEU/EuwLqKkb7c0sx
DbG1wbDkVQq7GlPJ0Nyozp8U6fBNrTSiQchK5z1hz7GpiEFGgnipGERqAEQEjS8gVUpfx4AJTs//
lpB6I9QVqoksOkh+H5RBi+XMrqzceOTbAJeYmvfLOZqptEd9Zix7t7cuqKiM5vLEvK93E9WydMBz
wxhkmj90jEShbMWBTgJNn7ioBnLCOJR8BNlFd5mt4KH4IDpXPcCMUSBuKbzx5sIcvJBhRrPlMgoV
rKm5sfw8mZP4/Q8NliSXAxKhzvQ/fub3CCdOY2D7p+c4mt8zI/r0MCuxRXvJ9iWdBVe6BbIYICxT
ZulqSeYg9fQq/tNGzrUvUel6ylbFHo5tmy71KK+KosKYQRRk4UaAzZrSGjy7on//UTQe7+Y5+Q3I
g+132vrCnkN8uztW5JmCB1Z6uIKL5jcz/HsiPTH9dDtD1jz+1b9qyyzjRV8CStMBEVb5rmrC+5Ni
exq5euYnYKwv3smqjev44f97ph4gVZ6wyq5JCyOICLpiIZbPujrSVzrMdW8pY6MY1m7L4rWiEO9T
63EzSH+eEZFEwibtaonNtpDnnL18kuiw5Gzpjkhg1z98PdgRUumyMe2ejzVHvBpi+FKM+6t9Nsrv
W4KvXqA2nt+dcu/IoUk9kBKU0TcI2CW188O4mm5XeZSRXmTepMK7vwh+bhbwI4YuiCMLKltmQkVv
rW7xVqAQoBSmJsiDnibc2MsTj9K03cFzH35BMOM9RipXL09jWAlkvp6MwdZmabH/p5Xtjnyq0rJq
M/qjW1+YN5xaXM33pB20H1TQdizjZg7GgX+81iA/vsj3VeY7s+17bNg9lUdHB376+z83bPPaDVkU
VpiqbhnogtLCxu26XAtHChy1so1qIEEONnJoo2VSEtExmh4a0DNMffBb/0fi18N6HEpOMw/FU1dr
bZozfDj0+YDGFx6GTC0u9pZFwY7kiCI7vG6ZBN95xOju6RUDFg0qGKbbbYakl7JJNYlE0EhJAPc4
9F0cqt/Lk0X1iDXQxpY5hRF5jKxgxVQUlPxyfej28s0ldiQeuU5KFfOQNd7uCLHObUXd0bWFRYrl
J7QBU7XQMFbtb2SLlPC5X7dCv18CLTv/X9oacgqKIw+deFWz4djSIbFe0KBm/0MYGFnTnTqfy+/J
AZKQwvVyJp/OgYyfkJSBxR6JdT5iWmIu+CdyimuqLujXXZSKFv+QHkMu5CfaQVDzQnDo9HVCBKas
Wti1/gNIPZAeihgiPHvRhwYinSMOvo16LSYC+ygg/FaFu3UC1PoQ5i8of0zAWZ11Y8DvnPWreg20
EyPw8sBNNTUWGMhK44JK6ahw4DnByXT8u9kXYy1iQVvkRxdYLfCTPo57CjFLmi1GFA+Pr1Ct5bUb
owg99+iS1L+QYHs3Wm7gmxEOgL99jeP4/uIE7dpilpEQnYPtxnmYzj9B7bzvW4U+s3292ZZNBl7P
LadYdFnUzPemi4jUBNUbKHOQdXk8XNFvp8ot28nlQqm0ThBb/uyPseR/qAjISSSRJrfzlZXg0DMS
SosUEy65sQx5dc5KEH9zEQXBO6cnOvyn1yKx5ff+ZK0Uhb75ceaHWx4MAPH+l04Y/ErbPmwsPxFq
CabsDEgXE4QiIqM3cexfy7d4Ji3sHRBFUQ3kfZf2KTJrombQRIcB7yzYGfxwkqbRnQ8fmfL6evOM
3g6Dr6B6Z2RKEpaUQuvov8b6fatVWtldJqCgQabKgJnS4ZthPZDII3LBZwVpqMt+gReK9ADEq3NU
Eoky+oJlbxKQ2wC3YMnYOpKR4GXAruUCppsgkfqcfA2vCbMTUjpugVDjaS2qw5QrGeNczZ2DNPmr
1qdJlCpSOQoS9e2LyG/0cZgB8JmVobT3364TH9Dmv+yMhcu2ISRxDy2ZlIUAUBAm+lWgVLqhgPEc
X7I9fDlOwLS5iYHYxBNtPRZQl17JPppPIxutabHkwvUhgTwlSnt6cT4qzhb3dRV/esbtYi9cP9lG
GyAkTCzkpfLCAc8zKif74z7Y4NPuwga4oTeFMhkmdA5obNryOXHqr9qbDTGbOyd5sYFR4kGQoCgg
h9b8eG3sG1t20uj+2tK6PaAXEpzELE9iaCjb2YYk/EL0F6v57wOmT5Oe7k3T25n0fELw5UtmGh6J
W1c+aqjgdh5ISEG9OWplyNvZjhzB554Yfg2UkCgdBA8I9o6RR/9vTtgPcFfOQSBgAZrdPZQo9gnt
0MTnol5TeBHOTTB8m+pTVDluVKNcG1d87P+ORyuwPZ+LhHmsgItHg9tgh6uPrP43XixyMaEjM/F0
wNI8PU2ki7L3uiUbADkWLjgyI9RG/QVGiSNKiYznexFt9MTjILGwXPEffxoSz7DOA4YzSalCd2qU
qXa/9ylFI0z8BpeiJ1WaEOGVgRMY1/sh9jQSOLuxgJTRy8gW/qbE7ng95/TLeSSzn/VtGylvD4rv
9jy/Jc701TIKV1GVPMoXK4Vh/TarWUwXP8y7HA25oS/cUD4eCnFKv21y8pzUbhk0NgYqkggx04t3
nvUN8tcjArLiwn65Ge1BUcNNcUaRndov7akC9BuARrDeyTyPWZR8hEU2IdTSvlM7ObQLa3BPnAPD
406xUyKPfkxoOJtTfKteEbsLrO0+0zltvq1OYc6S9DPs7/kPW+QcOGmsDZMOs+9YsvCBDBodldWV
/tAHRMKOuJVC/kxLvqm4mnqypw4ggJtno8KQxA+qj3AczqnyFJbla6qSQapWXiBwsj/xRLbSGOh5
MYDxRjDDY2K1PzkSlvtOnpAssB+LZW1F87Gf/f3S4UlZK7KD+fe5IEMWcdHDlIWDkpaIW0s4CNvL
r/Ldv5MmGy3liq8l7hQQYje1zGEAX0QjoyjDNfbuAULnRvPEA1dP85mIkMJR95XYykcctjhkUTH1
2L1ZKFwD9hPHaPO5/vEGZuCT7ujtIiabeO3JZwMJ2P00Zv/v5AtQBznUxVYWTEdfZudCSk7/uSeL
+fW0p4QbBRspjEiVC6mU5Cn8wLddNO7qsEHqedgSp8WR40EnNNw/4+oWF15txgSlDQtw3bsA2N55
OU0ObElOU82SJmHuvcgVGOtWCcLcpCuncM5EJ2gmJjUZfM5vOOi79nPq+A0f09tbfytJjyMejhb6
0qE6XR60BBhNw3aYRZ7fmr1g3pIsV8OgxLdU54etJStCtyiZXjy+N2CcEzMx8kijiPWUdDE2A9De
4Osj7p2g8YS91T4X/fBQdvD8QPY6urBAOttPWjDjsbY40K/vuFvDhoUcSP3Jo/NNo+J/F/5FOGVy
Fyim42bEvjq5F1q61cq+kaln2mBxvbT2owuFF59s8zu8tN5KqOKmKG8bPnza3tlgpJuKXIsmBmhw
r/5pF6sTit06/cUxsax4A79D9MNEzkSOaiJJOKweN6pcYOERPyNTZmfYsGYZCp88pp4joGSRxKBi
bdeKTiaHuBJ1Jud0SZV2P+xRb1QXI++ul/kfaPSimTU4Q/B0b2cuEvZUGkI8mDey3s26gJy2/hUE
x2w1OeuRGMwe+umgUbqKcZZgyY3tEuya97uYUnGyZL6CZrHLAmE6q7j8CVTTiqs74nFLffgkoPMC
Bh4/qAWyYR88co5L2GtoqQwjWDoX0g8k15KPxevCIqteoK3o3Aw112U88shZ/7dwamG2uHhmflus
mlwJzv4Rh+mr2HooK2fTK1BWvZQGVCHTGv032uEClMzJI7wSH17Jl15G2Xlk7VrzUEVJ0+xHZ65i
tDgWtVYzyKcwpb/5MBb1zOcp9tbMxuR0rxE7oGh/pr3Wsv2Jrf24dHCZ0JTRoPM8gyQCjATIT6n9
7U/cJ1GJ6gxBk+8tDiIEsBbQYyeLZz/92tEDuSA1l2qlE0m8Ah4LCfQA5gJ4faPsJzLCy4H1+jPp
4sHUm+9eb4W86a6T1RJIhyIHVNd+1oyiwY2dy/NDHl+d5AsnchKhEGCDjNu1uKCdF10PMFLfFiuH
kZB9EuqHix7U/64PLSJ3IcMss11+iq0aSEWGgcpZjoIGwyMDrUehjRSy38z19XayX/dHVvGPVjqb
2ymm/FLoDulRSM3hB1nwsSECC7z0/J5MGWsKNkBI/aJ1oh2mh3z6kYcNk6E2t3vf3WB5AW0No0lK
3ROm+WhEhzODgMeZucSGy3nohygy/+plBcSrRgg0O0jsRLPLrgX9mx8P7BmZFzBxQDrZ8BHrZSo9
wdzP+FG8hPaBWO8QSsX5/76zZo9F85AFQsdVLRGkhxUtMItPqaesxNrqKgPpJ+pbVcLdoKTYUmn2
N065zP3J6eA29mXitTqbl7NOgX2IcvedE/xGGUqzMZm4ReMy9ll2opiMG7whu1Db6BvLHVzwTkgO
nLrozF9LUsdruxjXqFVCfZF2bw8dnBNbOtgKimbrv70LSfft/zwK1nASFPRXpj+i8Ld2REU4+nJe
YEHn5gzvvau0PJptZZRtCporozO9Pj2DNniAR1ZpWX666yWW3EN3lRITYUgjn00hnhoFMTbYPkEW
2pBT+j3qpiFFd0NkgAP4DUsue+YcGq/WASqnrSfg3YRiGIu0Un6YBjjiIzBzALGstkfB0ZKGh7bb
5Z5C96vKkq6PWxIRxrjQydm09o1Ay1z7vmA+AJ6qnRWYNBUHEhP5/Y1kwPa4q7JNLAbOyPZsCllS
0ULTVSw5zlUT7FIac/S81HVhHSlggGW0pmY16RkkDLDYeu9IbQzFD+REjlbDQOUCuoqavwRbEYy4
nN5UtOojMTDOX4AWeOmPhiYPafNn7mnmeu649fba4nQ5N9+FX7Pd45ULQ/vJnRWMRN6TGiJRiuK2
LADtVW2r6SMgavtyWWRA22uPqRXQrIfoPrrxn8ee2RA79AW9k9GMCJyM+MYjiVGpjjAmMg3SaMFw
UQMmG+Lwch/Nn50jFvhIu2guCGIaSRxqrCa5VofLieO4u1fywBW+dqpiMKcPk2RJ0JvNiTDpgyIa
w99lhhogoxYE4vf6ktYHVYHZbQZutX39NFAi4LO9I9dZYFF2BXkgYFSAMnEUg4feq6zmOLfEKTz0
NSHNZ3rNkn68FWt0+xmnW/clrvTVvmSQcD9h+cEfA/oCnAf98VSF2qJfgZcWY6Nz5uHHs45L1Vcj
T6GjmoAyoDQ65VhgPeSRYPzZa5bADOPSjwUhxb7S1mpJIyxAcZSfBDyd0k7+IVMN4ePKzWio1f42
wbUF2A3+C5F4doXB3vxvxNmf5v/VQf612Q1rqwOSymr8MYjijhPRi5Py4/ngb0xFili9q//AaB39
eJKCfXwi0+b+/INigL7JAJ/CpQ4SYBNF4kIih7DztWqKB5A0Rx3Y7Ng9X6eaKVgqtAuiQ8gWCrmd
n982uk76ThSxmsGXPR5sKFZnHV4jlfPMaRknWCSqc0P848wv7ZYh0stUhnDXmEnhieMTIEXLZGAb
KFKe5485WU+YWtnNqhAlYzoI8NZAYlYZVg90FtfZnpfFQvtzyOvdbQsDRgT0DjMQnns7QjD5+UVI
ONh5XdvNzg7ADkd34IjSMarkkOjOeRWJeXvRTO8gDNUVGyx+TyCe2ZAMDppMbMXkTxCqIj9GJl6D
bgAovr3ixWK5uvXj3zKBoflzbO+Yrp9Wnesqwnbk8ZFyW/fDifxFIy2b9w3qEPFfmwPutu7H1DEu
VkFEffI0IyJnnRSKsFnjI8BROSo/QtHfHiZMfLwEf4an+xRzP06wbfqrCRKWZ/FVTsU74wQ2hGkp
tHOffYpRc7CtjlfbeWDXSyljIkO98rdVYsYqtMP14j3D2ss+I4ANU8pV08VbXdHmy0UcVlV+9tBK
o+6GYFrO0AyRooBDp+7pXZri8xMpw3yWy/L6k5Sf/iZyZ6lAHD4v3dez7gtK5zjiGm5hZhYPP35n
83r3PBR26kOqsQVf4Hhl7mBoGNsNLVvDqEMnKIq70KcnAk/vDe8TrLGw6sZ3cvH7/GMJ1n81W1Ju
92/YW9lVwZoov7TISR3zR24We2Wjk6yyyp+ssCqWXwA1MRnEFNjHD8ZRm7AHoOlN6vNy1NH/LwDF
TWmu5n9fDZiIMQIuSJqmnvHtqORhifDa948vJTaUQ6CwWNWaQHhM3QYOhlgt289w29opqzPnMdhn
HpozDaQcObYeEOCiYv36A1pFCbOP/LBCqmm8PThjEVoOMmwPHacfdM6sj+o5op1tddsam6uoyLFW
UMM5JzUpVl/7/6slJAgrSjeM4uIXhdR8DkV/mtZSdXlNOS25njf6t6rOO+lDg13OhY86mSVb5Dxg
TmjpdzbIXJucw77d3AEIC4Fio4CVeDn/MWk85vSxNfI2VaAc1e2osggCZvNgPOw2xT3K3CsP1nrk
lLAY7JNis+TS8mzA7ATn03uU0SPr40Ox/rssBG3aL5ub7ZdzJPGQSdM1O/b9qOObyAHarnm0BtXT
pMpARADHQ1+lc7wwvMATdqyV7WBwUZmhigQYk596w0CuHI47d5XWbMfMdLcKJ/JfeK9qy/xKIOXU
lwbhkFj9vAvb9AcCd7Fn+2GLe42a27h+TyAeovSXJn05BzCSkdyJBnF3spU+BruTahREexeWLVnl
+CT6CvEcYRNfT3BlzeRadymbxyRbUMIJZZJUbOSTYBNL7iabWgSq5o6qrB2CQCjHiFG99s60x5t1
5sDtwBuUcsuMKzh1qQHBYg81rQnvpwnP8afr/vOjeWOC2EJx6Q4dr1EIoAW26uHemUbvKAysoiJO
zkYBvuTH9K8tzs4Mq8h+wsExw0vnybZHUAp3NGf1+FcwNpxX+dzuvJwXGedyWe0P8EwSmsqBzujV
oWwcsRIZKFkimH81F8xWAbuINYX3kbAHqyW/RrPyQDG2+CEb4hH4vLnuCS7A/agQWa9mzndzfBnl
bpVezk0vJ5wsB+6rnmOwySsNrCCflGZC06NN3JbihCGmf/7/rHxq4433zoffNOsVIRDxDDetOumN
QA6SAfS767ltyiIUO++5ImGx1ptKNIzYkhtdcX1FF9TzN6O6H8c1oyr7Y1CmvKfvuzlxzNgGMSap
lVTqyJ2lEIhVK6Xqb2ZDV45yxfZpBBSBlMmNk7f8k0eCBBeVluu5QhS3qFMreuMmOAhRHuA3YMHj
srhhdyjiiCPybMEsoif3Hx/K4EaT3DbeEvnn99wJmf86HppLWH/zlA7OPCCavLXgZ4padcG4DsYF
zeFRsiZj4ELV9dPVW+s9r5lY9MFY9S8a7bfzX1uaFOmS5iMyrOAbGRfig7VeMToyFPwaegNmfYs1
rmUK3qY6hK9GM5z8UjXl7b5miSpEbVMT7QkKph3wsFLEpV9cmAWDWXMl8eCljz+E2Ds+0CKs75cL
QKeiRMYLkDkNl++22/04E5AcmOVaSU3R3d0l24Df/U3deaOWn0lG/h0ChT7mVtffEmehNVDAtXmQ
Ny52NKraMfRDDvrUWsvCw8ILA7IgMTjjUXcXWZfQ/uNpcuRdmySnjqHv32rg92oh+WXNtqfbmLLg
cZ4jdZpWCsH1h+G2F0eC+llypMUZEu+iUSIheBOt0h+zNZgTOK4VZ/csFnS/Ss0GbZdvwH9dSwQZ
EYDK61dfQekikxsmhbPQFZ9CkFOXhJFR7SIhzbdXlcdNZ28YKeXQ1Xsivd0PAqWeBL1vrvW4HicB
sBwEA/3TLOMoG0pHvjev+wKxx5BPBGghOr8UKs/ZiwsUwdNImiFTsDXjDGyDFRvfgOYslihlHtfD
JfDLpAi+9tfcIRpik3YYMr9KVWZMhoZMlFRXwK0xbh77QLRpsqxM6cOVWphkSwz2Cc6Ta/0cIIvZ
RQ2oZ3VXAqtAwWcfWgRyimVyzk9dXJnIAWFHNGx45dN1EvBTb7b7tw525Sd/u3PImtfMMjGp5e50
AWCx3pd3XKCbrXdDZheRJZhFBugB8nUsQVCyEB0kYZjncfTqOoFHr2bxAqxhF7iz+EzWAMOdGMeH
MkcYQwtofOtBPCN+Jr1O4hoaqnX45ztuCfJaQZYzzBLYWED9XIv7RXOUQQrb1bDGalgzD2KPiGM+
bVAdQQ6cNVxgr+7STNe3T72vhfEHyBdWovA4yhushDNnU//y6PJ4b7xoViKa0MA2Z+/phOaLbFgl
7tl9aZyfecy04gut7P5VEbgB3RU/Ppi3ziK/4mbetMa5PsgQNPR3UoolJLNkWvTU8iZHRWaxptxR
qiUZrDVEMfeQM2K01LlgRYtUcs3HA4fToXNKYd2AGFttceJqsbq2k5HAF4bgkrxV8+8G8ezIUDDD
mw+lKcJEpp8ujZvv4m23NuhWe5CkHbXpHfXkrlmbWLnNkcJK+uskZR2pjZQBc/TBetZbUpfC5bb6
488WhPRd4I6zEdtYNCQTLLvm7dxUzQDaJAWA7DuwHR3A0tOZSpCgFw88sRI8nLrEAAzEUkN4vLzc
gTkyjWZmrL1179MbFhnGeETTAK9mNKsA021jbrZxWmFOOp4e5vLjziAqz8h2MdXg2KSJkerZO4ba
bDW6uE5YyFJYvHVkmJUyIYQ2+GsHdRtYHuqUMEx2/WhKWMrOg7ITUEP4kJrP8O/VohIkhV70xsP6
O0s1LBpbU4kI5CzTCkshNHo8+Xk6IYQz1ScCzS6Uuv+O2jh1rA8y9Kea9lzmCmu5mZjmrRnSmUWB
dXg7QBouvj7hLrv8e2W5Sgxeb0XxVv3aGI4FoZ6uCfF0/nrEGUHH9EUy6VwrvStMgNoiJpI2mDiU
2EJXL995AQ/QXvbJxnKijTEkZKlHzfg9bRw2hatw+BclS7+5GrYg4BgEXJarNPSrJJctBmMwsVvb
e1DjLohCBl6Cy4CTC4NbFicbqi4GA6UbGw18x1PGw6NNAo+oi8gdgqNgY5lXAvWz2Hm2TmvKV/vj
A4qCDSQ2GZvSWrdJw3TL++WFbzv3NFwBLcQDcNDcPLan+FC4whWY/vb3QwwyMlsJJlTvoTLI9Nti
VrpLxIYuKNq/RMJhNvpIj1Mw/4zaTxCa0R1ejQ5wCEdyITO6V6+/8VCb/OvEQDb5Umoj/LbZKS54
iCVJuUXueSqQCLxuGvLAxQuGgOGLOG5Mx0KPkfF040jHCQC9Xpc/D2HCmoZ7zWk1+6Fs5CYTkUaZ
HfzmWDTfJL7HA0oCou5jLJDgPPIz4/gNJ6nZCZe+CkSaesbGOuW0AtgbHQBczRwmsyHLtITGbaug
uC/gLQFLHh3x28SZuX7boPGOgt6kD2ktER1B6g3SVCIkZjnN4dchWYPVVNeCjvsPMbHgXabyQLoj
lSS8035xx9dOOICzl3CZUYhrmGd4VN2oUKeFynGdDd2cKaxt7tGu1tGqAlfFf9trVhvufV/gjqxp
hBwazBIx+vXt8ICVS3vSdqmoOIA5y0sjY9SIbAhFENYU0DuplVNOyJh+wUlQG+je43F2Azm8EASL
qwcemkIPTe8zHLnTIZhFf6qUQueNkDDTUvLlKr9iywPKfMTKDIC9c0yraywc9YK4X2NE2fv6W90D
6KBOI+cSJSfOiAkMn4RmTNOQ+z5bTzPltKffqv9bg/xiLkuLpYbcaQU8NGq59Rmybmr40WCZppSu
Uy3U7/LLzcmSS2w+7Rp4CaiKrzjAwxHVy9AeDBG0zDn9Mk6hG/y3dtKkXjCQG8Js0vsBv2HgIbRg
S+JdwcREuz61oSHF6mdsHj50WJlXuC5LHYEWsKzTn+PMF5eLKBv+7WAuv1/RT+ogJfczm05PtAvV
Icq5YgFmdBjHVd/f5PVW2ZZr4wkDL4WMlvQhfbS1XaAlPU9Y2CR2zOgghFErm5sD40yVARUIItSF
UQ+yru6EmtX2T5Drrczw+fPbiXGJcryx8pW2ZLF0htvcNLrwLmy8G7ACqQfkMuO3gz13zRrMG25Y
51Z+nysN/aMhRf8elbVBVFHNDkOBjoB9PW9jFXijiZNCqm86gfqwz2seWrOEj19QedUvKphpBwTZ
VUtk0tkLI4N1XKRcq8m1hxzXksIMxq8e/EY2IdXIP15K/NzULDM8yE3B4h/dRr0bHmRJJQ5lYtU/
yJ9Stc35loOfJZ5j2QOya024BwTWKZTig13eBVWO8Xb1KO/bxOf1HmXhX1QLUay4/f+cjgp60gHH
gGDtQiUX0IlYgfjFOncQHV+UzCZkpeeylGeKrUEayoguWEZ7abWA3T2xHm7y1IPHuqXpWUFH4eTN
undldUB+pLwXRNa9EFn9Uf51uqv6HJnaf2h2YBBZmCFvMFXOhhdBaiQRDI2EiQRCUWqwsiG0uvSG
scIaP2/u8ehPmkO1ElHtuGVdqu/ghdIvuwLDCyjZRpyFoewfjD5HAMt6o/UMAcEnf0viK9GKIOfd
6BRl4+L1UzGR2mrPpuN2zUPFYt0rN+iFzbNAFDv6KHdM3OsskWR75HFXEZa+a74niFruTZB1aYu8
VMoEU8NAqW8PsCdppXUK7lIPxQdYjRwwIGqZ8/7psPpr9y/MtKIzp4CX6G9OgmmatVAC/P0atqF6
pHIT5XaTUq5QzNbHYQQGE8U5s3/Ovv6gDEBD5yaA+pZANzu2idDY0ZW2m8S37oo4JgaJEilGguCk
AJ+rpO0nl7/gUj2nQNMCopCuVsFXSZ9R4634eTrCoPirVXxybfB5fX34gdcgteqn3fGzQnI8Ld2e
wzEgK+Y/1rkK6JqzUsr8FPgrxnf8I+bYAoNZ0mjfe1VeXUxk+/D8inBrUybjVu6XwmrXNLhoc50f
1C6AQBWKwzipB/X1vSimRsvzdIOHBuf0AV7hJn/uRNQFEv49GRhprr8bF5C5JOo+Q/MQHiujU0gB
/qY0wMEPet5HoRwx1UR9VLmOzy1HWt9TPl4dayB75NYSzawlfLYn7MK++7F+TUwJYmsnawofcFt2
nyu0soRe7jxBz/rL3cwWsA/jR+Nexdo3Mjgux9/XwlmtDneUpGOgN/gDr8U630iVI0kJPq3If0YE
ZoHcNrwMXhxEzTT+t6Mw6fPn6F+jEHIZLw+lUVPJimgjBb4rdOLvR+oTqKwWhpy519OIbvIxYdsc
M8aq2E5ag1vRFXJtiqgMA/ClzR1veKQbKiXl0yV+G5EAmHEu8zboTYUq6Z34FVbj7duYETFiq12T
zAXFUd0JbctKVMKdGhmpz8BUn1RH6Vpl/7iMLuQrBy+k5KYhYWRLvYjY8sO0aIQis22/lqQPCrQL
Us9XRGtZTn1Q8BOQ9dgTs4X6u0ef9hHYu2VvfNv1PbIRAvCrMiWRF28eu2jy2FKR5Ow28+xtQuWg
OOMZ1dXpSYMRGOsd+NGc0ZAJ97HYgtVjuxhdskqSJeUotCW9Nfnof1dAu4LaFHNFVgQ1hnEIlT2J
rMtJsjnmycW/7yHatJZ150b+yofrMkudFz/LoOu2ThbM8lJhUjp/iXigVYbVmETH3lkjh71Mjpmt
OOxYmr/IAqy0i5xiA9xNaoEy8cnHiC12vPGPv6cGQav9mADb+gwHB+WrNKBtlsgkoy0OJe2G8NiG
k5Luvdl/Xt2aYa97HIsEYa5tCqNtWV542GgOYLohcgyOx1bna42TJLR+J65OREAUiUm2qirFuv0g
UHplJhfVxOlf4DE+NYJK32xeJCOFP60ZCwV8UIPAtKJudq1eh1xFwaZh545bpwxxmwKGCGHC1QEf
t8TYjvp8kziiPBLP3D99tHfSZCr9RiaMXIDfJDmnnxCELdHVvr8wdKQZ8K6AUy9kW+OiST7yhl/9
vQRLaU0Iow9w3yoKqk0kt5lWc8hLhibFFwJq1zhCXS4yfYv/dR/US/ixeLpFIYno6Ig2fJF117FP
pnKXJ/6qWEZJ87PYcys73aM/03unnQH4NqocAhVr8vHhqKIi/gSfbH0fml+oqG9jOFl4VWhBI+zI
5hU9AicsmqhCgFpybuMV8ZGRU/vQcDlwoG/LVB5FQ+KixpPf2Ekf+Go+XJ9hm5s85PZJLq+tagAo
nPiUa66nAnS6ooFcxU1pzHBnrdWlbb79/69LA6lJzRYllR+761LP08EgktwEazzaeJhVffashqTr
FeC2vdUDcb28IW7VJoeN5QFn6cKPoYTCDPpLB+GvBIjBLzs0/m275RHpgYLHiHvDr5IIGDB6lgsV
LHoiJsN9C9cN+fHFshtp9AghwwPVXZ8hZD1K0EGlWs8fYk0Ln9b0pa/dx2sIGMVx2CzlBhnNmcjT
vBcewIxasEVcOTMaQbcDEaQ1VZx1ZBOdOXZntZ4ZCrGJjp9oZcrZvtficyO6Hsv6jpyk9tB5nHsW
i4eVZpywwIzzhIgbn2A1PaYFdx1FIkj9sLyqGAbTSNqmzgwG16svJ1XaPla3QtRvrRditiB32qYj
p2NHf3YE24FPu5PJU0vmPyUXto1w636UoFU5GxuQraHyfS8+NI/o8HIz7gl9sPEkueKkXXaZFj/5
q0D+9vsvKhass0EfnobSWiI4bGqjwSqwkSC1pFO3HfZ/Zy9RvP3OjMKeFrrOcYm6Afq6X9x3Uhqk
sBRuYot3v0rok+WFbykIFX/Kdn4D67woZ9rFmrkFnf6o7T6SuJwAJr6mS20qY3CuSauDjSS/4D59
8x7yXSkv0EfaoPl81j7c7LYaCmqNyhIF/gydM3goWc/mG3J2HomEqjNZFAa5TRwFz7bUjYPMndA5
4jJJWqvfVd8Ymq9v6Uj9toLTPatT6NAc3qJ82WkNeUOZusXTV4vhGameKcZ5H3jFSF4+jzw36MgY
Woj6jU31C8P9ZZLwxBRhJ1gbFwRIFnhePyrEwwItdTUyUOqUWnlbS7sNUaaGPe8g3rxALbCpcAFH
v+IeBdIpVTm693m5+y2cmbRJV4IBAhArk3MpWkkj4EdZcrccaDaTuz2bgKNAFcFdAWt8PQ1L2HM/
sMlJaXsafb39UBemfFen3g6vvzkIxHXxH5Ft7PKPgpgFX4Dgr86NAyru1ipdH7tJhp0g2o5RgG1J
BaOFUBnfCanP96M28+9Up6VW08VqeXEMx62uPvbb5Ns3HBqGQZwg3nwpHzpRp9aO0glkTeEU/B5u
UbH2VgzZqhw5E3UOg1kC7j2RjliifCr+0kx+aclRCSp6q4DEFtpo3wRi+9EBJ3geNps+XfxbGKZc
/x8xo8+8nuXXwVLmzc3wlaiiUCK9F1r0nrKIWM5b9XCUG0OAtufTIE+jRhOSS0hLaMYoCW2o+CU+
Q4tc4SlVFdfLQCx+QD565DGFL8Ev1Q3VfRcPwCBNUl4rmmMKJHEBjP11hBV9m2KyKdh9enDHwFwk
HFcCaHURPhT60kH7fGAtnPomOUt/4JCunUuPaqzxvCH8yiyP0pbZUFgD3l0UxuyfeP/9vJw0jwMe
Jr9j5+dt6a4xypkH7d2AtXmWsuZtTGTV8tiX380jhM7si5Isht214FHJYdQ9Aoqmcxe0jdLfnkrW
DMRNBM8STVBFMhiXtnTaB2JIlbHw0IiRrfqFqv1Srpr5hNryxg04YXQ/FTTe+QLX4j/tVI4dKAQq
jH4mrj7gZyRVDAKZ5byi2rwM33sHNJjDOG83TIyTKEXJFay56Oz4Fc78BNp2Y+uvZ8vnRkcX05iw
zYo096VqnTJq32eJVnjxg30TuN2kVJ8+enUHAFDvQKgeveQH9BfPk+2ZEIcZx09X4AOg5jeNL3wc
9xaWlJOIW2k8AWc3d286dReyv3QHywYGiNNZfgGVtmYglujjK/UPB1+UGZbXx4LqlXQrHl7HbTwF
kwfpuRb2eKsfBdW70Vsj7RfXNjDe74ycFk5PV43lzHKIhnvREZed+CRAeKJI22XTpebYtq/l+d3v
D/JgbKfCoh44BRohEkPv7Djm1qVz2LJv7BU49QMy4RBOseXsuSOFaqstmhlyrg6sRxK1KD0Tncji
5K68lwAYQ/nz1JItCx1m0gxJ99R6BLg5+PcFWSPaRvbMpfSdIbRhee8HRmMGgcS6uyrb15yA51OD
5ITCklzkQi9AzOz/5k/mTJgozRa/E+HlUnMoHLnjv7jq8UAW4MCV0uvLuTS6LkTID0/2N3KkA8l7
EOagvgiRzDJJkuCqf5m7aCaCFCsgTJA5VEdKkDKxGdrDq4TNjxaLqAK6z5Q+EUhGJMOGkcgibAYt
uYDK0d5tvUWwBYRQ2y1mtDxa8NffFXI3J/0PDTl04jMkhzLMZ3mwnmTFeSMjy1wNs6G9U/AWWini
j5miOWKcOoDmG68/Tt5V191SnGgys9cqMbJ04Wcf6iWGnFAv8nf2uzynBYEW9uVEwr9UkpvmiTBc
IHO3g5mK8VvRl3enbj1LurrYb8x0tXg/gHTsoGO4aWb2723OQ+z2Og5LYKVuC/LMU4vQ9IdsiROn
YBiuw3iN2JlJgexCZMU0x3U5znBm3rD2BY7aPNqghW2ciJKab1o2f4hfqDQ+LgUgs/D4hhUOZLBx
coWXMVhrTpKqarvJvSQpjMRYqfWnVrbrC4urdDmYOqM0CELHyEISJXrgvkcUvt8xO5m/BoH7R2/Y
HfdpWPektsgaf5Ca8h1XGGhC+qCbs7lnXZ1H3qV1UH8ZqdmUV1nk4SWRFYSTINuct34vKp71Tk1D
Q2JvTZBxTuH6xaJ1E62naJAl1ist1C9j/3JgE0+N7Oi1tshPIfc6jtT+9xvtBqWlKucwZqw03+HT
beNKCvWA69O/dnM+dNrDvFS7DLQcYjTSm0fOGxDL5Kk5XFw+hpxEt+RHjRrels2WJuBqEr3z8G0e
jwbvIo0zNZE+r3/oorjjzAkRA/aImscMHk4iRilg6bVHcg7Gd+VxYSO7w8RWcDe0IAjRwsEcxkPQ
Z2+jSmh4sDA7yZqtLnDEgkARwYu3WkaVT/exVd6itLiTBmLO17tmHy5AttEZUP0+32S9Yekg347M
EVxjeAFotdrMyQhUdOSAJlVL0rihrWZtqV2nL8JmMGE24dzPYyvqn8ltF9JaGKmQgbEQoocFpxao
JNoJk5PM8eGjb7sUF2Dhjklm6gPuu/HDbnmfAPCj69fUQCGRV+9uT0tRWwxqjA4zx2+M2/QQcnuR
nj4jTCWxJZ+kT4VswJxkSdBXcQGt3FQyp/a1yChjdgbxjQ5uQO7cj7hNiMFJTtm0lQj2UXnSW2d2
TOuJ8Toz40/NNBB0dWH0o38VAcwtiChuIwYyf85K0abHIzBARFCZNO9orUjN0kUXchPVVvhTy2Lj
UvxiLbRQ6Bwnx3ngeYGOYwM4Vf8RvTyeaWGXjZkGJPMK+0NZjvWqvfxdyhnpOe0+boNrHtH2l0aq
SsW7LbREnIff1d5Kzon3gdCVwV/OIeko0+3SQn1XZ3ph4dLdh/t4SvwOKKyfw9xpizKhdoAzARl0
LsIPXuxDy7nVRWhO11vllvvwYUFF2/tuwHbgybf6lQ/JsvFssF8dwUhOcWsG/ATfXPCuT7BwLF4B
ZYS/m5rLgVmkZFGc8u63L7QHEgqBKS3YRY4v+hh+v+fKoU1D/rOM/2SvuUD98WwlzY32JEo8o/vb
bWDSXc0a4n74l4KpKEvvwoj9t/D2DfwgvgOnZcTXQ/WzHCwOMU7KfQCEAo3gJhMbkv3zuLDRYYgu
X+dJqFBF+NMIZsJYmC59zDh9BUYsQoXN4JiChO2u400iGsTiIfcFk4MQ3Gl3qSiLnDpGgsxv5g5Z
6IyQqDSXXGBFxplDaIoLGQpdYdz3Rh34TyyJ2KEYE9UJogQntDw2C8q5ca5MqSqdTn1ictIz50dt
G+tbMKP+BSvO+a208GOt5cgFpi+LClV51h8XTZ0HuwplrlwP6Z+65zpSwgiCVkdignoIvFDkzSVB
3QteLN2FXIkC3uezbgBkT4j6p+3gz6PrlI8X4rG76jcjBii4PtUaRuVug6bluFsR8nO2G3Pf1q+k
Re+2AosPGYlXC+M6KBMzh+md9zLSx2FXO8s5t+fRRfKca34BADGHGbdzMc9RpBVxvpJtTdW8pZp1
Jwhk8m57iyiazt+wVXrI9D9svi94YyP+wVtEHx8rZ9qvnAV7mswPN/QbQZjpHGUA7pRTueT4NRmp
eoXCEjpd23WZWbIoXFv77ywx8UAzxIKWSEQUkBtTZjG5BflLwcooaErorjfdbJwyUsRx9+ujtpXf
ArkVIYEb5xfHEYQ6bxuVzD/by1WDDAdCazEuIe0Gh9m+bh6k0pon04T/VrkQkP5hMxESK2In4x8r
UlfTfxLd+SS25DbjKKvFBYaeYYNyCfxxfH8WQrGkQuNc7xzJp0rEZ6fVP/ue5bcELwXb9vcn82tv
rDThmohl2U/Azn7xDPv4kZl5fXzOw4f9TOGbs47RkEsaQMvJ9MPeSSJia91iVTzrUxj46T77zLey
WI75/Z1QHxc0SRTsbun7uAeURupNoDBmoHHlumoSPLa2sCKT/aelRt5I3CUxvV65aRdG8NGHwMQS
L0f64IW0LClM3azVJKT1rIdcJlXvGvIsbP4g+A7Dj+x6KfE6EM4y6SMGPnkw/1fu/FXmMtd9MH79
6BwkXVGC7llI8Euk2Vr6r72iXuMIv7PbE7plz2JjoBorc5qYPpt8+KLmGA7TDIusMfaLDoXasJzs
7rG5c0t2MZoqXEzKkVLRLbKQd2/5ZOXltG4GiGhyEmdrbe8NMbIUfxa/3v7YnmVFHavmfr161oz9
OBoNOvhBFANSq3AWVk2ZaATBw22dM6YqILdV6vv2X+YXpRdkPjHF6xk8cVa0FTUjMCRCqECbR6pf
4NT8LyaNl0Jj71esJ7J7BzSJi7gd6pdvwz0Q+NjULsQoIrWyFmjikfTTvWQE1n8BjUn9RRcSZipz
HJ1Hnn0uDDCAX+mZh5TCm7kEVwgNK7rDX+yWhopr89mcxS6UY7T3m9OABBAwjBbbPwSR33XnQq6+
7/vTpnM2E3MvoXOF52110TcPbfnNzf2SNYm3P3aDgM8pvuPC5SNeESHRxWu2Cdqr0FSQDFMnCnJp
Sf02RTLE99SAWKbAOnWW2OnlNEAa1SqFF9aJc58LkZUldamxAObF5tgBRzCwcXvYXq6voNtOrmfd
Lxl+m8W4R9CJvZjq+ffCSdmJtipnE4wqAdBVgQY0MrDuDBqrl0xUQsNt6JKRzZW9AN+8C3L79gt1
zl4kDnh6Q2juFs/LZU5YdaIhy5XB+oJexKAwaWyxTjcQWtg5J9UtgGP91/lWtgQ9Iae9YADrvNud
j0OVsx4Fwk8SfgNLeaTi8rtF0BvlY3GLNdvza7TedRwF4XfTOgqjnIoriGcFlCwHeFO3M8O+efK9
1jaaM6jeHbRu/yH0Ezg03eALZ+K8fj5TSYSHb+dlko3klE6/KmhZMN8UhUdNWirwzjsJaZpEBbdt
VQurU5IrkQ/JQXwhCJRoM+N0BOUtbtA7OAGx4SoGvBodZH8bGLHn5kfeSr7AYAHbs+ofNKOTQm65
CQaDH0xepdgR65fQIe74DBsQuV/NDKEPLaDE/r+rTB8U9SZzT7MML1R9o4Rmky7gea1FV7CaHV/F
ih3voqdYkFyU3iqd5cUgtIWhSsR35GOcWsAuf7JCBEeZEp7+fjScF72r9xprxPXnBdbfFLBL5goS
pfzEwzuxmt4fK/TtQdTs5USO6ErjCCGEZ6W4ZCuBUqPGV0m8l6Jlxh3EVkj7EuluKnMrOawlj6fy
Q6uggPmiPyGYuQZPMexvUMi7t6WSIASBE0MGxoVUju0SRmNJXtBEDFcAnk0DbKfT0LyFUHgwa0Od
6409AnVtOdCdqPCXyM/3pVUcNO3RefwzN28Zs0b7XWw1baXvM3Wxz/uY3hZyKh7ZRViAqll6SYZF
kCZkfxhBKU/fsuWO7bRKIG+FZAsUvtmJEeBlYi3iO4Sqn71ETgD51/+6M0SYUzA6fhEfKg8+BGBP
4el7pwUbi2xaVjvCzq+JYCu5F4TAU3Ut/NoNyq/l/At68EDYGm1dq8euZgZDnxe4W2h5jEfyqH+8
qQ1MS4/5p/iDHMvdwvsF28osokPOMyJ9KBwTjg+bgUhkPNx0tge4GUkPiO6ubs1/EPzOrXCGkzAQ
CEskz/WYxosjpJUAPNS3vTXtGRMsaMUAL5WrbNCM5MC7e6V8AZowxYRpNN1t/T7ItyuFRHQwbqWW
pM1a/M4F9/9J0nH0kSX7VhhEjLShlKPEQUYez+umICUaMsp3XY1tc3vZLEBF5+rdXM9I3jGkXzWW
SCPWCepge8aVBh/ZN/GQ3WcD4X3dJEr45ZidfJSYmmfcJy3gPklAZGqRP1Yo37DNIOwArOgMOlgI
Xy/+TKc7JioHc4+H0yxbgDYYTukAYTrWhiw8alwx1xrDjNVWiweD9fkMkadOe89Hsv9WyW2a6B86
aSD9o7NjokCNANJR0zUZ/0yMOQPy8PViv/IBNVOTuXhuzn9y3UtnbsoEWLLkUKukTWigk2V9VKuB
hcLD5NEteKpqFAkMLJLSsqG+h3rU64s1anir8icoaKfZ1nu+IZ/KmX8X235EV4/GHgrGnOeU5BaQ
bOlp5hsI5ZISbpXDDqPTB30LCxWdwmcS07UHhAr7nC0suQ3Ix6ryeEevUpCefJqNNADbLoU6ma8J
DySL+WfEWeL31lmf9kSkCWb/0ZwB3IgOgIlyd6runBaZxaexuY0QeazyyozsJBwO0uzjD3OeOzib
rnDwDSYDQgb+FZzqtbAXzKpzpnik+C6oEoM7vKZPAe0mUN5380cAMY6AtyG4w/O9JlNyYkowp13K
h1ECbqhodrXWH9vL9l9d/7s2Opcqj64YGFXeZAzLBbwlQ7a/CeskdLDC23M441YO/AIkkgh+XwPO
i06wjf5FjbS4xi2om7gWdyDlSApDCoegQZ2DnMNDQZ0u3AEM2DoFdXgIsErBbFcUY7hJ0tO+6+xm
ob9RRkAUHG0xIboudcz89iaKcn/zlHrTJ5KGma1jt5WgUwB7nAdjqENQzR6/DYvAPWp6xm4fRZ4D
N3hp99/vbpIxyh2uAezD+Njl5vcp45nzk7hvcjDYCWuGuPDWkXbZpWN/Oi6slmcWUzXNEd8LqgKn
7l496VlL8V/c/fOF1AepaCsSQkd3p0cVcJHJ0dADrEpVGjMoOTqCwGYjVBRWi5EkUQQewV9YKbs3
91BtLECIDqxOIHljReqULGM5Wrjrzid4gELbQtGP/lJazAFkPlyzOfKVIJGBV6I2iSD4w+Tg+vUW
vGTZ5Ie8T7R8EI5+QP16KYC4nvdpOcYu9q6wYqdhZxivITEpfBdrddqYuGKANWC2iR20PWvinGYA
30oKwBK3lAlZ7uIwZiJJnx7JuR3I3E/O5ABsSg0oAs4vXl90tLZ/xVZ3kQIj2HHS1AmnoY5ODJFj
F9Fh55wOVBlxubn4H4yhmQHWVLh9rSeWeJQEjJF/DehifnGbAtYtW1P0D7HqEpI4gm0lCsnDvLtF
tkZ2goOwtqtUJoaFBTd3hGqzDWM9Q0aVlhJq8Zd1E5nMRCB6grnblbYMWH8PPl7cjvdS3026ljy3
BqLj1VHHY9GdIdnS9bUiUv0Gw1Q+RydsLvNzqaEQD9b2ypYamZ/RE/CMyhte8cTaPnCfw+mDlCUA
3cOt5n6QVO5FPxnSaHpvjaMt5z9gCsJ1VW8y6c+5Rv9JfuDfgtXgkjCmkKiWUjoXTCos1iKxp6cS
bzJ4NAI5oMq4KJN/qAtRJMpCD/+TcZ6+4YDvsXeyr5u9ZKBA9fCRNZrE8Pl8HJ3cZkCYS6DtTGF1
SNlLgJgSGF1CZKVtrllrwvrm9IUDK+cp97eMT8lC+PV30cy+fjQgZY+HBOeW0W4/h6qVc3/yyqgl
Y+3pi0E9VsMed/oIx47rwZfyowimusm+hEPkS30vxgErL9tF/V3Kot47pnTOQmqRe7BYxzaSv0qe
8Tet0bXEPfcBVOWtfVsg46YO/7aM1zoibxyXb9G2VdOF84+ncFV8RYKxG5Wlf7Nmby+G21iBmLCT
yZZ8AL7v8SE85CXoT1TZY28gh73eJN0nMvOMPtz6dm3G0NyC/m52zKlZoupP0a7mOWd4P4R0Iwt8
1+pPZSa3Ocnn2T4iRXjIqOineNfspsyoGBq4AguvBDIT1ZJfw/MQeW852JlcMQORQu+zljvGTqtv
bkKRiHftkjRWsA1UaJpLry7kfYpwCgUmBkq4xRC4R9oIy9czOF4ktmOZJiFLx8kuJsbeXQuAQ11G
M9ifW9OY+guOD65cI0poga8zDct1U1AW+2UDNzTT6NrhooCZqYeEkqOyZ+ZhwMlRGQSaEHCF73Ht
CIWfBRK/NiZMWvCv3jn34V51Ocrung64LxW7SD/8hdFy75JifEn8OHGQvqBpHYv2K9ExFQVja+/2
Wa9ogXbDGakp7js2JTJnO/e2en1y+AYZKlkKdTfC8vkQD7ESxUZnoJiUnjTlZXVxLJuhFxQkY1bp
iULbAwfyZo6Q6LuD1dBflsTA77G8G+xR9nExfodzOpdpF5ut4o5SfWam9ZASBTJ3VKOpMxLmU4cU
Ldx6qrDoeKwaaZ1Q3a0kfciCsM061Hv/uJk3wTM79PnmRajHZwbGE8JA0vTey2886OcRgdgjGKxG
bbBZ33hEJ8VRqZK+IQiWp7IlQH5EoptlT50wENlICIWedrxml+EifmZhYTJhmqsCLnZOwtTaM3P3
FZTSLH9ggCem/D6hZYYS5QvlI4OHr1R2HArEOK3e/YlBJwRwW352Wh1IHnCmWNDWZn9vgIZijgYX
tmphV693SLShbPdNliVFadIfXbNHihJ722HxE+C4kFefnohv5aYP4RXHZPV3/Cs9fo1TyYvU8Xr4
9oH/UUg1P4Ote2zq71YjyhdRa54llAIWW6gkD6zU/w72YNvR+mP50QcIvs27psmgggW/lFTiTrhI
wHpkn8uov67D5xEk/9Wn0RcXDpQTLYVd0ebAun/iTc+WAATbYYkdwGOJC73611/7h2f9qyP2YoZ2
4NBvbRPpDKNEhXWkY0tKZjG/GjRCsgmxxvDEJh1SMpvxLOk3rvgdDypuziox0k56YoI+cAcMqi6V
d+V5rIYhQILgxeJNVe8to8b6agkmgrdUF8wtezWwdWTBF/Xx1sZVAl6bABOP1kSaY1Hn3ntppN7b
uGlC0ZOvbLrolGNwuMxSEoXGI3G21qXL/J9l2gthSvMp/6zU8OUSK31mdnUO5rlO4sV41IgVxBPm
1huJyGBFtnzp/Xh0yVxXVb6e4nrDBh+geiasLfOkRly1nN16EmzuXW24/A4nB8bv/qjGqoo4SU48
qwYmZfrwf6cEHvfozW9IYGjQAsuQ+c9QoC9XsXG8J2d7V4WadLdRMUFq+or/sGFEh8gIKtRmIHvU
u0+Dfq/U+Brw76shCX/gPkZ7RfqvvgxSQP0BjIBkYwXOgQEzZKezo4sca0ZLKsXA6n/c//JwDovi
u0QMRCMIYduAdJ+09eN/YF3rXWhjIFEHteUyrbboMSCfqjRDNP/R/zj96C3WrvxFkQKHAhf+npiS
Eri7ub7eote1tnlqNNSxcBkoqF3Y+CbBKfIeKp1B5+wOgCShyaG2VXy/sfehA45wmnh5UcJZD91U
zLE3FcTrEgyE+7Y1aJgFAzbhYROF6Clp9TtpYxWMGz7cSAxeewwaQW7pXRv0cyvCPT24LkN9xA9f
WjgEgqtP0m6Qd3IvUqLdont8+4oaKXzUfd8ijLVNyNu6OsSWLQxRaA4pq8FJUtt7eoThxfBMurIW
3NDTXiGYyaSp88oARnoejgBVu4kh/IcbjalKrUwNa54Gpw5VT1+OE6atTbuhjGfkxAaSuky7Nnc0
zWoh8Vyxv91p81KHkpm9WzLg1mD+7gIqQ5r8RmQtapI99Rvk8Q+FAJXKt/Y+6638tFQa4QMvhg/m
B5k00mHarI+N0J2OWby3xLNYTi0ampm4B8BjwstujgD01R2LkjXMt9/U3tp+Ya4za1uBdIlEq2kv
f9ZcdyK6OvPds27RYwDOimb5IZHO+7tNOsK5aI7UFSDBjYM7sdKQID6OFQpA1vL9JrWEtStkDs9t
HjFaW7JL/HQWPBoZZi1obRYcGrJOMXIO9YzjdVQhmoPZPGjiOgD9WwRVnCe+K1pn3ojKv5snYyhb
u+YQ4Mh7N2nz9+fTvewf6fp4zd45Bi31opXw0CYxTXoMr9ezuq0nSPMQsX8Ql7A7a+CSCgQBZZuY
/Ak50RT4mSXcMmtSMuVC9MBCUEQufc+Un/E/phsbbQ3GnREE38tObkcvg2S+5DLlIJ/0vpHrcUpj
iqz7dcRd+TfDqKhJNVU2ZpRhqZrnVotlPvneSjvfjxlQsuX/rSR0QysYjSXPGZ3LqerAQQmBSjII
HqVbmCycMZlCSELRqwcDP0whkAboe7sRt9QUqSRqSG2e2Q7MszZpsuSgwtJOYqpPtgWVfsVMnpzk
78Mf6Gc2kQoj8c4rxe/Xr5sdFdx9UzgK2vMvEJh+yI6IKFlnXrX4LWYI6D5iXGBKFKlTdaLGnszq
ZYw2ozeNuXeMpC2FYdQSpB0bYy22ttxGWtPm8zYnVKXYPLrFB5l7vJClqll7X1a4NY2BER1x3z8m
LF3bLKn7vvcl6TWyMpunPRfjWcTLsfuCeICz5pfKb36iQuOQ+jxXFf0nEwiQBuBl7idFqTFCssSF
+49AR/VQRTERt3GTcy+pdJI/ZeUGl/kYVajZNG+TKf6JExlTvjFnWlOhYnp6OZ0KnTMj03GyB41E
OQk0yHCz+fQmGoYAsoknflXb83+JOAA6OadrbU1F05Y8zZ0bfatj+COcVZEGLGOBRB/g5h+groMr
raul/I851z3U+R9yCAUmLmhuZOCms3BXFMrOb0o2aWXN8rKfNaImyCqyg+4sF76AdE+zH6/Q0SRI
1rHStZBenbYc7fcniYvMzOALJYkHhiBMDb5HIi8XLjGD5sb+t+qjhS81/5DPBAQteH+CPv3Nar6s
PR3TK5nbpJlBUu345rq7Jlf1eekDv6dB1OK0XZkfp/0wa4ixjbsGtuvdh11Fnll5lJ04H7YiiJ45
s/F2UkDXa8muT0M5sn/yw0OCBepctPAwdKbTJ2/uK5dO3IX5C0T1DKJQTtddl+/DvZczsul/nSdF
OByIIwj9G91e/g7gQ3X7ZCzbXgjJe1OcOU3/znJ9D9xMS20WrQPd+dJRkapS0/GjOmxv67EgaO17
RGb41/kX2XOD0m8VHiAv9tmkbPF2m5Ic56nI3z+L19leVi06bQcuwU4YVON0Pzdypl8ypysWvy9L
mUsEFFmDXp1DST/boyMjIHqxJ1dHll8UMpAbApqMIPK2I+Lw1Ot4sz4+rrDlDhzzD306Z8Z6tLW8
cNEpWICwzI996G35iNPbLQyNxWvOgi+HErcfS87XyoGz6OoXFnio+cnd2ViYor0AqJ15hgPd3McP
T5gwupHkoVyd0z/nKxC6POn0QbhSMrNH+3Re0iM594sYBhq0qwPb3pxUlgqMsy84/ao4RQVa9Vnq
RuPrD55ZjGKd5Bhl9g2qQAVpKjTekXiY64lgTjT4KViWJg9bbxt3V8okIkJ6Qmb8ON9Ks1m/zz7J
aYBnqMID6WmTKjldyqtZWq21ObIES85mXSR8DorC0/dBG8N39zJjpgMGjLtLUBnpAf+Gs6ZhsGsG
nWk8kpdhMQqruRjnzukvXIFlBcmHovTsrZxZmUTiV+DC9R4CAM5aGKN1Gfhny0ooJYlDhO9ip42S
6fqoKpd+JFjeEMmGOXlg71XgOTqPCOUvqxbRxeozY2iZvU/yyNqAmJV91lVS2d1jogd6ipopwhfE
gnWz6eiBZEtldmXD2sK2Rx2mc8IqBeLn6+9BJc0OAhqj4pREBQUDcbjRa/EZMt+wH/qtyWhkxucL
H/rvzPlaX7y6udbvImZtVPSYv0B+fGGfdDSxVr23nBsih8YJYTo6WfiH/RM6RBX2E1ar43HzSgUI
xRXrmLTTCJ2QbUaYFa8XHjhtJwQlUblI8GwqbTKP+gUfWy/JJcW3M5WHzOTcRWlkPix8N359p/Ke
r5hnaoJxGmfCdnc8roQGo2tl9RpUZ/iLoNWsXCTTFUkjsFiwTY+AiOfaezRWdJfdVYsNS0ohqrNG
UMbURwDtCqK29mNfjn9LS0ECIKgEXuW0PUqRAheGyKnEAMSxZA7iy9tL5i+KGFcYDo84U7kHdmTV
mhLqSGlXfxps8FFWb3YE6vcAPWwVIpAciPshPfxOL5wiLrEEi9Hjzkdr7Ue9KNRi/NYVyzgnVv72
GGnqRP/WsUTfptEHAiZt4bkyQ/dwgCInUGgn/2rUgBtZ5HkJBPbM6HH78cz2VVUBs8AxIskZcETV
FLoq/+RyiAsWm8TL5aiGBKGGrCqhLxP4ihW+uOzrt96OA8x/q01BXbuQ2iw5lMMaWAKa5WZiKPmf
EPcbCjjCUAVgfYtSN2ht4inOYU2/b1t3bkzIusM57B6EK7xDe2b1PF5Nfg1zsZ7bUdQ89arAHBRB
WCIz4XR0u1cdqd+RWZvUtqqvbO8RubdpRUfKLpJx+3LERzBjelMxqzm2yr7XnQENE1CWC/gEsty/
otqwtMbc1eYuUFojFDY16NfloCI0KAhrCru4/6KayT+f/4rr7EwgdqrAGZ5CK7DIHOqJCsYhdkf0
bAlWz1jzwrxusQEaQ5k6M4eN3pFLgKjD6hkHqNkLHMHVNoaMU8Xl3NpU1I/uc+1jSR/unDkNcRW4
Z5k0QW26YUkgPyGGm4Tkqo8kuAs3xubBJ4KPm6mqzE+0NFYVcYQ6DENNn2D0EJy0yTVZkBGP4FVX
+wdMpSMJTcnZ7ZbcBdvnmJeKnuvzvBgxkb8kRkU7F0qPpXLaWLXNwE4kp3om6xU2yXx103gMr4vI
o4JvcKIX4MphITzdtcaJMYB1a5O3R2h3YFbNk3wilVS9yIktl+tgTpdD+mc82HB0jNklRX8+TbYn
9o8NfldB/Cj4bt5WeOS+FzMe1GJe19iksETJLnoseQl766E6x7BQPvK2J8ktk4j0lBPwidNP7YU8
V2J0NEhw3D0IQDCtv/TA4ikZ8IU7iOUEpnUdN4D+bqhd2ghkpu9f7Uz8MXExoYHFlyfW0Lhz7Q8P
dr+O2G5BV7u+CbTPGwVMnkEBkBGHMt49buDlAP2m9qd2uLd+Rjg6Y3XY83+N0vA+VQ2sebMw93KU
wI93dzAQnkktQp1i6oJ549Q+7oM6mNgfYHMAOAA5JYuNLANlRE98jfDdkMrtkDJoZmdVc0xNeJxc
W2e6L0Jwz7BHrISDhYN3KS0FNU7bUIDKDX0oGKZQ3ijicSVzebXS/PepBFpT4D7FbjWoux3BnGF6
+o6CSnhZLSezLL7B0hVZ2TFi96dTcGW9uDVI5Wt99Dy0AMO9BiI07RHRv9z/4yozMoNx/7mQ+iSU
l6gmWZOUt7KfEP2+SjeC+B5q7EjJ2XYEPq/u6wCvTg0pYnukKId7XQoRftp9SESq1JGjSDM3i3V8
+lY+g4b35xB43HCQO0bDbiXyCR3/9FYB2Z+QZIM5BtCSFyQZMX5wvyHATr7JOIPi1hBNbV3HZvam
YygxcpAA9fqUyOi5/M4TWEIc9REi/s6j+QuRL3PcyAUBfwRYHx9u/goX1d6qcHVQ5ptvg3C7OYcN
6LIuXkynuvH2rA6wRUjsUhD5RGjb/YIBU8pyXNhKSY7vcXuMx5HMODAZ7bZwMSAdxYUswPQIet8Z
agkEa7vE4tbWkQ+VBPXKCgJ2qVDS7ApGptVDJmKBz6VHgJZRdphbXQOAu6SFVNuqqgcUehTtJTgC
92bQBPPCHfXCH4fLDI9yYrUUijO76DMvexI5rW/Hg/9U3EI3zHiHiu39Up9SavJakqOhs5VoXhjx
dco45Dweu9lQeX16vImkNmRLuj4tUICt6IXbnD3CWQu+TNYhudyOnHpLemMCXXWMO/9/doKlP2ke
VJU8aTMkGUBHPmcOXA1xMCTdtTKL7AsAm/FlsyFHqlDA+tpis3S60M53lLy0pZVnfEQndl4Z71Sr
+hpvLVWq5dqFOnoPjatZoN5OaqUPm/z/gOIxRDYJ8rI5r65xa2O414T2Wz4ar2ujPFrNEI+vFDt5
GT2VLWOtope7CRV2s9vnf31OZoK+20lVv4q0yWHPhWAHy6LhIW9+VdxwvGWSMAmO2v/FZAC8GfGb
R5duwwc4SC8jw4xxIrU4uRWoCg9HgxGdnceR3MHzbsBDL3Ih+Rale4ycNjltA8Usa/V/c5KaPKLi
RiZYvFebf8EFVW09QHgNp9rI3C/vekOJhP5B2hG04lsUEABdmcHW1BktX3nVOr5bjLwF9yi8ayhn
fzYcRmW2CzyjwhYxqg4HmXWPP2EiuPJRO6QCyVHJc3HFD5jOP6bWPy6mXITgLCEOqwkAIZuEYvGu
LFUBJ+U59zokiqkROLTx932Xz1AEfOZM43Hxez/5kRePSCk9ET34+hmUXmyyxctXdaMk9008B8TR
NLY+xOVnMVdS8xe0V6NEElN7EYWYlNG7TgKPJnkTtjhFile+v9QWYBY26UT0NKSOhuGBCY2PDmaO
NgKLEqpJy+9nf08ZW7pgbQPKa1rQ5kKVAoOx7zabgL3yOBBkdHc7xRlSBvE6ONr6B6Au1XasGsax
FVdDMaDEHTUvDiD9jqzxBKXw2Qhu/hY+9x9fvj2x7+MpM4wW5GezfBnnnKALg3uE8M+L1FRxfr/S
rH1YKg8TG+EwQ+kDZfZKj3HHCw7dX6AJlxNi4nyje4fpytWGvch3HHMYV+KuT3Gj50nM6RpbLtcD
ZQGQb2b5or/7rNnxVtRWKUVhk/0N0kIjhSrleC9sNs9ChricybCLXzHridZy9y3XjRHOgdmxr1DU
MajGfHGWX4k16qpTXfhy0Tu+/RP/uJ48KixfCZqdS21PsrtHczi3f3fSVdUSc/aHWlO/1mjxLQNB
rB79omqykg4Krm6G+hslZ5hIzRXGlEvYcy+ylx1r/Rzv7tfxDvfZE+zXiCXyQUrHd/sFdxi4ax0Y
mCmJLM+WsqKGTds53nsQmfLxlGAOI+CO6noW7+wViqHdm0Qay7E3CkSzxiVNrU9J8zOFz97O76he
AkNUBSdOnzaXSBrPa+j6aNXeRAjsROY8fj1Xsom2jsH/mfR9MbohbOO6qH7X3yUaQ5sitvOea9Mc
cZB2tNSAwc6bcwzh1Y9myBSa4FnbNpFgtGiIjrToUxLBeoe4BFG57Ox/BFvO5XN3WzXFDgUVZxLD
QHP3AekI3Dngy0Pk3t1yrTADSxE+hqf+7rG2NXQA/vhWvM+VO9ppKndn7C8e3Gqf3aZBXr555/Cd
CvWrgSatNZdMCfQkTAJa2I7hl22oyhSMk4grxsE6VPN4QoHVZQeGRbWBYuvjH6ySnByNi8z7gppp
aNRVjWuZrpeUHZT7gNLoC/8f1G37/w/hjRa/7nnSGI8W+JKPu/03O5GcWJg9HTjax131yNAUpfi3
47UmXdq0JqvweVSBGVritAzjaW6zubBoGQszc/RRVNIwwSJ6dxJlGKsXsUhctKMU0MQv+fgaYYZs
PcCf+/KoFahnQF7sF0PsKISOD4Dozv7lhD7NbhtLlkgK0w9e3mr1H33FA1e+juUsUBBc0NfAdjHs
WkxOL6Y3QSOAnjB/uf6OZLrX3ztUC5OvGCrrwLC3Tdf4yAe+7UnSLof+gPGKCzWf5dHSX3mmMyhy
Qpmrn3XGeL710SjtVeyNb5EgN4l+ThGKvvqt5z/AC7qhfPgmtXD5W1/W3ZRBzZW4QRICrwikqnCk
BCb+PyBWgCvka38HkWPvUmIUKeS1VOgc1qOiuGECnURKQ88ywCq8W8n9IEWtQPDnY2K58KmzW5LY
0qNi4IOz78+f9nWXg/gc8hbVfAIUgDktOYr/dfdbzaFRD3lcX0OyecghFNHhQbHCLQtkSerm75Qz
Pa5a1w425Y9bVmxCZAzZdABmrUDi2Kpp1v3PNsFbt9ln7zh935Pt81yfojHFG9rNbvcoFsCiPVEL
nS+KnlyfVSUXaZ7PGrUIBNwF1zbFb3p8Y4e2IKhqRjUPxm93JMjV9mVkJDNB+W5L3+IWKfwmVELz
CtAFOoYp8WJKySYlm1FjkJB1HQN9EAUX8fSM82GxEALNGmPrfv69y6FJ3BmN7XJP9FoSFpxtg6LD
OhjlxzgZv+qSl/g4P7oLBYIyGEuXHi4udHsavTZURsH27jlpEXLmoDMOkRYaWy4+gGjgQ8F5kJtl
vGkOsP65Ps9EzatrA61KV3WSWuwD5p7LC6Yt6xrEhy/WH1ji6rpB9lv6spNvomB5rXf1Dp4vp1+/
3MuSqBQip41UKXAllsM0rK1x3PHHtakh24X7yhpP08fWWjDInAUN1gtTz6gIV2uSF4yrXlA94qh5
2DMVMz6aI07+6hoXhL3iOJKRmzKtpj5vovguz9pbI7Rq17PSOTYrWUTI6ARi8RW9x9cYo2IiBCyF
TV0S3QnBFQ0MdT2UOXGJQnp7A3hs6x93uQUbH4+cd6e3VlDV+RpAVESWByKQv4Gv36h4JG6/mlXL
W6dgBreafJhHoVOqH2QcJzglhtgIpBSDidIAQzRVnqoaXQ7gf+zptmsd+o+kMx3C6Y1KOpQBTNya
zGu84ST9VUz0Z/lbcCxfZG+CaDO+AuBoFT8+VfbLNJ+eP4FXD0xPyI50dugdS3gSpHuD+VU3AbKi
v2gsbmsZLdTMUyexeafupeuD4O/37jWWgNfnXaf+pU4lC8JcoA6mppOqfILxUrx+qIp+XrVrExXX
wJZa4LlgmdLkMJyeqlq8kY1bjtEd+DFw7Ba+B8PxZi7hG56FAKC6xKt/aGNUpekhyEuB6BYhT6Qa
T3Q0LlCOxCrD4csxo3+nqy3a5/O6WYRFfIZmKT6pVpTuO46OPjSIBKTuqqoAM5Hsar8Sz3OA7bZp
DlzpnzBPvz3upxIIa+h2fr95LtmnwmcNLbf2Rj/Wq6Ppuey5uZv+AdJbNN/smZUfhQZt3OhSiGFK
TnjnhZa1SeL4dmO3R2YGh4UTdBeXFwnRBodbYRE6AKD/P4uz7gAw8bV7/pVfL8ZNJeziFCNe8KZR
pIF0qyD8kZooWlzcsPmSyP3dyRr6FcaswmwdCNdEead9YzOMGtz6MAryW5cxmYRZdGH9sfRImbcW
bdvP4XYPtCDkLT5MqYkt5KZhqUrWoA+7K8wThBkzsBu0FwVnlkUVLcROE4e647qHfFjE34rGrnfl
OerbQybiAutbnyWNP88g2wiXc3HemFi3qXzphznVRrQQDs2ElvQ3gm1a6DkwIo8nqRqJw9OKrYzh
jN3JJ+twCLOXcosKiXmcaHv792NHJ63OupyK+/iq+1SoBi6UpLKGUhK5NmQ1TXn1QPEdpCm5/Slv
BmvzMDFmZ7vCQ6Oo8+QGDbnlI1tiLCESdd1mA7sULOOynpe8+Z3kWNb1lo6T50UzP7zG9EVcCy+C
IGNNQXODGXUIfWYfwV7l8s0EEUA0qYgOdghEXO1ZwGnGvvDyQW03qwRQDW3iFqR1hm/oic2CZKUL
TIbsK6zRIZya3XA0I30RQVEmSYXjhPcFOwFW9RFgoCd4NWbh4EXiGa4uM2+buZplsNPDOkYMbG+P
Z7poPDf/1AZ1KlBU8DyXXOd23rqNeOc3mqurhqoQ5AWa3P7r3xG02jrZJHnEvUmeY9kl26YjAO2Q
Ukit5W0i0mxcT/4Xqh9+y9HgURRhmnGRS9/5BN1ZqyTtLLyHXUI0tYd7FjXAExnYxt5t31atflsc
UnICd6JgBXnXWsRm5U9py7GdJjDjXyo8leKqfTOHK/xYkCVfP8S9yl+jMvtLCoSAyqZwkwu/KYNL
X9BEZvhLOeKTqIORGbW8MKFn97nCxYDP+hMA+nM1zQFk6kle+50mOIBqwqD+/Cs9jfk+iX5ukpGq
whILgvM+LBYnXCnaYnw++ppVi9s7Ro03hoop2o9KIl8bdVYKa58RudAzswqWKikd2i8csz5znPse
0n+WkIjdjDg5QFH3XLUkwRbZvVCV5QAfgy0H2EsACplniie2IFrzV9aO9EaVePBC3OMyCEPAVEJP
g7rPRAxOsf7Rqwauxat+p3Va2hfdT5GfeYbP1Poln0RRBWRgzgj2UVpUxv9iiiJbp1TbgO4wzrxV
uMpr+oxgOr+vnfCfQ0ZHe9l1C3OSdbaybuWu6Trz5JUGdqLJqIcmed9b+YpA8z6S9yQD6+gjZh0L
+dS0hMB4IF4nfozciocTm/CkoQBBUb2dYApzgwq6UStIPxFr67nY09g4+nJFzfQ77c4AozTqzuUt
eMG95Ltq7/x4XL+l7mnt+h2k8p7X+ZR5J6vmJFNT0MjqD/uiOmFOh/nG9KkuEFq/3MNZEsHavUv0
EO+uvBuHKhQARFr/ufPEG4jTVRlbews+yZzMk5f5k6quO26HOmPJdfzZHo3fqDA88ZhhEr2+R2K7
63zBU8LEX8cOBjUA2h5wCHrBlMB3EcWq8Hcw7tvpjTzACJuY9n1Vkg7b0ZzUIH6ohkhfiFQedq6D
fWYtK88bYJXiA+keXf0rEZf2KsOSpoeR3wNXIT3y5INRq1htwBzKYRh+ae9yBssaakQFiSFM3PnU
c/HppQjj60rfdo+RAvMDKXHA4xE25IBvJOZtg96KgvoIXnLgppPDlPcpZGZmxO4uP7tt1LTRvy5B
N7WzpFtFi3UNJrt/utxPbbpZFrxPvKWPhrk3anl/mIsNzyBvxPdItnZjlgAoffi0fvfUKlmYzzwz
ZKtzkiHDsqNzUUAKFb0vKVzhZQUs4UQ8o2d7VJm9D1ziWX8ieAYfo/8I6ACoqK7NXm2KGEVqNoSx
5mO71ZK3l7k5r3rKSQX5KAe5DHoOpgdeiZU5rJTRHfgWYzXkatcNHxHHPFVEyHkrfzXxp66dPUFM
qB4aGMY4+iKCPq8g0HIoN/Pv7sMxjoj2Nlb7n6fJ3VnN0h9ya/x6zEj08Zlwx8NjMLNRxO2UmGNt
nuimQtisB3MHpiJM145zdN1CvWQS5lW2svOKxiUwlQPqnyzQ0Hgjw4P91cMRNX31XpirsipKBn5q
uK30oVgOrrHDIeu83yK2QYlbzOcickC94uuqzqrwDhI45no28FStosqCzCSc+XMEv7+8SUGnZsSx
8OwU3oylYy8WGpOgK8EBaPzMb5qQuwSu4amjJtU2EYaJSGucA3TTqVqJr8uQFcj9QrBTstcsVwPj
6RZcIHCr3l5l4vWf8MFqSb51T3rcFiNlzh9VxSt888U3h1+DqXeAZ1lBUHaHZwAyQucJdTM+uDnZ
oYOIzFmD+dl2p1v2RSEp4Y1vUjMXiDoBZ/M2qKaS5MqEpd5vNvIgSXTsw9LKKBA/sx/KkrKYPX1R
ATaLAtxtSjH0GGSZUCEs/0CbbnLbIodIyRXHT25cDIJ0MpnI5CmKFJ3Q5s0wCm+Fi8Ntz5q9tU+r
GB/GalAqXb4Psl3+XlCYXYY/r1ybaq/rvITSN1S32ORsvM+ucP0x+u/5YpEmj1k5JfFVJL6xvpI0
oyU6f+A+hc3YD+A+S24KQ1/KKGa6hUH/1PGnp6cedGuTpcqQh1dmMNHu2W35hCHyf47Fkk20GvKn
4HD2tN85Y73ueJ26YLJNTq4kgitqLNnR/GxnhFrKC0h3ESolOoNJmVx6la3c9cu812s0CegsGuJD
wrnE1vcVAROIFNoy+ffW5sjJLptTzg4HPl0oOWtL1bHy51FVBkWB4li5D9eQca47RaS77rmGu6jT
/FVkXhpXMfnovM9OR1Hg8zrfVAMSIVnW4/yik4GSYJH7bu/yZnPEeokJHvY9os4AV55vr8aOeAod
26FR3HIEYVSrdmefIR7DPcRX+LcemUja12htFFmgCJISuNxrR8xRc/NMK6GOi1t5anBekw2DeZiq
UgMj3J7uojPGYH1uY0fqoYAI9Yng/SrgI+ykxmVNrMk322+NocP47HsmDzCchaJckCrkCNSssSDC
hQsFty1tSFUkECOXKejrHVq0S5GXDdprc62NiBB+LUpOHKsfIzDrow/M9Rh1wdWeDwO+E7508HfD
kbyCXZiB2/O7Lk41s6imZuIO0LmF1olUoFzZKauLTll6u49sO5c7tvY8vgv3XjvyFyjz2AjqKV87
xlgcw4FtQdV25U2bvMy3VslmYTdDl71Hy1xrVitAdehE949L00eRirYCaMHXvpiothb5VKftngOC
7gUtWkXjsMerwabWgtXC7cgkOk2Cfl/N8nWsrZ0mVEBJI66fb0axv4h1gip/lxunEYPXkN2AOhCo
xzU2yqDIbbuRRprPZL8fK0Mhb++CC1s4KM083YLscuAnQnVbnwNAp2xxVEQSi3gzBBk68b4uMWEd
cowp6IxoDfUrjiDeSvMCnXGTB9GsR6gARUo2KfPAHmY44VUlZufGapXyLw7bxQE8cUibqCRCVLDK
UaQlwi5Ce97ZMSMJ58CLWzI5HfSQc4eO7BzlbsZGPAlrIyvVI5n5JB7z/Uj3QYJc2Utj5D7cSzWU
zsKo2uHMZ5n7vwyMzilBxnT25Cx/80lgglZ4S9xenEQtJSYtDuFrbzGm9SW9S6w7gkPn56d3uhH0
9X+aBhyEJXeZjCxktS44vNuqWzO3UjPgRO85eAQlBg5Kru4vmSJRciXb/XeAGp0TdIqwDd36VAfa
R/KRUJKoF94mt9FkoaiwCVzx2eDaWQoQ1tQrcEEi3YNs7ypqhWaBNB1nc4XbNOf1Ekiz4JRQ9sJE
weIPMJgUOzz1/VQeJVjX1w2l+q14lYK/yo1A+cxV4E7WO61hY3Cf9306LvaOVZKqZZD9FHMCUfgU
hEubrzyPjM//ijTFiRFMoKzrMMNulBMbPV4VLNL4bLgAJQ+A3l8zLjR/TyR0FId6jZTgo1MCz3Iu
Z8lSiG8dlJPXdZ63WIzgEwbi4roAqkpoqf3n73dmES2S9tFDqULXt47XO+0r+VUyRz2MS/WxB0FY
QAbFOh21Lk9ni13qsUdimltMOhsfck5WDK65E8qD637SZHerZQuY3Ioenx62UI/VoZPFlCgroydY
EaTdqknIG17oDHwC6IUl6qs48NhFaMyOqheAQVHi0RodDw6+eVtEFDVich6vVWZyh6cTtuUw/S14
buhefrOyFkjoN04coxQCqicGCsiJPmnEzq1f3eH83+wNp1m+1fqYO9s6ECXhC1TOdDuKMs+Gh04k
Lz54PW9enr5PmJVgXreqZVOQpjoWg2ahHKvyjrNwQ8dGAyLKqGwi1JymFuUd6ai4LFmyCuwW4KqO
lZzlMkvNN+Hg4TlS56tiheK8itTx9KcJQUrdseQeHHWd9m5Xw3zU6ePoLgdO5PxBMsJ37QsRT2EW
K6M1FtAtc/2Kwz9DaXCbChgG8aKpXF3dGyKL7WZeOxWGLrfMTj7WLBV2NZ+DzMpsMUxwCe2amr/1
+rl8rBqUyduWayAmL8YwjAhFi/T0a5L8+rg5gO7o5jNwp93sWMTbKAcnY+CuGcjbQro5XlxXvBet
zG3gvcyEpyiWzkZKt2AfNFboyAKMe41nLbj45WMeSAN1CN8/xjC3RNYiD+6Hfbk2Lab38B7Jfk9V
HlQ+QXSeC4NBFMgwRotiT25iwBFc5yd7wlJ/L0cL+MNx3sYHqdAVLiZV3OxqXJEkV/w0ifO44dst
WPr1EXERqn0wecP/uzFgdUz/cf9N5KRYDCP4kmMlZcCJ/2Gx64IRqZBA8qBRFsQOtXedVClCxGOZ
FpwB0PZ+thTeavv6rq1jjPoqKEptw89m4htgKQeRLFZ4NkDJSZM9M9eFynl6AUMNHAKKdearVEor
/jsMeEWca51PMFtarHyBOwOhJmB0yvrgtyXyLvXUslx50cMdN6m8JRoEjHnElV/JNzcXDcr7mud8
RWPzLF9zWTgf5ZHMjso+3JPeiGGdn/4GI8MocivXrrh2jR5IyDJ9B/IfmUOMqKSFbK9l7C2cPeVX
gg7FG6gW6zFPZK4N5xrr5v+Ww61RHVufriH/+A447zfiTzkBlo/mnUAhvQinuDhJtv+IOes/VzAf
Efr6njjJPBuedVF5CHtCxsYTsFfjPREBsWkCRZpw7f7YMqYqLALgSX1L5ecCFqQX01R+KrH2AkoB
HRIp/50mknEBFtUofyvC4mcXSG5SxOyuqq2uOwwOfcMptIJ5MRE9HyhqEPxB5FuNlvm7bpZoJT3Z
e1V6OgaLsm+9O4Ha05gS9nUZYcQ32vDxtEVY8Qb2zGvXsE7ONWczd9zS6zJO3fyZ2HnZ98uDLAlb
fPCnZJnkAQPw8RrQS8J/BJXmboA3KjOB1ruSVst9xmqFZPOnyci6uvqFCHuVmPouhVL4mFbqFsF0
oZfMGhAC+YWSNOZ3gIYnKXxfGYj/mjcAOUk7524jMa26/2gF1RA81nJvOdWgPAus2lj4N0MGRh9D
WfOh/WAx7H9+D9icc+t7Yaf8H0r7s//Ax1Xu1duePSCp342SNWkq7kgZaeRGu22dY3YTIqfxkPsM
ZXQBtxPoNBtdrxP/IIbQxKXsHbuID01AQVIilQiy/AMV8U8FRsjbmAVN3Wa+PDrdERsyTAycWPR7
zIyOvVd5XxtHH4BeYHrlpqWALCmSHowinXXWtstczRBRX9OeAk3FqIimna5GH3DkIsMlnLD8SUbH
g56JehjyxoYib3zuD2kANtbYKMe0bEVIj3siidmgLfPyqXQgqVdGofK4Zq6ngyXnes7Jb5lKP5UM
3FrRbW4r1abn/cItZuMAFWpdUnXNv8BrUG6SXTH4eYtpF1QboPvR20bneTXfqi5FY87BQKZgCdQY
J1upwH4RUT3gar2DOZjSl+yDhs2JVoAZyl0W+9VbQwOzF8LG5x85iX/bNZM0un64D7KMX3rFX6JE
qrHnvmMSOdalNKYkyUGBC3ai8wLLSPxq7gmrJw6l0Ju6TuxexSPBxm3QPJFMdLcx5ptw7co8YRnw
Z2hVE3Fa9wjAX4PlVW6JW1y1AsyESFzr8k2XQ0m367UPkzBjIzJwiLli6Lc3qolirTaBW4tK+3dI
J5BSggOXB0Qyq7cgTnVKiWRAPBOoYuBxhU+haNVZVzzr+e7bQtAJ66ZcFOPTmpUCyIqgCDiQr+5r
97WypwuyUqtn38QVyvB5VNaC7ASCv5ua55Mgoj8qc/v8pr+sLWG9mZoywRSE/PEIY7ISj7CJ42z9
Vhmtl+qE4jaHHurmjRTvF9P1dT0cZzlYSG+yJHL9Fk9x47DJZKGvLsoWT9hNfQ9YvkCTYdE7slmq
cbFVsLJZeEMxS6/RgAAZ5hK4OV+7DhTX35cGoXExT6A+M8gLqHomboZIWD9f8UhDaS2rGBl3MtiP
aBi8tb2s2oJCqBl0//InoW2VZPZML8kXZqhrqGuutIQLLVkMl8M1fez74Iui2hqb/jSUmkipgh6y
NthLe/0nTqA34b6OmxSk5NrkLAMxlNNWOen6LQ9JWfLKck4SSJaQaP6lXM3SiDeQFvvWXPG1XyT8
LsdUREJ/Hf476UN6/KtMVWG7xOpiLUCVS1LLoECWynfouDB9VzaPt44qbjvFVg4J3U+3K7lq1z3m
eu4tz48rSZYcw8oAx/eWnMZBFFYTF4wIHVYEgzEVKS9v8CuzekbwUuYq7cdEA8/uMb7e+MCPS0x7
YN4NcVRGY0kXKfUZmHyxozbS0IlGY8j/0wplrfRhDhvkXAtazELpGL1fbSzALA5+Jamz5H4ztn7z
nzoRWDUFU0GohXXDCmrb7Zd4K2zlMvjLabx3uXxZ6DowlZ9vQoaBXaHSK1fKNLufTQn48N+rHPUQ
XbupjRmqeQHITa1AUDMjHkVSYVCgCNm0Pswqca1MPvxXKOvCt3j/unfY0UeR7rf1TyfwBu8Z7edG
xwhRK3D6WRvM9jzOCxMkjssy1IWIsP4Q19li7Vcae7UQuMpIisgXGaiYvx5flmFnrgGvCCIL4Uu3
bFMSjj9la2SDjr7NPDJ0DUaWV5pLGiGGXSYRmIp2eX7oVnYUWGdrjSe5vpGK/4GgUvm/VrTCIxot
IRMc6QZE1+7CDCZabyiFEr1ButOyRhFRMPveN9WgpEFvPCitiJRN5bCiL3GJnn99+W6ZOh3TWbel
li1WC+Ekgw+QJjNuB/ET9qsjyYh3/ALgEAsMU7gB0Qk7s6nTJfi+Nrw/Yoa0hfCspixNyN/YpN1r
2DXcOhpLC/VJm/fFeqeHRg1OvrjCGNEhPfe659/UAl0NJ8ajsK/3FhNjEXEa78ytxM/Lxb/aizX5
bFaZrpffWxWB/h0W1XqE2F8eM+JDU1KX4mHDqPi6OpYFeosG82h+dFeBQJuEnP0PSpcu46kQJmU/
G7w8Jvu73AJbsS4t/EoJQS7vS+kw7ItgqoiY2cVGuHtP3oumh9d3iGvTd51knozg1F13Mir17Wrq
fGpfhm3+YhxErBwU3VLfUG/R62jnCI7VKli/8rSUr+fwl0iVD+E2vy1w3BYHKbiwnGJQRXKyQyMD
t7XTAEs0moXoKrOgo1yOCdOn6z55AiaZmH1iqpwwi6HK2hOM8gGdedFacVZ7zYDTy2B0wTD7ujEA
NtsCZcBHrlp6fGuXlAZqRFBlb3uokeQsLSfmMF7RbnCkAwdkPtyUPHyOiCI785YzRmsTySY31dYf
b7Wb/NjKstADFEZ/CuN5kEDa5/jtsDLwDdWR5YtmSkRyD6cV6B2ScabaRf98Q06IZ/ILhGLaQEwj
E+sTujDvzx/2FzFmPyJU+OySp5jjVUtcIJwkklWL7JV5LnQIWOQvoCk2iC5xlPLvt3X1kCFRGQkM
xVRz7FlS8ZheeGmjN7Zf8UDDPL+VllptvEF3ikl9JR9x/2wVH84P0Zpln87jBKAmGOrhfsFU9zUk
lWU9gWmGUtBjGvBZseaq6GcpFGAdd5owfjtmOVi2sQp66TusanQzNVut46NnphiSS3GBim2fk5ib
DdHhNUJ+Q2GfyPO/MGL4z9wYMhV16OpuNxKkkwumIZMnyAeddSe4gfTeTPvgzv9HFGBbAkYyitWV
IUSE56oMpzI0Qw2BnCeLKCnHGfKCWao4b6+hIOXoAzuRkCKhOYiCDTr0ZxFMMAKqPMP0fuAK7iS9
TpobhnzxG6xzGalQtJ5HtcSXI9d24GluEsO5Q5EKDeaUOpnnSU/iI1TzyNQvrXFIne+h3FQNMHGB
E/LvMqPJOcc24dFwHerQRVDHzl6iF1A2n+rSyRC1kPWMZf4MKcW+qKhc83JDxlJuC3ODQF6kjEc8
jOEZyXmEYNziFcr+FU5oJoRtsZiRPFGL1OI9XW2nhLh1Q9QnhY8Mozg1poLpUBonOr42EZgx8aI1
rBFS6FfKRz6dP4habUvn5RT9ude4o+RZK802m1Qk+vNJqEzwGxBcIPIu2J3svHxaE6r73xwqqJOj
LnshDz8luyPCZPO+SiaYtsC1CI2Jrn9xO4CO5PunHR+6JhRFXCz0VpUBrBN0OeW4sNf3VXeZiH7k
nX8MJbICyuozyLnR5MUypGcEE1gkh2PXom4lfbRJ23TQwhfLjMTAZwA9ScTy7RjNx2/W+G4ydAs0
HVmbSDatdSMacxHwt/0JAcG1TAw08NI9MtQkwpAj328eg6U08ob90sN9P8FmLBNG7Ksa54JRf3RU
GJKpj3qEIQurhavE7LY/oNrRXnY6+pNZceMXFpYdX6FB2/Xw1edZ6peVVesbwhIE8KCzVxFs7uFY
0vO1e1dTSjnaY3ogMHE+MyCsSKGP9lPUyTbcdoplXM+mGAJoo+rorTFvZkU1PfyI769aQXGTDn3j
pIEjusovUZmqxKI2+LzSvUX6cgQdFpNdFPC9alPJONSxEjjkGClKdJe38IT4IU06t3QMdimBSSWl
xwg4OwJsb/q9Id1DP3os2eWFSOuP8IC8k0Yxw25InRWbharcNLY+ZIRKahuLO4ZmihjT2WmC0Y3a
GEm0+pgYlPiNkx0gaWMfW2our1m/CNqElgEdU5u2VXvhBVFN8yMQKM4COj+VaRXmPJH3UePqiMCZ
H38Arbni+xUDIlizFPiYZoPuR2sg1gY5TJ3TgthSLdbPp8NHx3BBES9Pio7MwnanpoWkZqNeEWYv
AfNmgkl7pZLS2lLZcjK8cFyVYV2euCyOMEXfzkuOhmMqFayHqq5yYeyc1Xr/XUESIILdD7P8+4oe
LllXW9a0usg4ryt2PuU8AdmPUbnanTLvoluzq/B3Y6XbxMWBaIxp6OeURId1HAnOwjktUzInB7M5
cMwezY0LmBRmhCS2ENm/dAZ08/ciuO8GuN9DtIoAZRWFXxVbcFl6TrSRk9ptLbDwbhs7Ju4I0jEW
o5gF1RbTli2f1H8r23hK8eGFJuZ673lqKmBK1j66D7G1nIhilTO+flfM8jZUXN8ulYNZQZNuaAd0
2tX8SAy3rFEtTf2TGGuWH1xXTf5fmL3uwZKDqHh1ln2xoJMM8mDp+gY0kC/CKveTRH5hC2zlhpKE
aUDnQLl0nWmps/dCftT4WAKGeLnaRf9az68wHy+HBKmAHc/bTOxxm61VP7IfWpXpnMabhZm8y0gR
zz/gCduJLjte29ca79qftZECMJG2R66PsyZxy+um2RnTsqOdlW+JB47JccuHidxxMuNVoRZSWY5b
ZGm62ZCjnU5mcC8mrnggBskZYAOiGCQ6nUN1XDsFXTEWx09QL1AMSLujJgD1QL+P2jDs6o3WvlDj
P8Xw+rvp0u/TQrkzB51Q++n1DXVe/KsGoerTvrm2817ofABV/X50YA0iXceLcRYT1bo2rCIbA9e0
I1gi3W8N4BoJrH95XycJ96JoCZCgay1ooXxweSKcsr3s59BC8TdE/aR+9cfEcCTiRs8T+Qc37X8N
/T2YXGXwZmxihnPehNHpy57j99ZAmSLk2NE44SpNLAVcJki8HTRISYN4KAuLHDiHIQhAhv7hNA8M
+3iJMz6uw/75aIm9UWigfRxBiaWbuuz7ngAU/JdevO41K2XvNUbD313tpXpn6Q+b5Km9wvZDamtk
kNalUm7o+Igzm9ogE/29p75XCBjqizOInAcdCwdID/Sm7KPYJMhbFFUuK6qjobsen3i6lPIG6ih5
DJ7M/RENCXRfBFShjzNf0I4HowezgDLNJHRmgbCuJTYM6oK+PjzHrHyJ1QLraq1Mthe61siM5BwE
YvD8r9d3SzT9nDU3drWZn5yYnMkT9tR5/34C3GZx9G/8ctFSdfKzfyRi8UTHNzXKu0/u6ZcbJI3G
Uoa8wHZ3/I3CG3stMLX/0lmyBifFZbvKMBL6KuG5xx2F488L++NuuES8k1ry07JxE2jSfFcdCkD0
BMlzG3/oc0TIGe6ZeOCWo+S4X9YSAEKsDr8Z1lWOLERRuc0Jb1WxS0zwE/EN69+T0JWuQErPZu3g
FKVbIofCDmIlfG960rl3MyM6l7N+R+ZtxckAV91LYXAZqotVIjNiMvngc8T26ws4KOuXYH3bP7k/
GM4UH1N2Wr+Na2gsacow2f5S3o4xM4ulOl5iOmPLOJGpJYbY/HnJpqL2+CwjSj+YxcHzOS4FMXPl
QQ5QvOK99+xg6wnwjBxAcWdYcrBmfkY5R0OXk55zAk4DIKVbaS7nRgDZtIsawOCCRwmVQ4JZn32r
IzgtpKS6Ls1h2trDPeAodxr18BnTHu/VSQg9R2aVGzon2slplRtdjMLbt93IrMJovM89I5fTZOX4
1vkl8TEtFZg9VRkE2o+t/ri71rNvkFQ9YcKqP7vwS7so2P55j3AUBZ2YUMhhMn4ida+ye3QhJPR4
g2xvcOtMlXmxTKsXmR8S5H41kd1IWwj917gmoi3c/vjXKhPtBQJl/TtMV9TAr2EYVVeCHprwTyEQ
x2yjlvsyvzPpw4y71kZaZVG6x7/4HfYnFjlTKv8fgjojxOEmsRi2iVGs2BaJCK24NrUyxBPgu3tk
0LlM+/uESi7Z4X/mdhwtNgP6E9d8xABuc8HhKuEUgu3vpdpG/KnJHbPN2YSiF/viU+WkYFoHhVE4
lGkjjpZR/tgBpqungNjZUdBw1JFCSHlDW9xvDTpYUZkJL4OrjrV3sOEqBPCT3D5K9HFOAxz2w/K9
AzwsIEiBQWpyHFbiA9qiDmkWG92HaAMZyIjtjqcOkXnd8SE/AvHlmjivbaRBg1P9q2uvJ503srim
QZmbWulquNOyFYaWePu2m9D3VZi/gl9/60vT0q+g2lbOzL4t3mdbYXHF50OUCB1KVxq/rAoDU/Pm
m8zvdoHyaxyublJAkXzRCIOix/gPhIR5dzVnUQdlXK6RTA1pAoeIXExIHR0udQT3oGyWcwlpa/W2
Ubwh42YXjixm/SDoXouqqHmGCp7aY0yLjKqarOGrklxVShQ9HZ4dDbbukU6g3HwZ9uCYbGngBrdo
V9CEhqA75Pbm5+PmNtDmCSetgEX+ptrqyQzuTEe8Kh983zqTeKF+FR0zAMrBm4Ipn8k1EdtajYcA
C82S8qArBmhRr93G7zGn8ZBX9CQXzQV6NDRQKkWBt7uuKDKy+O0IIAVvKFJO73Y7ldl1JhQ2WbEZ
ri5qKuHO/DCYlHG6+hOP4zD1fgPI9Q807bCbY9q5XDT5XFj9QRUiekpaC3HhmMdpezAJLkLAwvtt
ALa9qOAg/yGfrZZHKAaQAdH9/3FnNXJ2exfLcGTPzbR3v/PCxiPs8Fpym0bODfXNPhSEoAsjnCOa
vMQMjepYujqipb4lPF4cMNSGcaGPZ18ODJTTZtQJK6dbHxmgt9Ig6iHns4d70RkZXFLHxXTmBX9Y
VWZZB1HQomWpzDaTYldQGJvCTQkUsAhqoIK/zT7b8+HwhyUwmPDXUjPghh2gXRH5i9VTLqTe35xY
sUOHBMzn9r0URel2kLzQikvbMMfpSh0//HGZoRBa7wOGkxwIPEaO8RD2qznI8UKqLEv/E04ZLmEO
CqzYCFsWv6GOhL/X0dwl9brkPyrgeiBkpY8GPc0vf62EHzkf+d23dPhsjN7nhAy7CjA7DQZGMZsp
S//6Yme6HobLAUGOd4Me5qM9VYOiw/cXb8FlJVl72WSsfDVpC3KBM9qCCdZkULLszAQcGG8tni8D
N/15QYgAouxushvXisvn2swU8UHdDaVvVDRd+lMi+ie19BwkbWXCKgh0gS+IOP8p0K7dKTP5JGCr
IesjIDwKh8vnoQ81WNdDLEYG9QhMArJv6LXq58dGuB2fpICqFJmxft0tS6cQtxAbBFcHdgnSPpue
yzFibZogyFtbvcSU3VwzIWgVzV8qcGP9+D0IloLQos07DjT1QSrBPQ4AMMNmvkbkDj6ScsVa5sBW
a2XBcqOYGR3QFGSVDePtOx8MtqXkUAqW2IDQaFkqsxWVhng0fhrtmgdXXrhSMMqjcoMEe9ULWMUK
RX3G+QsGB/yjCqDPggjTzOaQ8fUFzdipzDbMi4EAU5vZRcZlxxa1JNgbYRj5tqp/pY8qTqCTOQWI
tdOjJ9+SwbXq1wGqFZIiCRJwenJj6KqHCUrpQ9GhGHMvt5i8+eD+HQrnkZjjRPEXByIgy7xPOFlq
NFU4oTmwY9aPGaSollT1c5cbPUdtfTWHp7sxGbNhUpeUbl0VTz/MyohvBbbmWJ3k9WH38YkMDH4x
+GV548JO+dmxtHDpgpt09vv5OKeXOwDag0uVIMmidwB2cvwGKIP00PtBY/Mgm4np7VQzqHJB1Rwj
vHMpFQ0jly4+syst5VntrzXFxTkyAiqfqngNNmCNhFfmWH2o/lKG3Aik0+WU9QBxtKCVtqsupyq6
5rPlPJi4/kaQ503Bnd+WAkp2EDcZcOBtsVb0qBqzzDK5uaPk6XFMZLkRhHgerpt1sDnX7vMcTJ0x
pceJiZptsNF6cxmNqeCEzvXFzUZFByn21y/OxoNZny30HfC7jzcf71IxNTkHBT/aNImigDdrAtPd
xq0qaA0pdztBXt+tZ4GfxL4KtJPlcSJIOqBOsBW+wFR7ontPGewz+U3uE8G3echm+0ucvCJBJkFd
0Q5JG7Ng9kGNt+ORBwSlGvVnJET3xKaHkkVuFeSuGzJFsDTmhb/vCvj0dmdm3u/zeQt8HEFHRx4c
5eva/risXidWdktu0u6lDtp5iX1ekp0YQGSV/vPIHFWAGkrUSfJyWwvFpp4LQdU+M6nMqS+9PZw4
QUvReQbAooH30aOhRRYilJLH8dHuF/rU3TqtKEwgFb/GyoCtTPxuvxp6iOGMTjyDBAf8BHAn7dAM
4CnRGxlDNXLz+fXEIH3lpGbDDXoEU66nmma+OZEt+17pta/h3UhjMwajkHA+8+sFM7wRwU4Uiinz
yzNnTMmSu64SBYCipkFZm3GY8/CyfgY5R/2Tl4TeB+D7PCdW7lNxGmLRGoz2FE8PXbCHgMwq+bJJ
3cDBmCeKAf9RAWmUdxXBUP+h3fpn3UQlqmKw4hjPKbl3KpqLqA9zcLWsysIDPb/AMCgxsMleQ8bO
abjevgpfwyzXKn1DUal/IPiLjNyQcBeRPdU5YOmzm+EyLPW8hGzBWv1GJAdg0G4rzP3C3UUuFkQs
YvfJ38uHjzrvAaFF1QwPvE+A8Tn/ayU2bYJdcrYJs4ym/UpsWGIvU1d+tI9skM+vm6b3lDiBOvf4
VIIUrdUtbBXaFGr6X40+numBttlorqfm+R3DH80cyYxPAzY9Uz1tezjB2tRdx/p7uF2jDFPitdIV
bRv1be1/mjxNMSp9cHfkgQrj/NexRDNhBVqmlRd/tgIxzUrHMI4p87/4jJpsgsgdy20MG9VG9b8g
inFfaMK+1GnL+iAd7OPtFWCEh9qEd60weMqDuzYYJyoBfe+3yvhVYdltm1MibTFO+B/8T3Obdfs3
I8UTLbU1HbDmXKZwieLTVidq4W4Q69FYsfEDXKJBKvrAx72oJREzvQmGiinI4y/5LJsWX25ZZbeb
uOtCCPkPE/wTAyeOa+EBg7zPErHpzGLHcATDa/ZntH34aciZNIU+wTL4qqjdI83qtL06iOB9Vvnq
loGPiHbVcgxY8yoJVyDH9ZKYlJSDvyb9awhOePMYAif4aUaeiH8j60JSTQRqhdBMV80CceBq2dsy
r5V+Y2qry1dvRFlfwBGH5bioZ8McuJpVMdOhPs/ZtTBkvTq6KTyEcQ1sfUI7mbYb0p8aJrUXFtj/
vOGHS/pLv3c0IVrbqgAJu63xGw8oQoIAn3v7C2DPVd5Jon6PceRDO0TxPPVKVTsxTDbApX5baYYS
mrc6Jz0YcZF970o2BcLBOrFc9fyiEGzO8hxdhs3MrtMS8nKEBbBvFx4fRFcMa/COSOPkTNx82zGj
UzWqmNC8j/ogngpNOW17XxEn5BVsrqSNOViqT4Vs7rhjewXPSy28QdiX0K1vR16UtEgN/LfGPRND
DGzaGLzQP2FkAWD8F3uBIXoIe8RzEuCZlj8P7pCZUihjKcGMvrGMMxqlnNR7QE5vMFJbmiocPiGA
r8mpPlYY+2K1tNbgllO7cMoj2hPj8OKwXrAwUoQhU41ELV0w5R0zylimmcNpizh2riVDTOf0CxBZ
7jHc347p0Zdn5sfnvKSYDsTuTmIAwfbtc77Mxkmco/Wu/f6LzRZ9GW1t6OGXah7WVWlWBVfvGH10
8jOY0DzzJeuvFsPrwR2SE8zGyyJIRTM3naymBiLjBQVTXaPikGcYFUVk9z6a1/2PIAdwJz27IrHL
PjMcHjgOfnS0Q5Co6yVi7OvBaaZWmd59y1jd5QI741CRxVsrTgr1RUAXiYcRZ+1z/EOSso7XFrld
ieY330t/7rER+vNeiSR6qqK5H5ap9gK4VGnClVptVlYrKOxYejXEUFVad75ecGvae5QQaYhO1ucD
/RT/fZciSJmb55m+JRo9CO+ivT/LDz40j9P6Uy9JEKUnVFWWqb7M+k+r657+FD6FONLlCq2nJWIC
ZeUeGwYTgl+b5XOvZ7g4Oy957ySuyDWXBrRMuv0K2Fbh3Teooro6Tzc38REVejaVRXBKl7bAr7+U
y4d9jqH9WkR60JS9w2O4Ycya/q8Jxk7DU2rteAiunXa6bqF9v2tF7BSmrZJSf9a4RCYiKgLEj6GS
R2GSMnFYCsSqoHfCubrxcekQOVxA0HPODQ+NTB+BQrpA4ayP72jueNzz1MxfdHqNQ9ry9Wvovr9M
5yKTPtJOA5Dm0azGldVIJrnKAMPBnPuf2bPP6EcnuL+MyKjP8rKvWbszglO5k8zj/NCj3GMWaw3I
PeobKJvv4hxHxX6yNuNXwCggd263cu9N365Y9b8xphQbVU7An0xZYcfEYRMF145idA9zswzIip5k
SGt2mALFQmByHub7y+rsxzt8YcxqYsg2kyMvYq4j1iNsLqHW6FEBMEIVoThTFDzipKypczF4Cnzn
BXVlMk59HjcNnOE2VJ6Np3xIFht/LkR3hHqwo8kMn73c076Z3mYlLGWgwuq63vUuax/u5V/JoeGT
hRWEtCbAPlNjxGx8BY53vY9kSeW6zuZdjK3F4rB+KWWyhnWBu0rCIcE95DPOWzyozArxvTBUBPOX
tzAVBhasO+RARtUbjsKKFFsAzCtNvhronmSP1mfu2UHybXXg8JRhOTSzwmo5xM4lIlWQ8BCaPiF7
nv4W6486pt55bbOMkH1P3DySeZPCzxsndnnK2RNjbsivgr8vS3FglEO8SJ8WLYn/wfTUKeyzUTXx
xDZ+m/IKM2xyMZgdPNFoFYHya89DxsxHprrOJpngT0LfQqkPsPgaqBITH37EXLbQQM9h7LbN7mF9
McILCiPXgmKnFUZNJ1WZCm/pj3jiPH9BFi0+GqUmIFXDBvc5YuFH+rFeFzNQiobbdb+eSIsjDTMI
uchnIKWspmPJvywbaCddZeyI6U0KvgX7zlxnM4mpAHKX2Oz/5971aGdfXd27L6rR9GkBDgvss1fb
B4vjFWCjaUuSpQzbSdA0WJBplspLQ3g4UjkS/uL73+uKGjzN19dNDeCMo/0rfquJiCxLSVy/52gq
UwIs0bE1rb7N3vrGGT9jU6GpX/DbZjFyQ+SSEr9j/SyBKCiOgQzDlseqFkbtgaBJTrzPF++XbRkW
CqPHHdI002VGIULVwXRD6r0gaBiQJR6tahETv6UvyL1eFkWDPem1cNIXi3EMX7ZyQwF0yKMERTk6
a8mQJlD6aNKU6efPrRLbvDWz199rswC+S0mQzOlNDCdHGWdf+DT7UsyPrrt/fUfOaLHNXNEtnN2o
2X4KtsbsRtwqfv9mgiKh1+Msmk4u6rGOMMNUFrABUrG0EbmifnlgZheW8OgtD02Yh43P3iVcorT4
vj87JbJfeHCII56566nAfzUtfdYGYCdUvP2ZUgIcl/eA4xD+gbqbazKALkTnUO/18Tj5CWsO+SRh
Rsta08KfJHGnO1nqwvD76PzbW+FFkV0/ELTqc5ESrKNroEilPw64Qh+QIs/JK7/2r2kCqygRAj9q
M09fHgogBUP7S/7gFVonJZFoMEx58OB2n7U0pnBwhbITDG9iOYplFUcdkZG7NBeAXsr5RXADXdrw
l2o9yjP2VSJWOxLTAzsppdMvPMYvuKFQDXZhcQgM3RxFKmA6u4mR1Nr89begYbrdCKR/bCyoP0l0
PhANa2BrwlUPSIq10QsU3ZxxfpHzfGm6AgG4yIj1ZjOIh/Q2vmPc44WjoE5wlIoLnC7/Qp5nCqPx
mTqSQg9AOm5ylBuharDN6aqSlnH55Sa5fEhsTQxXR0YgyktJvIrO58lHz8j88ktm7md3hzhOaDv6
r7WA935TVYZ5Y5V7KRPxzT/FrcqbNE7SEGOBq6Fz0nGMcXSjX13DSBn7XCojFHpUjnbGKjLOaKcr
n9Csn8j2JtgDelNaqKHxQPS++jojVEAXLW9W8tB66h/h3/dTWX/LvjHIOudlkkoORV8fDmluwwF8
IURO6w59u4Qw8C/aBIzbB6pw14CNsh6vq495sqOElJS9rifaqDc7w66S+01cEgkb70tattZX237L
uaHcyOjW948qMVXfGq9Kk1LXi65xd16YDvabUYXr9a14NSFBrT5c6l1zzsdl17FpyDgdJrRIf36H
sNIaGM+fTcE/cNifleeWLyCHsnW+dRlEay36ewduebsd++WmqudpSdxgigs1/qezdX3aV7sTH0sG
yM/ADGYG9JDQC/2YqWo34/8F4rBfETzuSkcy2bBqRNxk6Wib8/UND/uBjcACBc/m8SrClgHx40b8
ZCWsVpx1Do6Uvy44zuvb5qWMYL56IUs1Ulme055865h15ecmqUYvnVzsg/QAMEwXtDe8xaJlSITh
Y7FPrhHbos2abSQZnD+XgzmtFjnX3pnevx+XNxmFh9HcSDtUpGhW2DTOum8+xkkNIO+NPoa3f3nk
8t9OnnrokhTW4Af0l2plYOyxzFqz1JZho+BQXHZwe3FE6uBBFg9mPCOf2psAZokCpBgzbfQztTE4
qb8wO8/HK3USnvAkjjeNwgITWrKAgaNIEasQfPWGMjw/v3CYsbJkERZK29gGJgzQkH0MoL73o9Yr
g7VizM4JYXH+PPFs7AzCPcb9n/yCw+lvalUYXL3yHXpEVO/A1IKSM/zuVwyLfNdzmJnu1muutsaD
mGEgWJTYI7AVxPP4Isfpk/vOewpWPn1PKnWIi32FasF7ssPZCs0JU5eVOxGXMENYigDlcWXl4z2P
Uk9uTfULPRCkKycvsmHfcmmJE6je/EE8keDLIs0QrXJhgb0b+PsTQDLPHzQZoYy9pjZuZtNWOync
06e7ydGueUcY3psE5akaVlI38MODT2Rt1FRlvb2Suo3Fzyk609AnQWrCYS+I5eTQNnb8zqCqHVXy
TwR9wD1GFmTKpoO/M2o7XwLGtG5RtG4k7K5uw/hty9HKQqG6CAACSUy+v44gfKAhbSNlJ0RN9nQO
1u187Ain5nO/4SGDNTL4vTuqa/NgaUtjwR0PTL+dJbT31PWVB22OdCrH3WzNBm1zcVOfBUe9euqv
zQrNKHXCiociOnNM978pi9wPcz65WnAGECYPiOEkdUh+RUaM2nwEn6Honv3+7B5q/Gaf2S6L5TBm
xha2ij5T+HaHsJq1goke/io8TJKLC+ZkA30vo1kY1E3UifdDZJoyLqyLawldpkXg93sHWP96jQdB
hX0TCMXqASJxlo83BA3wiHcB4l3HD6kkcxYo/N60casHEzQADBqOOZFGABs7XVsfFNpLF1uV+bCP
Vl9FGUPPotZTJWFPjEuXMA+CarvouCyuU4QC8CLuUFo4Q+pNwo4Zfy4Xa4c9zOyMnlqrlGrPsTC0
DOi5POIr7ibfK3VCT3y8B6/83bBVo9/5IWpSCm1AmnL9BLg5YV1Xjv7YQ/GkxfsLAFESAFNdrl9A
rQd5h8UmqoDwakN8g6o3pCeWywP4aMN1UaWyujmcJMV6RbSjNI9huTUeyn5+Yrt+2+nW2c9XL9Iv
aEmdwTV3BRKk4l/yzeLZyLupdK52tGBzE5XZMfvs4naFBAbD4HOza9vd9XHSwvQjz41ph2BWxXln
bDro0aVlRO8BomRCTqUqkojnonUTSdjm+JOU1LOwFdIxhRMmUejg1GkVyHYyJMOuCm50pjIHubDT
SMK6H6ca2TDN1Iz0TqOoHy3+eMnW9vs0rFnxgxnFlnrTyaxDCkpvJDk/PES7m1IbEVKGPAmOGo4F
l0ZZUWC292ccRvpyYZM36KOhpEIvQqEjlEKgRH07FVKi9zVJokKmY73lH8puxBDG01y7LtIqpKQ9
GPUoX6PkepYvDTH8SVri/2pnW72oq2FUNCnl265tv7KyJeX/9f+fGlFMC6h1b6G6UvoIt4V/hImY
F5xJ+yXRNOeJgUfbm5lKjbwqIdWu3ILjEsUL9e9GzKC/zNWAsrO5+4f3VxxWoeNNeX7XVSoGZcSA
bGZIj4FkgS+gXSdUamPvjB+bBS2ofIob3m8qIIccnplaCJL46D6KMrSe+ogKKYCxHDD3ryve1q7/
0QmeJcT/hKfSlKAaTrUXILl+MXKTYwqN+yk35DQU6Oi/diNYNNUPDgm08IyhHW7gcAuDk9JwK0WT
GV49TSIBQkRa9O5V2cZNjpubVy5HJJxVP31FvaYmAn7JCThfdSNPANoiSvfQecDrxTjUmak3s4bB
FanV4va7aeToXzCqR7yqJNTqn0G0AP/vKCFlxHZZo5yYwg0ulMVxS3uLac2iM1yQ20RncHCSiIZe
bgsVYeAtANjtLzvaSIXH9mDpL+0r5x3dLp5Opjxq6mpaGoWAHoA32J780wO8qUyf1clLq/Z2WDs6
KGjyg+OmGir9mdgIyh3JKXl5fUwhVOhbGDW9yOUMRj2J4tlcijLHhj69iNCoT8KmBbAMOrki1lBR
aTa6c7fCshhmdIJHWNuNImYgnX/2YI5tR/VZJFW8XhHIAu1vRS5TiCTi+cqx8Yt/joPUsdbCNCjr
FbaCMROD7Tr0VFn5Bs11gj25p7YRLh+GMnfPphfLoyG3XmdsRslwRDwPSO5oyVn6Vs0ICqS3Xr2Y
DWl/OPpCBk6i4poa6pwf5/0blSIWaQRSH4+AtxhS05WYF3PRlHQEsU2iWxy4HaoZKrWNaEfHb35W
DAsLMgkmk4NW03IZydviewHxVJN35r1zlqSTz8Bq0nuApfe2vMKG/EaqS8ukXk6bwY6Qur35cWOB
pmDQmW0KRoCwLDXT9OahrpNIqOSF0re7/HXQLNpQ/BuIVUUHseRjNvkQF13rANIx7kvUfDxDBHNy
4m+a9p6t4H2c1b4fpdqvXkmh3+gnd7hJFYJURzMh2ow3ODn2hTJeaO29AEthYXJAeWLFwZVFQb5G
qXGLtwHymDRNGDu8eiayFo82iAq80jOgSpiqs2p7/E92Mgw5vQ3qDpBnJCGUEo/4GyxsFgMsOYwB
E/Frez5ehvjY2ygSLaDppfZ1MrC75bzk2PwYCp+o1SDWGWFVwSPfCEtoi4aKjpl/FiKcNueXG8y0
58A/q16eSS2lE2ENTNe8WuQW8TmEG47anKzw0yuzbyv/mM0Xa6B7735VHzCCcKZ6AVX7i+0HL4A+
eRXtsKdbf9U1Jrr9ZnV6y74QyJAaJj3UgUC/+cSSMF7htlwMgoXTvbrNxl/eC6T5+QgKfiWpL22N
66Y4HvxdHqvIXcsp7X9tqI7fNaNst02O+IBgrZgkNK1jdEOpQTRptKPGUst0h7kmC3gua8Row4De
zyMmhxf/X0FlM8P0/qccnIIWl3EBx3QlvOz76SR/7grZVzy1s8ugVLtFGwwSvhsy9z55Ylmiyllb
oBhaTSFq38ENX/WtfHKvCOYyLravpBhP708KaNu7g9FZJGfbdGCb6oyPvi0eH7Mh/hOsR+Vu4ZOB
k2h6YzZLRL057e1dorN+oHh14oi0joYGK+Cn0ldaa1o+dIwcxTCRFZu69OaB6fw6GmhZUn9gaX8h
ooNXPpcLdr3vkuEKAnu5p5c53f2eezOu1EszYS519eSlGmSqtKG0Ce64Ih1K9zIwuRHG1++WZdjp
UFhrtK1rix/8prEhLlXWxeJud99cu2sZrDmcJOhbDQhVaCAvJ8oHWNNjUvN561/EGFD73vyy8Van
QKqxtF0lqS6yk9RZXJM2rdXp379rkba0rZiyj5zniVl+Gd0IaBlvtGoEXhaqvJTG4Mlcw7iYPPPu
GNhskmvMVWq2s+Jix9pE5+6nsiaCZMF1tsUDZi/gteDguy3W5F3N2UKubTsDSesQ8oJbmnhL8BuJ
o6+12KJuuXyyfSHowCd8gCZHotCG8H1MguTinVtHGbmREvab5CkPBIxGV7tvNvU37ZtesDhUfXbj
U15SlLvrMXvcnGAI+sh92cuwQXnWnaXrbJW8s4PFF5Mc6Nuj2HjvFAPIr01Nzl5+QdtOleHYrWOu
1nio8O/kQWb6Bkon7tMh+EqX7P2v65+23LYHC+mxoge071c+mLGk/2ygrYB2WEXBOZu127l82z8M
v44wEY+nY5fsOKcsY7C2nq/Rp2t/3E23VbD01G9wTcoIWebFvJJi3/ZnQdU2h9YySF7gQ1dD6L5p
4INktS8hxzsMiJlPcjlGTo+9JGxSok5aFDp8vVMJBK1tToN6GGugq6F77Fefy8YD0MIcgqw2Nh1T
YRiOt0nM5eH5z2oigXI+mFysN2vC9z07V+URCKI8E3skd6qamUeZkoiCTj16CBrf9Ea5Of8AKcoC
F4A3MpvyLi+REYXzeenSfoMI8NidsmyqfTj9mZ+lbZFoSeyFJkuSsbhsw6ku8p0zB/PHeaWKNXUe
Y/jBeh/Xw+szadaB/BawuJ2bOXI6uuNJsN/+fZriu5edHlFkh21bQCxSjYbE/WSJHG6bb9NqUvCT
iGCJOybda2gTyjJWrzEQmBF4Iou6BHA+uPupF82RJ/B6Y9fyZU3trepVvOYDR2zFdUhZTXiCg8+I
0Lv8eGjG1Csj1fkGYw87ZdZwH6jsk9jun5WVAx4qFiuCOsgMDcMTI7Km4EtpVR9VGacP9sHZIW5s
K1KjexUnlWM32X/x7bOiK/aYvz1kJB2o2cE6jLn99J0qekhteSzFGegtObZPsvhw6aW1GV94yVDy
o+bzGPbD4iG8yimHEDqSYJfuDrUgwP+EMsOaWq8fFl/Xpea8z/5Wew6voIbHFkEWgh7II7dguYtW
3Ta+eM3p/nOxhQL/hbcoct6LPRHdfdPF1NXFU4TgUvHPSlpnvmRR1URaPLYrbnGdAfPd3T9tdwgL
RmuKk1qm/5miPcaGHinud4/yBLEQzLPr6rGCtzYSXOk0igXW9rKbvG2/587I9/P340jMsq0JljQP
4qOuKB0g7Z6Q3wfXubFfPiYYU0ReWfTaEdyd/zM8Tfot3fUP3CL+E1Wikz1fzZwISH/9n6LKDR/M
2s44x4wG9FyKgovggLCIuOmHv0cQtIPFDal6Y6TKlBpuLnxuM6lvoJPvxrniOHAA5X3RKXVRFGC2
tArjme+z+jyAUbUiYQjB+BzLdo/jQ5FZ7ZtbNYQ6AWzzV5L/o9TWF0LMLTcdV8sTX0Za0hj7HGPF
9EJXynKT7rjUh1dIc9d9uazCmJuatOOEVD5I6fh+EzwhVm7qvdAchtUnPrxmSPBeyoUjeA9s2etQ
IotzQI66Mz/VdMujeeKhXY5OT6ykiNRedcpxA64Nh/vgdmPrcTjK9Uhx196AgSuU5dq3q+MZ9Dst
8qv2JU3JBKuzLzo2fT3TfXZJSKKNjsyvZxRo2gMIeMuEQYz7NwtqyW7VrcwamDb/HY3KGw7JuGOQ
tpDahQRVc+ixMmxy2AaD9QJeQSraXBQN2WKzoTOOUeRSMq13WYrGSES3qd1wpZq+crH8ni78RZ0c
wENfygdCEu7sFaD2Ydrv3v2PQzFrJlNS/dl5dpSna0D0VcxLIxfmJNcAs1Ag6/WsYqahtjyE93Zb
93bN1eCnVC7T8TDWjFO2LXW1dOwZnd7eGE1QIU6sqZ8hMFd8FnZcC2EtTkr0BPZnanfHyNPeRGl1
Xqu0OgetxVeHgv4voEP5lkRlI7TMhky8rF0/WZldAKoQ2M3/VGn2miXZUJaB+aarp1ILC3QAl4Nn
6UEUKjIrK3k+EsF+FYWPxttwr9SKDGJg23hMpP3XqklbY1/nxxHs3X0ivzd6o7/CcOll7sMrjmvO
LIGWEj1241EGb2SbAeYFp+YKb2Eai6Sukkqp5BPUHA1m73xhsKJa83/zeoGXkhnmgwG939Eo/aGJ
lw3SVdTvz0XZ9k3NDloP0tHjKyX5H49XcOCo42YJc2R5kGAFYq7R0I572Qlx33TkT9viYTyVVuam
vJBY4qv5abTzn4E88wyoekDUGpJ2CM5FOJ3KY1VUoHLI3ufMsOVHk8iJ/HsYtzwEaSPcxq33DjPx
/WNEsDWlaupNEsyMG9ExGCBpZ4wdZz+IrMe3XIOw3CfWoUgPt2bIIjmS1IsXOp2huBv16ufaG1kh
SqKk+ZuyAiwVXkdFWOIsP5IuF1n0yR1dRw1RJP1UijwgcNpwSAFRvaW3e7DGs9m1GY2MH5rg+eVW
arbDK7OXPPsI0gFM6Ml0Y2PM8MBj1/kckl+/1apY06BICbVbj9ZwQ7n5PldDjOLCtiU7pMt7OJ67
hFSs4//nGu9iUA6U9R9/QPd7cKVgC79Ikn2VBSAROonCCn4BPVNTwvn5h8dwDMIor2AK84Afvp+A
/TEma0mKnzz4E8axD3kmFRb47o93ic+8HCBwSYVu5uqGXLYoF8mhDqP5mXN59nGKZGLxpRJSrAWQ
j+xmeA8BT7HeD0B6q0R4CAoZ7s+NHbcE7UbGPZBcj5vKl+4/lRgfmw25H5oqIXKnFfo1hgr3+RfQ
taNgCaQ1N9HHz4ZEFsZJ/O+nU7wUsBludhil1jDXxE6Td4F+wktFoxytI64AtCpUIxFX98WgybSf
iChPHOYRffObb1uRUuYxo5wfENriHQDaqL9tiv+x+G5DC7ZDUNFs9ot2ECKT7D8/N/PLT+nVCxmB
cAdR5w80oSX4SRMSI53tSZK2azccmlKRNebJo8mqDJABg/lmQnnqdLPPQUs76Md002JYtbtiRCGa
jl3+O6dAYsuY910UIdBKxdIJdAOD3r+41AlfI1ELjWkQ931mXi8MCYxjkv8qGuGOnmZQg5KpWbAW
0zfAG6IjiZF8BM/jrqBmwUJnobByL8MQA7Mcy8INbG1EZaj9gZwCckSfLJFVbyUCuFO2MhMEdYFY
2vDdJNFUZKd3kGOu2SB/JbpA2PBPsKhogNsPxjFcJX+gsnd2hJnczRot4x591tLmznYWWGTvBYXS
bQy0hmIoubuq5kvFx58XUA7eMPFeK9uAeMlOqCaTwmI49mMLCY50lsR2ph562r/nWXa9gNbBbFYq
ao7Evg5rGhc+PUAYyHVBLRQCYM7+03Sgf8ZvhUe6GhX3/H+hNLUksxez2cuPy/6d9CtJoEHNGMxD
8n3Mt9rl2dG8KA4+bV5g3DWd+PYLBipVIK7A8iG24U8V/egcVoqmxwrWha3E0z1BCHJL7lpgcftf
wREeEgeD4m3PM04MDBMbthl/LQrFk7N6LJSyJ20i2emPu2dSzCYo9q1Wv7HgOURDfw8OaK+STyr9
KJdcjO/3Crq4Skg3PM1X2lZDllR9OWfcxNzLupSBYOQzaeQpi9wv5ASE2Azrvn3XK09pKEHLoje+
198AyF8uJJ3vKWr4RVc0ssgn8xVnvrjyhkESVyI08pmhVSrI06VDbjdsiRA6Oubn5Bwx2uV0PrZU
ila0MLZzvVLTNcJIWwKIuj2XmF6+XSh+3bc45fcloBNWqGfwDvgAan5CwUd2FLsA+XPhfUwcA49e
PPz3mTPqaxbO4VJvTZq1ltdCqrPhEU7grhCHOhR/LAwpBgZ1SjQijbfBQ7kSbf50F59eBuN2ROXM
W72laUaIfjw2+OOurT4PojVwmYAjwzsiiSPuayHCrSoyap0RdVlA50bShwQLH3LdUg+7yS7/7xVD
QCk00Tf+K4VRq3A4NKFqyzTTMgRliVi19NmuYyWAqAjX7c+/ji1pr97Z+FxkY1jsf25I4GDn5S3e
YF8Er4qHKGwiQNOhgVia/selawYF4patrUvKu7T7PtP3GzveZBxnw3S9ns754i1VxIsbWyAqQYYv
avyac55RSQo3T7ZJN/2CIznpg0b447TKl0ZblwOesnD8IcqB3HeZ3z9MLz2sITo6OP39rBemyDWF
KaP1cX8sB1jUfWipP5XtjjTDSZywV/hqfR17jik9RjcsbTWjbID+yQFw+PRVEdpxjEZZymPEQwYk
TRUYDrf8a8i79pQnGHNPHZ3XFiWFQr52uPImpX/tNhLk3qMS8c+UsD9XLCZe9eCUqz0Ec4VDIbwr
75Xl/LVw51EiiG+3OK5TYL5yz25fXdYpl1rUVDMLJCSmLFNDlADuPKwJuTpvUJeFud89xxlt9VFf
ncMczaftHw1sCe8dyeIP6r2Et0YoaDKiPjDQJ9Pdd0qRAbZ1y3jIu8urkfVNmg9Mk4chYYXwK8sg
vCgvWIqRTgudd4cKsZ7PGl3lYhrSajapWGWAMgJF3enHbBI6POVZUUVjZL3C9zjoLzt+Qsc83yzZ
KsNgcxFD2M6Y0PoPgDGHrJskyLAt6BZmhA9yb+sGyx+jF0fj/IHq0sM81Ju6Th2QscJXgkuYI4ns
x78HkARDdIM3MpZGlmyAXc9vXipoMENFKK5V01jQddZ4ro7yXbscN1GHZq+xm7IpSF9WCZP+SR9W
LvKYm+hMzoXbwPE353qr71cIKy657oXQvagMXJOu+93TG0Fsl9KQ8KpjXRkuh45jHi3ntCZpULMW
m1aJ43loOBqsi017fWgBeVm5YdGvUZ58BgMjYMdvEcXVntfeMhdMWRfU/i5gYfIGNL8fPamdnlEi
DUsKJzDH0/ISy9G5codxNv4qvQPKPG0wCu2LIfU87U6MDNF0P5xcYUCABHkdZlgcjpP1y7P4nXzf
FEyn97f+LlVZV2oCJoaPI85g/FkF/MqYPz4gc6i4q7wDXxbfbiiZDw2wwR2r4eZLronqckkty98B
VssdChP0vJJzmCKc4N+3eWmW9BupH0NVntSoMTsuZiUJ/S1eW2eM5n5sQy1hLCaRL7QF1QQSje7g
fzmEJsBHEyz9FAccGlCiKp0uHZdfI1kGn6UWqJWYdLo+wK+HqlnIHOlSKTVKrUco4tF2gQMjwwqk
tkbvALJonjxZ85hgS9LzH54K2VzWhPYpEFxoWP81lOkgAoajvpaznSjErOPBfSvfxH7Auu4tAgyt
E0y44u21WcuP29XMrcmTkOyRc2YTohdVMQDMrPC2JSdIbzeXCywqp4XqK8amH+1GRP+FuPnYcIuw
pyXeo4jEq5BRHT/qVIoHtBra5RjzKjJD79lBRcSkCBaM7qi/nDOpGk6osR1wlCSfEwQEjwASgaTA
tOG8Cojlp1X9FtMviXNIgTuKwMlrpPwYnK+XbrdNfdNN86oLW0ii/wYeHpF5hnZ5PeCsdhObFT/V
8Fxmi6SV89t47ng1ns5GsXadOlpNMS07AU2uIYEdruDdSj7Rs0l9JggmQm2XzjBzeZ41pytv6koz
UIzNDmOHmJAmX6q/cUbNzjjnNBTriFSGUu6nrDdkpv4g+TvYgskJlEEBgeRDUefzbn+kdYd9EpZ9
ibiM2qirPtNtlgo7nqa/V22GiazoBTlmI/umUl3/HUX65itVIr8fVwtaepFsg1E6XVxkEyttR98M
OAdw1SJkTwxvmUxtdWUFEXfxAcLf1fcFjjAi0ECiBwHKxAkX77iBYyeNkzQkF/aKyFkg3wHsAQiH
e/qlMi9qkeRd8mR6ur2QLaJQnRPkCRP+gJa2HqX/Pnuye8iwGdPs+AiCR4QeaRw+PssLaKyJI+nx
cvHoSigS8Pb4skDcvOgVCcrkdvWo69qWfJdePjbsSIRXzOVjBs1vadM5n4Z4yRKcdTQFFZ24x3Ia
h0xM7dnMU3GytnQb8XYrr2UUHf07QzWcHc2LYO7fHYhIWBnA4NoEFcroFhkKTZsAp/Y28+jO4F8L
KfX2bsrhHroKNQS72I3oTMxoBfQsl61I8NPaEfEVIQFu9sjNYoMSJ1QNicz3zGqsZgK0JGd+RinY
+JkHtw6fBlqiqoIR3JtOEn2rBlz3fhP20YcJX6/TOKTuKhXdJjhPLem3VinB3j0cw1zXONt803V3
yU5pfu1ORDmusMIpB+JtE6mKcQXd/YNql6mX/3d5hg57mdy8HD8NyqZh8tqzIsYPWU74LuuIHT7w
CqX822cEO5M1JG97wYioEDHxyE+yKIFo6+v0+GcntdZHWM9Hidv+xdM/1UyceZWbJtDvcML0OhWk
IHSRl7YWgD9hL0E/LpnzI/ouv/ErH/v7GrTsuiuReZGEFC7zjgNemkrHARTpnHyDuKrwKARkbWMi
UD7xEtPgIGP4HDblycdOM9PjwDXMZIGTdygNCx0pATnAQ9tx8P4O/+J/yomlSgY/Vu5JRYApvmW1
90rQMy97U3kIO+v/fW3zrv+LA+2iu2KIR91DCVzi/JxDNcA0Qd4pbqi5+A0SQ+QtaQlOwU3uzqBd
Gk681/naNuwBEtUS4PErrIhxFTPkxLBMtuzVsi2d44q2qvfXTrvqLh9/brTuM5T94Zh1k6+T4/k6
1ikPItwVHlKacMOlAp8a2seJ4C287huukhWpe332XlMvu5y2zjMlCGZUMRNaG1rjlO8p0l3XjGgR
VcPT0UYB2QnyKn3Bvb9UdcPFDBBAjSsow7gEiR5QjQJdnrexwCXDZOdGgyLM1Mv3bkVpT7ot9e7h
ziujBP2yQxzeaCfU9/tuijxQeOXIhcWVMXXgBtms3TQDXiT1nHe4COUsw1ydaTUPzxoh/1dRc6KH
i1/3RGov37yLgKSECNO/YBFUcIOcLf9vz35931Zje0SDGsUXoORll9EF8plan0sewNOGkaDsQV69
cFgpU+Ub5hjWdZ22WjeEw/NC5MyVTfnIRrqkTeJxuOQ3m7gQlY3MyxYzn/KnbQ+WIM+b/FHVCUWO
M32jkYIAnIQfKFrMIczGWb4pzjuIm+uLZfK1Zwf22LDTGmPZPkjxlUtv6m23CQDQLtqBd+cIBOuJ
cznxtbPx6w/o8BtqJ6xihcQfEeRCnMSe5GeCS3nn7+Lt28DBAUmCFmfjF3zy8KzFHQVdcAkcdikS
uzswCYwxMYUZG28RAW5z36Upzk9jHbepyY8ZFR+h6+l6Su8jkd3irCsKwhsnEJ2K1VdS9A46zqP8
kRhaW8lTSIkp4LUlElEr+r434OKjsyiJAhTmNWQXd0ZETB7zQiluh5fVrbFFRXSfBqjp94Z1Y7pL
HDDeqtLk0kyRKSXPrhTNY/I5fKNbeP1OnBoozNVlII6T+CUKAqX6eIR1pxIsM70d1y4u5TZ6Phz+
fu1NyB8UutKmjkcdtF0Nowq/34couIBU/CJYwd7AXMNVLqyHa4Hzz3Emf8uiXC24eKKmloT2sY78
6WCTP6XeoQ/Qk9l4v8p75reBO9mfaK4xI/LEBJSonZLrWc4p+nBko4IfvHCjeTn2krZcC3eMMRwI
zpLY1dro870skSqEFK3ysRqAPGnUfEwUUzOKX/SL6zD5eda+TzcJumh5DmNzlxiBLuIJ5O0tsYcV
SjvkDNSHzQ4aoT2WSP9a1DFp/GxTY/dV5ja7DJxJplmOyCmjCrS17rtRXsHDnFwoArHEZaK6Eovf
YqWUoZ7LfbLwlBwlGPUKjaDEYLb31oRlqJQRYVpr5u1YGxN78Z+x+j55nuBSESk48tI4qdxzog56
cGHXsfSm3XOxqnkhTLOzHil+aSXU8ewIWQyZlIuvfzWP0X6J913sJtLcdVmDUh9C+EnPVU8Gu05y
IeIBkfNWrSw+QO8zqQwTSERaxls/krsAGJRwsrNs73JV0H+T7ec4edmy6wrxupkf2Qnuy3StjD8R
wO+yfubzex7YaaeSFqdtol9Wx2iXjFKWTfuRAONE6/hUyp3n1TBgPk+LPlwQ0nSNqci6Zmd1UfhI
YPYWDpXqor+xiugc7RS0epEsnxV0j6ohd5APOKeeyh/gNqYOWJWs++XgRAGiWPsWRpnUJVVlQyhh
aTZVwQPExeC6GMwvAusGs6UJ7znW2+zgM4YDakyKtrci5bnSRrvWpwJy4K4pMN3yq4EO0wZ2oghn
XRwqIxdq2vq8pPeKsjZxOo5VHZ7CwETbDNkDUVbVDz21Wu57Fo4XoUFZnoTmgQxwTe1fpWXzXHDW
LCmDGtWRvkcdkXn6XVLe5wr3NH0t6hTRQvKAm+xSp5ZDkGBfvgS8HrF+q2owOEXmuptrv/2VuPYm
6uU3CsfCehaciCh1rb0kW1bT9wGbBOjiBwN0FrhS2Bx9i1BUlzRIxqKvNllVPK4PH61sap2mYIa1
yti/Sw4M3B+ntf+Svc5mPEwUzOrvlY+X795fe0gZ0e3bAoj/qhcorS/SXdP+1sau1KRlCM1hFbhR
o1lJCrkIk+svLY3uvHsxOTWdsGnFcPuMNKkLOci4fSR0ACSJSt1B5ETItJ5LrUPX+F1OeSrfOi8e
WpXAYQcEArHrs4J+VjX52+i+6Zfxc9Pl3ZES7UiKnv/1cariiWJzn2wNeZi6iXwFUJdRKbfQNDM+
CIYZ01s58g5sI+q1WRYDcXzJyIfH0vkhZII/nqfFHBvYKnFNoR141lcQcDBoRvMFwhcLmJNsadoV
HmZZb0PqbCiMRzRH7qxhZDfbylMjE1PK5z9qCMeZ+GuREmrPBfhorP/+RLJhKKmdXChM3F7fGlPR
2wdbdLMyv7xosauoXzUuVN6l2J/tgkTd3wLC64Kxr7m4tnM+mkmmNkVijBfjBQ/UUGv/W6joP70G
g+oUMrPce9dk4XV94i9pPq2ZbZXzqxfM+ZMwnyS/HFbZ1BpOuH6VdpVMuNpKJnZCRN4lnIaO0+Ae
3s5Gf2+za5gklBycVgkTaNt86IorjlL2cnpPPMsZAPegLfdDXtKyq2r04BYFrB35tAuH/fmCMWgY
pp+jtK53drbe2WoHWkd31Fq6TR9vkEHP1tCTw/1IReYhoj+MVVdwNxmVEgsD4FB3CxbmT9G65a8l
O878KLrd70QjnVl+fXpiLWBfZd/ULgauRl75LWyMtQjmdOIYXvIamjev+GihkpNu1m775HAoDzHw
JREw7myK9d2goZFr637DYJ3lDMWL6h79hv4juXRLfayB7FKMnttegg69CjDxkCR4iWAQOpuDw67b
BWOqvnpokkfioG/FTJ0QkPB3JnDSNQ2y0FCdJifWP5fUui72eNaYbtAXMlDusehY0C6pOvGkUSEJ
LRSLsfrXkr7uYCB/LipgAwVcUsqGnw9SqKdDTNRilucBA7vWeiUS0QWfPPX3DKVSo2GPXNUJepHZ
O5bWVaNHoWOF0mz8qrnZuAVHyFFR7/Lj8xwZ1M9xxDnIeTVwJOWPzfmNbSBuKpNAjw0MToE2m3Fr
2G3NAkD66S5Xc4MHMLmcGiVetcAk4ByoC7ReuAcnUYPwaIrKL9p8ekKthQBrpR+sW6rXruVNHkJ0
IVXVTXhYZF1FtVKOYi8Jf9c5JS3tjKM8MKHxEdEsjJ1iJUPZfCy33wcU2/akplfhm2fluzaRTOM9
JHycNXopdpJ7nOUzQZHi2gU5hm13okceR9H6ScEVPe2LEVZNbjt5ONuNcdiMsID6xdEYEf62br+u
YnHzVeqnbfe09chMyFipfk5A/yXv/pybVtuystYdPLsJcMQS+b1X9zd+3+B6x7WjLQeScqabamU1
X3uB2IY7V4vuw8xZnBYw9rsfof2gV7tdKnkgY7ThphEuLN30jpPtNyVyGj7jgxru0UJ+0ES063F6
kkT6NQBB3wbgKzNzZCeXRiV9USioPvVCBUESh+MbKie22IgUtz2vWmx0RC+ZoWH0vuAy6wcj4IGj
s0NeomNcNUDArWulo+Pk5yriP09sLGs9gJxBGPhlUA3zXi5v25RUYlFU2uVnse4rTYBUrMWD76Is
gc+IeOM6Dbl2eqaW/ilKw+EDmlXsKmstcDSP3HElYJRzQnAxXyafDDdoVWaEA/FPbOVNieUHrY7K
j3ViQm/iBOTTj/B2PJxrhqs0LCXPKYffI17zl5lE2Qry9Q/byZZZ7QeSqKarqJCZ5J36xAYYTUU+
eNnL4UfdvaJEcZhCKDSl+dorvMkwQseOpCck1WSRJCnGTOSEhapucR+qy3LYg1JtrnfteVvwXatC
KPyRKFALoQei/Bm8ckN9HmxISuce97pwwSEr7MKBU/h5UguhUS4QTBFwnnqZPgp8HZGTYM+DqmAE
244vtAvgUyWTwAcgKEIr4ZbZOJUxomZx+ZJjd0VSPDYF3UZG+YvuJz8pplFpphRyXRjF6JHkyhrX
92NuLbIXbMb9yrtpF8BXq4dJviPwN2EqL2oHiItA0ndumDWqbYPrVj4TjiPxzKdfk6w+rNyEF0n7
1cx4W5itH1ybL8gSOMNiyWqR6SMVZwAFD7+CNpksR8iZWao1hUg4yOP2Apv7rBcGK5L52gJDioUB
GACxXarMC6iwK32h65A70c4THfcBP/FwCEiphy4vDlSB9q6OKBzxq0wszlnuSSjBuVBIVvjSNJgd
5o6jxtCCtlDBI4Et4uRzwJpSw5IQvu5q103vfLVfWaWt30HDctdKEY7J2NP2quEX3DSNds/Q7fxj
64NgN2PGvKe89yw71jWydcoosWysbCzKGP/OwmWw+bPiWKlAIkwa0nWBrHNzpBmTGUljxii+EXOq
yAAMpiz0uDzUHwa29pEawPehHSG/AyPT4IOZQixFYDryweY7l67sVF3jveHihAfMvYnJ6el5iQ00
zpDSPzhshtGUGXtjyYPkHvGHLUHtFVBD8Dgz4bGMofdctWwXokokIpv7uCgikuBgNfM8sLxb3YbO
5IGevsLtFdUAzstnDX2FFv46JlPlYyRbTNr2ISVIJp0jjdB4qxMmzTw551cR40Wya340P6abS3P5
cl42+9hwGxhpM2FFw+6f3SWOQPj3P8q+N/YbP+ZAYCge7kcCraII4vMABq40+l+7lFcKYcCjDD3f
rEuHcNYki65H0o54KioB+wLRyG+AzU15fcC6FbRtPnBrBYjeemEeKT9DEV0iUoDOUJPhYEoRuTcb
z4qCxW7e1S7EU6kNwVfMaqythDfjUffPlRSMy7kiPUGqkpxMxYADnWPrrh5qcQOUS4I4v92WNGDO
i/IvGP/9xfEpplSJxJViKx/UqsqBON1754QvBh7MDpIs6nVeKFjDUjZ5TaDRJ1rn4jBL2ATFE4Xo
kA/74CSnxiS58DG7yVPuG8cvKHm+JZ6KGxvfZWHDgZ4WdFpbcRamoF9SiXkW/526YIH0eXf2qJOT
MODleu4OJmce5twM7ZvHCHqtRlcd9S4qVrNpPRyj7J4wSng8TM8/VCerKnxYTtVE3xVX8ZpCs1om
gHqrQeBynZtSaJwSHQixKDeNLODpX/pS5ZG64m2erlROZ7aqlD6zt6YD5+sKfd4fVZE7OQlRLkvn
zX/oNuc/F3089zFxInfjzwX6MpYSCW4GnGsjOzWrLi4GZwUWmyWGwrwUafACl89PnrN/ZPoFXAj3
z/brc+8R5X7YXlIvQExZcXqd+slE4GgwtphRwCSedhbN59cHObGFZYwua/WGN3Q3xbENCDhJ3AS6
Hrk/9NxysAqWw1O09ta7b2oZ5gzpiR5noRiM/Huo06bl2xR48c/2h/xLpEL43Yxa+f4bZOurXaGy
f5oHcLCln8Ts4EDi2kgTxIVlh9ZOWIixUR+IPepAGha3hjx5rashx6ZJcMTz34lWJm0yVy4M5PCm
rXUGzu3TOFFydBwp1cuWhdqvZ5t6/LWQLoM8l6oPlEf0bAXCOwnUMtyHpUuK/qc9KzKcV7vAXJ2C
1IW4mdvWr0J6UgkRaXt+GbWIXGjoUyyygXiaEduW0MWBDExL5QoFrSCCA6oFk9M/s6ZRQSVpUXON
QGTAegt39OCKcESrBVKWSCfc8YOoytpyreJxC9PTy4EFTjS1rcB2Jpvy0WjBhAcJkvjjBiKn2rXY
P4NZV2TCHOSUgnpoL8NW/WcOcofFFrk2zwHz2oxP6nmTUQGzjRFTGgGlksl/mxcapqprc5z2i4cq
cHhYu4nQOmZWs/VY5q0EokL3Kp+23osRGvgTrS1RjSzI+0vK6yx9zvHkVpXv3qyIVAIM9zUsB0JA
KyNWHQmmyh+nGeqz+VfFIfVroYmm8LEJ29fpz4A11EdWDNG//tPyudPoBmEbxEWAiq/FnakDVHG1
mEuRFVdmg1XXtICBB4XNJoEOklchg4u6RdxM3stOadwLDM5f6/ywnZ4kj942+ZXgqep54MyeB8sR
/bkFkmYyGJLpfY9Qppo1oCUxIv7/17KTlQLQQ2YsZmBbxChh/Dk7H1GwFoo9ug6BNJdURP7TAIJn
GZEocZ5SxKaYTDWq+YprLe4gZxDFrso9X+MYqJYEbajpTBaINZe2cKG1orldZlxNhVB4tYcWyRmT
1k2gEBz3V/Sv5GYuKvGmwDxqjL0rRpOteWbTxbJPhK021QgEc6QLiLI4gnMh+64JtfgKIf+yXCju
daG+nHCd633EBt+zQi+xaSeAN4gEYHFk9l9syLMabfLFBbQOXFF9ckZjGL+1l0PmMHZxzXCxlP+3
rSA8ZSNab6Wn5uGgd1Z+pb8pB1LjK3B/eM2cCUdwRquAHOVg259lXyZis1cRdrWYDWDC0kIKb+lQ
0vEhN+PP/FG8RSDwSLeerzfJo0VYG3ryHE7dLXcsFjG474WysNTrvHltTkD6E1H0RTPReK8CANj/
CKYFs45d/NnCJNeDBZSbpl1Eeqv7ae3R2VTg6SWyWg/SaeLhYx4DjtKXAJTX9I+Zb5yyUKRZqce0
LZYjraR/nP49U7uen5FEgDkU8Ucpl5RwtUdEQZLNx8PWpLfL9vK939scNVoZxe/kUl5vA5CaEEhn
lOjcZ79IuQlcTJhvEDkre0yMVYkBl2sbCXT6m9OSQjg+tfxN4/Ae4yetASpdRLfQuOJSrb95cciL
Ws9oGPSFXegQy9E1KPfHGrkLUqE4BhdzctAKmK56+WlPGwyCOnBROC6GOe5scZyXY2qt4OqRPIJQ
dzk+wCwOzmwpssk4mGuv/loiTezo1LfQ5fDTVfoAjz384ITM/mBRhmTlrf2KOBIablfnEh3sF4Bl
bMo0+h7rn7NSYKyz+8gby9zZLoZ0bMEtT7a5VKZceGrwZ/KOvaP3k+0G7JirYrtpq6rDqdyhtOjP
tXOTJ3RP33YR8oA4yFtFG5mRdPb1UeX1Veo/LV3clmLZOb+aT20mlyktLO6h5WVA/AqrgkUu6rZA
N5fuhQ3Ias862iIuC/P0UZIB6L8J0f6DkHiuJ3AHi1pac7AjKeEo4UpY/FHBzr8z5FyApt8FYW/9
Wieg3rxkLJ4erREAd4QPllJk8p6sJesJtc199UFC6+DTtWojsxzPK3hH1ghZBLeJqw22Mh3ISf0n
eVSucMLRPuraCIF1zvl3n1iQ64AlR1LvlqbhNn34fD/byDKYq0IVdugE0okxdLkp0Ir3Cd8S+Wf0
ShCqackowJOdhuiijr0ZyfQ349VHExuEo/XKpfIP0cgEePF11Woqh3kNrjRmbsEwoWX/reUhV+0q
/lFu/HI6PbHgpcU8Rrrd0ijT0Bl3EyiEy8zPGqGPL0yuSMD48Ga3sVDrl+gLX8s8WyW8CYCYfdeN
Yd0H3Qobg4YeZaixuqEXa+tq52C1cLeb4tclyaSCL3MTM1hyglfBgZ9O0KfkT8jYT+RlFLQcSn9e
ieOOwmmTE+e8UDwo/ct+cyWTvAPNc4cHdHUKooYmI9rxgIHAETZNi4xJZNvxf12x84RtLDoYmM9u
rzAgDaSp2QibX5FQrlGZqFQNj1qD99MYjfbhewhoZMsclc9DazJ8Q8EcDqzDrIf/1j8ZthVHylZo
uoeQ/TbLl69ZddHw5eEwLu3s98BnKnKwBtNmXFLthiNZVuUKwBIS46s977BkZqHZqo/aAnAB7Xme
hRpfsp66zCbQSF/qdbnbr6y2JDlcRGKm/9q07//0OGONrSdGqkXssbOUwL0gtP8Pwu+YNpcEZ5R2
PgAs/OdRSf9qYkF1J8GkpZ6ElHxcoJEI7E+P7lb8sVpNz7qlvKV1VzV15sQHrZPJzyt9Yi4Te2gg
FL1tSiSStBBm48hCCNl2cY72kpTKisCw24zizW3BRShvNNLpvmYI7Ap4w0NLucZ19Ob8l2olmlXe
HRqu5SzsjflrFlO8jfTCdQ0I3FWCmra022sWKpLSUYCAqFv+8BW8KO3bAA0v8OcZ6GJDuh6VcFlm
p4+ZptVwY/02nZvEwE8wFiTcL0+rdpTOFXxsIkrQbXsiMKdGChahcmxuwxHaYfgfa1TpegENQNN0
d11u7O/nY48M2O5ZaXIQPrGYqhNkLvbX00b/FYK2+WwY/DmOEbkwE23gc2bv2dL8zDpM39Ucu535
rhZxQ6uOsEFGI8NKlnPKw2rA+cAGVSeBvA0WMDiKS4drsz2/nKmSSmt+oiyfCgYgRlrE+TIETUum
HQ0cNDN/wUyAzxcQfFjDm3pPEGxR4D64ElLPOIycahjwiwPAKX1C0mKeXNmEaQ0LgQ2IOHyES8Bb
68nQg7UTUiPKDRenk4FWyoAKvPvAeoMef7ZDe9Ijl+Wa8HAAPwaQ6KJ48Xgflswd2avgdIc6+jym
sj2GhqNeinqKqKDxRy9XSOhCsi73AZnGTjVUtK3flp4TxpiGlgESoNa0VY9YxZzqIIc+OzePOzm5
Gci2OArAgl7yq3hyWmZUqg03K5+2byajSY19wfA4lSKsa/B2MkDn/CNqNxQqwhXuIx31Is1y9873
JF37NtspPfGQZBCOC533h1+J3CMiAl62+NX8ty4GXHc69a3bdC26SZtVlMCKxFynjuGFLZF1HuLu
uyq+TRrVCkO+MtMKdYbd+wZ3e1vD3PlMDbEPOeCqB/3kMcXGyOVsH/bbe4SD0YvQajfFNn4jJHg8
ciwh0Ta5C0pzh47Cc1kjQS/iTFMxaeBRkuzUDmUoEoEKjmbaYJyZe9P6/h/2qN1ZsLCD+xPqPg9U
qpdTUBL75GW/8D4EkVabkvysmWHh/yTZlfHroy5QOlhdyfrpZHTxjPtQS9OIe+/I5Af8d48YF5DI
RVyORRbjcLfikNqTPEEMlCzykj2scD987pYDnDoRvo5KaZoUfL62X31nWc+/BxY5Cw1QzlyeVqKQ
Xx0irlAPtIOo6GEQI2HmBdnjNsvHrtOPVW2+Y6n5GAm/IWhuK5Wb+bZ3qMbVPaidlqVAaeC4SlBC
ohTXmyuHd34MyRmvkwGJIOkB3JWGTDs3a4YWIP+J4dpgII2f72KmkTHb9DU+wLgkDp7ZLlRYe6S7
nWxuuXSUMNT/Br9fptRHID6qkAFvp6uO4gFzivXlZFXnUaCuZDwO1UDt1yORM3kS3OPK7DtYE84C
N4Z1rgXwYa9qS9PT2K/ujdaga7LHQI/cx8AReX6/bHlV0wsxd+5j1l9PcqPSJDf3yWdlUO9cw5u5
Z9tvLhVn7wzwb109EAY+CFjnSn4+ltJX4Ino8apB6E3D8NUtGKg7PAM5HLnaVWN/UHMzE1EVyOFP
JqSCpuuFpde3Y9Bs6/+hhb0MM1CeIE9ROkyfbhJyqgaZCrly9l4CABgE5gfIwqW0AvsLMp0Y0grM
FGahMzKWr5Nmn33R7exC97oUsDl4Pu1qOJa3IBnj6eSvfGRfhcH9AzoKqBIU00pfTAp39D5/GFR3
zmN53hUUa7uQC1jxGP8JpkG9j2kwfLsTWJJtFvNmyFbYkxLa4bjr+L5k2xHipxzdspUzczsyuPay
gGNKf5B62EMymhnog5TGmhBc6uu8Ikii8JDYzWPDiWN/P2Q6W0ajlHNYVtSaXXcmJs1qFoiqV5ns
qUCkrzw84ei8SDUCzf55S8jUrA5QKQN0OTRNvOc1Q+9v7Z1oeg+DS/wFaY6Metr99lL4St9RDGZD
XYdNbcI27PxGNSNfBpEcLMdLJeoP4/tpYYwvp/5qYJWWqJCOeIzyMhXVGRz94heGU/6EHWQZ19oA
x2NeSC9q9oNeQ5eUfec13Y6w6oKn6AQPTpbUl5YdBUUkBFj1lhGFbNmwmCvpZRpN3ZT4RgYY97sC
V5uHD9+3iElmpcsYPeyr4an5CQGzJvFiaeLir2+QFgHCknFsDlV3GevTp067pTzrPnzUeBY5n9cw
Qxzy1C0SRo659DGVhbEn8CvcedLkJqUgKqoLdYepW2xVejtv8LQoUNA+q0YwNb0kVR1FMnWwW9Ld
4VoFsm4bC1NFTV0F1dPmuT1iSSmyd8bBwB8zcXYYwCvk8PXcn9+rAjibgC1OCa7MjsoPgqvPktrf
/nwqJIZnrY3TltyhJyPzEQZwy0hvoswaKYOEXRAXJL2hmFvxYHgNeOrm6QcYVFSfBx4H2uS1YsXm
Bbc56U0hvouW9BerursG1m89/GoJibVg1sq4F/eoF0AYUY9SorPHAF3tKiz1kWcNBqPPgcpJv2B4
h6YUBCfPw/gpLG7mn1ObnCwFoGH0vlNWkCuPe17S6+z9f/9furD+2vmKSxvF0oyy+2mzaDkj0mX8
9Xc69aTCvkoTIG0vuX5VGJEsrJpbRaruogTQa4PpkKZjryr99SFugVR7Fl6YCNDBM7OH2NdJNMDs
r4kkAdnYF4rLk1LBgpRecGfSJJb/XEU5oy8sG+LCoMG+V0jkkb0iAWoN0kNUi1tHYC9RcxRCq9vi
QKhpJNm0NUKyk64qPk/hyIqDNmzTia/+XMTzTTsuTQUX8aFWUcDQGsvwuYOe98DhLhymj8j9kBQT
RZcqOdPt9PQhuEDth7w/Uk/D8WgurbKFPqnOtrjfuLrvPATT4WCQOdT9N8l+gQg4l/bCvswPZxHp
uyr0MhQOi4wu2EDVLgGkS5I+reZSTw7Bti5f3RhV+GKtTzFKAyiY9qlF0JbCG5fyfggRRzcRSmqm
PFTgvAns8ZGynJsbIzn6L+tKeZjv08HDZBfc1+4obAAckpIsfvSHD+egZ8hxmjHM7kgw5bPCQdeE
N4IV0v2KaSU7yIzBxToWwxfgaiJVR8YKEjoZaUPMAt/eHxZ889oIM3zjuHpluuPqz8pXuPg+y3df
vBfRqP3mPMYg60Os10opjqNgzXtgNjzfJlBb5Pw1XJpEfwlJM6xIG40gdHjBYnvDiulx2VLxh6Ak
i3o2QybieIGiSOpDkg0pW761CX4a7lfmgHuAM8DoJXwdB0IoMWmmuUoVl6A73h3O94PrzpkJ8Amh
Gam/nEM09/s2yerldIutbEa92Mx8alEjPJsgArIWS4w2hOQohzAjBS4mUwP/9vE7oV4fYYfnSnYw
cAasp/e4TzXZ80K//xYpMYsh7TiURFrDw2wvgjSGLUw1Jh4bI9kKWNt18P4jTdNqQAnjhuK3fG2C
pNYE2LSNIDLBqZe5JXrTnTPjN2f7emQdE048e5GgCBPNlD7VfxN+FBwvRhZ/nAoe9raQ6FWobbow
oJk4ozc0cO/gArUEUI69v0cbaJL0HdZh9YeCC2mN52flq1glBuhWEz5/5+NWxgSrUFiziRlTxT9j
gzK5xbn3VZaUS8PdA9HC1w7VJWxpP6NH1UDfm0NQpuoP1ZK3dcc9i5zGQLKwYP5WPL2fx2wRvhef
CNAOqHH0UKJKCr9dqZMxfd7+8yUAQ0/wo4qQkGctMx9r+uYC8Agqp4cG9f836bmXOC3MP6hcNzzf
DCU0i/voYb6BhHQje9ntOnpLbbe/ibjasZnBuZ/P4kD7NqWf0TCTLtNnCL4Hg899rdoxjVQgRQAL
2KEPqg2IhqzHtP/yBzA9KGFgigsPBD8753CBi3KqVblGdGus4fLXwjaDdvC5WG8CccdHSjPa8Mpu
+meOyMoWphLWYqxRXtxuDVTKakr+3Pfk9aTbfQvN2yAiX2SheDFl3iyN4HlwfV+iWKSUgJprfO5h
Z1jm9Vxu6ABWcjl2VDa63hd8LYzOme8tjwEkAFDOJslsOJQ5bB5gWOSX6758J2IDLrz0XIX3+1zg
pVFXrCHE3++TJAjWXlOnsc84SMMyNYETjHEym1yuK2AZ2N6g04RHzkJYl4REpDqbhjMj7aFUfDC8
8crluv1fH+0rJBf/nkyTKn0vPc165rUIpYRaGpwRzr+MiMbYTJzrxKUICmakd/2nOn67Clo+FQHz
PpxbbaGyKnZTe749pAlvXNoIZYBpSk53pzXZQuEfTaYpZNMfX4BZjdTrNpoYdc5uvEcrjyCnZa/w
r3P5omopUENhdSo1W+t+6iNW3W3+lWEvSRlfoyLKKHykMqsztWIDFSiQjlR8yn2q9qKYUoQoGrZ4
OCLQk9LdihYdWUCIKH371gJ0Yclh4KTiy+d3ZCm6FTlSjJylNPU9j39aqWwJ9el3+sB7bodsNSDL
0TZRy97f4z/jFnYf4btRMhIea2499kjoVDlI4PHHbewe6xfbhPLpbJJN9XUTwSKl3b/roTGijgo7
PBKGYmsbYIgU3Ux/BibxJMhPGcldgOCOyfkOB2MDSjPdHUU1wi3EQ8H+WrdQ9RvBYGr5/LVBW0SM
nUVQeZGF/63x8wUuQDsUV4PN7WRjUJtMk0mTQm4kcCKX83LCLfO8EZHR4Dq21f/6qVOYc1xpBnTP
TgRPYPQHdlcczRONWqcr0Ncaxzb8t5CGnq6TyeJzlr0Lh5P6oG/cQd0VEHLyFiuH/WtZF9fUpnfS
Eh96IgOhiVLG7cy39EwyfATEtalsFFBr4XoQ9KtwSUNxkjhVMt1koJmOYWqLEimlkFXWWKDZ62o9
ghxSaZHmqyvCS/ozA/a2fVdLllhbaoKsNIXA1Q8acsYXWDmfstfLb7riYQPHIMEjrkrQopXoViFP
b9OK3yLiDQzqsKe5MgJOUuHJgYxARPWwBClEnySVlgoRnuWxRe+ztRQWvAHb7KfNoidecH2peaeW
UjGuKc+M4Wqrsz10PktWOgDsyEIHrYpf5sqZkaqTHZzz0pILsm4z2WsWwKvbgwSuJZxJirK5GfT3
kWrLfvSjr0FVQ64hMPab1pHHOmd7ijuNPofxpyhVNf1MGO+8U40sAeQtPKAe5SivTpe79qC/BcFE
Hm48YyXNb5hq/2jWu/Gzh0S6OyzNqv3f7TzU2+d9YWDfufuB9pB4iukQehiSOVLxigNruwQ5TyAt
3k1Y7HTjB1epdHzSzGisvWIBU6EdCFNQ/95QscCh9Nt4qI++Lf69tRyC50X7rmMqM2VCdTO1z8PJ
hcZP4dUE3NvBJs9o7mlFhJp0BSNhhhZkNmScx2TU8QZZNUSu4k21Lyi107eVeHO+GzsE+iXRZWQV
NU8RMDj1WjH4XGzdCaI0qqCRQlh5YCJ1RHBjVxj/9+jI3u6TdHs1fB5GJ0neztXu4A+Stz1di9yo
QhfTKNAr0ZrFzJSUqXlikGOGGBOYdJj3wb5DDbcWHucEmXqail6BvOmEMcYD7hHE6atQXjZAIBK4
T5gf3lf8wtWP+fmYXgdl8G5KiBgzbCfFhhzlq2HozEl16sA0b4v9eizhMXuYnxHIuU6jF8DpxN84
anzFXwRb7UqL7TtTA30nIM/wyAyKLwXJtzrtXL3ruk/zD6HbUJyszNoYnuyaCqpLaa2yprPuI29B
EPEp2GOSu7KrQNgGgmAOFciJQAi5Sp3hOg1I1P1HUTUhPP2VJddDeWGhcMvzChNky1g7t9BHS590
OXNxFKgC4Fs/U355AHfY/D/+M8mH1SCiCpaqL5ubMnrdWzXp4/xh+j69WCiFtqzKj+oLgyMNWkkI
4UG+VXWaaeJSYdKu9d+Njbof4kaS4rAUz2uctXYEsDfzRpr8qqwzd1KenN34lSRj8QjznWxQfp4B
YhVy1VeNXy8ed4Q8AWKnF35hRa7ksuQzIwvcRYYGX5q7yJXvicFgg1D4KFSfsqoLjFO5dTmuXqmo
xHJHh2fTOX0ekdyAuJeWYg+A6bDqCph5hBaCdOxr9vaASukF04YIGooYd0rYURuFy8G/CxhwbkdU
gg45IhizkZ4TYgytWMtx4UdQam2tI4T1mfVz/rknZtkktm5m89xgQO1tqjWkmJ2Zz0bNxviPWLTi
Rx6/Y1ETQzMLAzNvJEOROepqMjIEIFJIWi6yZ2clFxB2d2DqqKqahC2M4WZjrT1qvoMX/0Wikw+R
UIOXuvxuE1IFqfyTw0XmcS5jQE/o/e9glqavi36hY41ZIwLJkJhOP2gMzYkVUCTa34nD068IUZdF
vT7fzYNagQV1c0FEjPUyVyG8R884w0tQJsvSMWid2fzRlLV+RJxEOcEXGiJoD6RBP+2fVohvj3bb
kkjH2fjx8SIQ86TG6pCLKCaRjwFIvPT0PHp4U0ly/+tNNyrelEaycZFZ25q9HfAh5Lk4UPWpzV+h
VBftXWwcYzF0cWNV3XAu9GUCbyzRPiV5Dc8bhCp8tIRc8jS1eWOfU3uyOywhFt14fnK5HA7xy2ia
Cz4hXbPyzP+aAyNEAuoz7i1wLaOBRz1yDd/0VL7nTcJEf4EjijL13GN5uu5Yf3wunsd48xb/vfjM
Ii2YoQxts2KkTLs6cZOXIw4qCnVgFpyzYuRgSUs+4Z7N05JJb6wxnDUMBbhrGEIr2QNDia2bYMN8
0/3+bES7VKTXOxhRw1Z+HzHTWPfLrLWRxVQ1i8dMYZUa48M+t6TTR9a7Pnt0SgHE3zzqka0R5QA2
k5fLaSlIaCxQw0koBtnvOEZ4TGkppB4WY7FiWalVBZIkf8oZlPg7gOlHWvqho/3PnXfNYLH+V5KW
hsA68vQHESnl0Ui7v2NIZ+EEg2ixaXdFK8DHWxvsrCRwpBXn30lD7OhsGFaDawWbq2OUlsyC3OS8
QC5CHQd+9rKgmH+v4z0TQco4Dz41LfC+wLyu0UCUkOEprgKRNYW+TIt9gz/elkLUV41ZNWOIwRDD
Qie21CPBM+jxkof7ufclJdPBUmq1LcrswEwfk2ZnMiaCXiKDTw/enUqB2kYburhqJSNTgvkyjc2Z
SMjYXCihQtDozvbumeqxu6uPfmuO1FgPAX4Fxlg/G8yCxIYLVgNLxi3/R4IgN5yf1Ea9BmVx+TUT
bfNIrB0olEeR1a4PKX+dC97KHPxzYh3jvJmimpfRYSB/ZqG19M3RfTgnXZ3YjF6ATDJHtL3QtC8I
TTqT7ESKMNWc3szl/OyN2HY79XLXAB+tSlV8kFOxB7bXQ426fkoXM9LLUSEOMqDQqSYM+D34ZyoP
I3XWp+EjPSYB0Fe0wJ9A0ymK1lzkhPXfU/EBreO1Ny/7w6Fa5T5/cB3BIGt9CWHYmXA6FurboQUn
CcmnnJLyBqfYmNXljULV5llmk8wEEyemZSC6C8Xi672Dl041vZUAYvz0ex7/smkelHYK/z+3cfja
mliccuYvOLpkBpb5p64PlQyVJmH8bkl6Z8fAI0phsdXfrreY94tY2xjO0botDcEI/jnPfSnu1mou
9uzVydtV0weyLQdhwmtcJKouZsj3uj1/+qInsNV4m1/8Q6SAVd1b4fzhiwf3u5ugV0uu1TyQHCok
vu110uVIAlL127ttuckRvqA4UZJDvWQ7p0j+pL6DlRoGklt6ICMif+xS001ATfiOTLh82ENRcd8z
J2M1X0RWDdn0njo98ROV6ePgNukA12sxLeClzEyM5g5OVcPP4RZMn+oV+m26nZehc/hXEIRLbziU
655InZt7WrJ7igD/4zoinlGbafE1mRi/3jaJsgnWquITjnCyQQ6U22NegQ84rZlEc4y9a5Sp7Aeu
oOp1PJgxOiRhAjOjbdtNrwus74fHGJreG3WxjNJee6EbSFAkfqIKSWvU2VchyAl9xxRkfbemrZt5
NpP0iIiye0dX2xAfG3bOiRNvjhb0yeHPTxdrr7Z5PBE+MS+wcQl5DqsjP4+IGeCDNHWRYFDBOS+a
kkeBt+pz/vikGKlgqlS3ylgRH7rRg4k3hGBUpvx0qpCnEpF1+PlldJ642dTPMrpA7GFuOzC16ATU
pOOazpUMJc5AvOxl0zkvWSqy3GpKch+Jgzdi3DJ4oeyUNMATirpKnoPgYYjLf9VXh4F2bH3yI/QR
I1O9AkPh8UyBpZpUO4Jc897gyJlqyaqGO0zfdCcxy4pl44k1RA10QPBDDPmrlDs08IYjywOJ7GJd
qJnHUPKt/ZnGinDXqrUkBimFNqbpMyZIq+4HIcSWqnp8rnEofgdbIyISr3Oi2ACHQPkcekKMRfSF
vId6LnjpSPv7TxiQY6LX03nFHSTfFGMMka1v1fJ3ktIcMwgzJW36rHFg08/VdN/TN/UQ0y5aj46z
uLlEDEbK2CZANb/U9K0O1fkfpfaB76jXSJIVVaUpbqMJOpJeGMcmIj2QeIts4Xi1jbZtey6ZY+8M
0X5n3BzroVjGxHPW7gykk0vU54LC3zdgfsRQ6S8uIZab3VdkIdNK8BDv2T2tsnBl3V9YBcNKXZOO
iHwnBIH7/y+PAtT1NVA/p4NeptG+CzVVt1djNdmBtkOLx6H73QcsnAjGhoVwZJYt+pCmAkh8W+ai
N1jdt8BxjISzj1cZY7yJMkSYBuCId8vo/sekRZ2BCedBGShs2ch1nEM8onAgsL4s8IV57elHQY60
XsZKde2gyz0X3Oid3W9chWRyWETxcdBZz6EfjR6Gb2tgvJeBpq38HlGLnlxA1l7L72OmhM7LgMW+
QmtPJZmSgmhda4QEto2RxbmPCbVmG4hjSXxyQfvtXQmakHPjdcVo0AD8lBIChXuQnpsh+qinqCEb
lqTDI6dLQQYnznIalfePDes9zVVJwWQsH0yn+7egTdvwqb2F6MXwXpZswznnY0pn9Zb8rPfHmzpG
Mn0fkHVjYvE7jle57F3hkNDUurNhUf7H1UH1lHA8pKsrgLoZrs5vPt52RuGMvqeQ5JwbAbqTZma+
dE672Mhq2MYxUd15NUK7tVA1Bl04Ym3I5KOSCLkuoomgtdVorLtd4Fx3uIsbGRUzHvCTxfW7UPcE
A1XPfSqbw2eEe4B7hqFTvtBJX6KxJuTRXz5xPB+Bn/yXjUxUP8XSsNtC07nNYL3Vht0lXj4z2wj1
TqOrhu/ZF40t5EyHhYIXTJ1LarBWaDy2vN0ACWKGzzFXW9OP1pbVKTMMmFrqnCinpAX8SgXL0PN2
sna3a1V/ExchTJHJIGeSBEg3e7q5E1GJlx1ElQQD1bWUa+YsIiiva8CAVuT8US3S4SRZAvoSLB0z
rXRcVk7hrs3JmByF8QVCcmvtc1j40o0k3XvCpUwhK4nmMiZ38DUZ/LNOs6FO9twn0BGjo3ZKmTsx
cSExCUWbwKwyhG0Sej4E8nScTITW5oYZ/JuUdS3IENow3Lii4MITnMUn56G1KNJV2fiYfKXjSUbj
d0Jyz+5NySb04FWwDY+B4XpmKDzosGS8VBO/L6D9H/UBWYzuvFWXjrMm+AEF0iEHEVeaNBNi1GBG
caWmUd71zrUeEeEPM5hgUS7yHD+VJNV5oIQZoGDCUE5yehpfwMqb2o4HhDHDilQvAcyOGPEwEZSz
X6a/jX1XLM0vK4mY0tozWOyI9viZX4p8bLNo5CtoWfoE1PZuMS54cw9zavRbIl0Y6gY046gfhuFl
KACNh3oYilVUvMBTCirfrGgguGtEYZTD/woiaot2hb1Cbl7vadGYK6YokJYQ+IuFpqJG+uPW35Mq
vYLQgQ0kxbGtjZep4Z/VaG5PEYzQmBPrA2szpIkDl1J8Ad81ZYcE4yPsKBJWdK7cvqf3PD53tnQg
W780lz2IGLtygReEw/8azxhl1zyZJGQUNuDSeqlhjE3saOGUvtENhizRO+XBRahz04WH8WvXCPHt
hKSQHxbgRnCweamyw9tIUIva+gHDh5nLzHZrdVAK1sAZ6RvV4Dvq+5hFv9CTHBGllVt1ESEVhfZi
XvWfWS0VBb4iNGly+jY4+tZlXz2NvxG8AU5G0Yf76mSxTogJbpM/YrIwU1/v6x6z9PEf2vYintDR
e6OaLQub2S5M5EokZEJ07oqlCg0lzs72mQVtNiBIFZlkK7pELEqa5Au8RTlbgSbjWbmFnCVxeanW
smeQjRdIICMrlGZgFjoqclC+V6UCGmEveBAzM3lesd+2Dpl0loXWqNmHwRY4rwW2of/H1I0PfRo1
+RO5oujirBAaNOsXsTeuD+95tANAGwUtyqjQOym90zxatggEepj5YvffqTcxpXHbQ2HNfGZ2SB5H
6tyu8uCZ2sFize237kAAVKH7JUjZ6/YKjYEeJoeauSn5DiUgp0lO8X1oCHCr3idW8ugi5jrTiLDi
KuLB0SGoksllw+UxO8zetjwMRC3+UVcGs4JDkw2TkjCYCvZddMyKRd/5WisOCYnnIA1sPScEVUVO
ZoSEQChSGZg9xk7qjA7StWwHdaiTCsicT+j1EbxgrMN7m5plwgCnZkP1tD8aknHYm+igQsuOjpjC
brLQGIo8xDq3tXNZT/NjZhp3QB0Sh2NumooUGoO/O/thqmdsLyLlM6U2m6v0jauVgHlP7S5q2sKr
MRHtW6yRqHySd4v7k8O+96g0FupthzxFqwfJX2riFknySBXp6tw4qga38kjC3eEfWKxx4PqHjEbz
AAatfp+p8xYc5tud+28eJPEO1ooMqntUQmLmfdPZ8sCoqrB5+mr8f8lec0EJ6OCTVIvOJtgQUFrR
CzpgZa0leDSuduXyVGW3e3aLmTHOT0YzgJfV6KxEj/TWTUh6VrgbyxNajsRgeE7znp8pe3GRmOQD
noYUCedWpvTvha9Z+PO3IXM67MWrCW7iqIoEdeLS3ZC1lTKvvF//ghodVA1IjkV0guVYoJ01rhiN
nf0B7wtpJlbMbNsPtFET5FfNLE7a0xF7Sst3NkYRmLXc5Q0YBzckW6oWOGgN/tU4M60e+NBg4DZX
m1y407T1Xw4J9N+VBxh8x91C0Uve2DqMnAVM6dhM3Z378TrWanCcwnRbCo9ja0Gc1/M4Pu3przda
1DcLTPmUN15UNLyId7Sevl5b5JsAA5xVLVUgYGDLh+uAowjlOKwvb2+rktH9WM60S68C0uw/LfDU
8cRpEdpOSq2cJYMmW287HkKyGPxiMmGAO8oXRw2O36TY7SVPjbxAWQLRGI6c7GyVXnZ6zzdZ5oCP
MVbxGCLdTnsSdCEkyzbyoQoivsom4FNvLNkJIyA2dcL93bcX1/jvqjpcQb6BItKnWACAEj9oQ5XL
VCMkZs8ZKdBt5xnW1WUkdAe0W7MkW4e9n681wXzrd1ch+mN1KSRUNgekxIcAmJe8n7xadbgXyHgh
8hNxmS82SQtkEBMPGJhwQMli4wsn8E7x2vdbX6aBku/gVy6qwQIokHk//VKiyLaquTW708mGdpaI
nJWu0PfkQUCz/OX2cYwlSdYg3Naskjumb/Xtc9Txnfi5TaVydJvK7muN/1OGV+uscpbCgFJq4afk
JBqfs9Afm3RiKC4QgVpq3utR9jgVaMI2JE/QRaSPsrp4j/9ddIKBvsvSpQHAvvlt4mjUwVWzBL2h
nLF0pgqu6noj4dwLngdNjTMrSjsoRdVDAFYOozPxEW9lwfSbqHe5lDSlGXIzIFNUTNT+Mx4DukgY
Ef99/717vrqEBjNnMeKn8liE0N0HtxEJbxGmdFAWbDh4nhYvBCkJAN8zCKZRhOg/seRJu+2fRpIT
eJtwI7U0wsynE9OGtamFAIoF6neDvGpe8Xuq3MeBzW5AuaCNERE+0uiHuOqtbmHFZz1CTf6dILF1
7boX7T1kTvBYaHVtXae+ogaHcx/S4LHvugf/tYWXwYcYtHZQDwFxsEsdg+3cUmDmqg4A4cAa949i
/4Tyjgv4CiwrbXMahdRkD7E8+V8PL2jPkbfEAQtqbFX183VZkhdeymNcfkD3OxFcnOnDF62vwhlN
rBIJUuGvQJugWqdwD6dxZXKx7V/yC71oLuasQmvR7g8g/sHnvQikyFsQRjyXT3zHLPFRX57ZkYqM
BypFQfwp6MRjXFfB/YIoie+7Xx+gBP7xLG3UVSu3ECS3bEOSKuAKpFTi/KCooZeJouXpkvuBa17y
hirjLOFOXnTD+tBIWXE2RErO8yvIROFHoU3uCkCjYyri4sgfGxltfZq0bX+7Jhy+CJY36AZVTP0X
/2PMaSPDsj9jPQ9oydZaZrwnhibw4I+z8QNl0A5a5KdY37QFedJ+WM28og+oemACDPb8b6FDyluZ
bt3kkypa5Y8+kBwfFBNyr0Tbo/TJAi/YfjbrLPsGdd6Crm0udeJiKBM2PbpYfyZVfCM+wtAE2DiD
vMqT3HoMI6rbaeJdzOspY5PU3TfOaWdvRJdAJs0Bzc9VMFApDYzdfKy0/ncxvc2+yQTJOM+Siy9M
dvNLjuO4pUjI/znsiwZ6GvYXUvKL946+3x1ptofR740jyN4n6+NU/13k5pWmon+UxUl/y2ysv3lI
U/yzoM7xjp+adSmZG0UW0BeoM7FefCJRRfLDeDA9rkiPlWpcftPiER7rFl/XYNSFQL7d5DP/9R/y
de4P+MhV0ElVPNWs//mAeVycRvaEQy5yq8luub+ZKW+bqDAeUxJH8le+bjrX/y43v25Xy0NKkAOj
/Fq5c3xKOd2Cv9aHXkirHXf69Gm54WupMQCIXOraUtbd6nv+DlMjPMtLqy3lCayGIo5qAQo6MR6x
N6sSkX8by9erpfx4T+ZA5FnCSImn/mnAANbxm4qMX8P96UJ55GVNeVgiRpn1iQzjgVgBEPzIGXF1
u2sHf2u9hAZXhNJ4hYCbYT67Yh3wwc0U2Vc/r+y8eu3jz6koDYEgtPM62/rdltD8S45DjBkZoqx7
NT6T0zBIUhBxpRSZSDTVQhRCtEgx8WGUZAYT2Z+7/oJftDWuZD1QIao/w8uQBvNW3U90Xqm2Rgh9
iGVYhMTbEEp7W4c6TzBoPjMwXX7IwoO+xJgOCUmPWFqDAPeTYENKXsPqwjWQil1yic1s437rS53F
i/qg/pTGsygI8dQI6/Chto8hdjIKTePrRsFHuMJWsOfAN6pdwtAMcVgwTAV2LatpINQVIfDa4frd
1QzNZRM6Jh35aoyrV63STmHLIry1k2ctLHVYxGeWMkgfrJ/EerUL0Ze810jhhcm125Lu/5Z4+MP4
WDLO8GTbAgure93hPs2Bx438LnZQfVGtfxheNzAqWQXMgSF2n1Q8hbmREm5LX7UV3+AJup2dgwh5
UWLI7pJVEJYfEBoCflFkF1v80aETX3AYqPj8FIMji6vz20JGrWeJsmmMIwmKP7L4GXNgoBik6Wnt
JHtNI8vSmB4UuxQErdY85Hpx3Xe3DE+muRdoevUmB6iPEyVTgK0xPvgO/3T28Ln48NgvRVHWA+tP
1loB2vh95AabIx+v/qj+HK1qejKYXLajOD55HDHxbuUOOoI4rbZtMi0xP1TiyL1FidWdyRwwz8wE
JBTjfozLEF0KiD2ll55ydzRY9W/9MECfwnSoazBwNXyY1M/U/GMaHLT5Xl+Gh3c6NFmhDph4K6bq
2WxqqAF4L6SPvYBfwSItquTqpFeS5WXz4pFOGa9+Cl7GqbcuyN+px+XfUPxgXF837FPqf/X2kTPg
T3OAPUyS4oaAJ8DzAs7k3xXuLqmSF82IoztDsNgPKVVz7E2LrlWvl2EGhk+LlF4xVFqvQLNBMruB
o77Vwl2YzVAFG2o6ygHeXqke9cxG8rYYHY78SE0kD89zNiEv5vtoUjFkTXHSWfzh+WB0pcyErBsI
5NZG6GTkG6nYRgYB35jdRvBYqoqKRF8tqj1cFhduiTmiU6qPUIkaG1yYIq9IbbP+4g1pMN/Jjdxk
3cJXxiq08wWUbWJ0dPrIIG3jIamQRffHt+FxqDbYgVSr4scCS19odLKJC8ul/XhZUlLVNlv9D1Yd
RbbfpJoTpYyupsT750UMEzu9ty+bTWBrFj2QrFWB2CppslsbcfHwyn9Ob05Pie1ycAqUfjOYlOx6
1WVWYbfCY+Fwc8dEqxTF6bIXtcAvqmCCZYnfAfhJz4f8NAe6pulNZzAGebgnjBr6YgA9FOQ1KeNf
GbvZkgdn77NH9VsE624iAtG/11pvIjVWZHWEzMTBmjK9nigaJc6LHQbc6QS5a2SXmb39nwmdWCvb
c7xgU0wBMB4mBooNkOnhVOz5gk5hg1awVrypmepqJpYz8j+QVejpBiB4X3tVVydym6RhktD4zdeQ
o2H4br27cXbQ0hx7nYuBSw2C8vg68dyS2jHGTPQdpU9iW/gWHy6ChZh19s0rfYMokBwjRhLXp/kU
MLn3BQzvEQ+0rVyXRhflHA69af3XVuYfj/wNqLRuZZmOfjofd3NtKF3mGT2KGwdaLFpfqY4OpJ8R
VYAFIV3BJwZfaUWCiOnuFfXqLtiTujdPy1ujfkw1bmf1tS8xL18g+TGcMUpjcGC8MAbNtGj/NlLG
yJDkEqQ4wpP0xTIyNI/u92GH6PBoksT4IKO1BnDRPSkhUnSWMGAZM8OjpY25QNPQr+0yKDsVDLZ9
QBhWbqmPKctKG9uMSIPDaGAVtDZ9i9j8IVTJXhTR6fizOJzeg5nGSc5QFm1Ff6pADJK9OgFhOZcr
9pOQq/6qdH5tzvRmzPLxMrtgbbQIkIIAb7J1Nt/saD2CMUA3dvYcBbTn+w0hYTk/WixZjT/fo704
JgtIOouaA5QmLuHu9zF6r92wPYUpoW8NjdVBWKAVYD+LLG8a2tT8cmCnQb89w5fzNAb7nNPb+Yqj
uqoXlNI9aQPS8yjM5ZEoSu5fAPshTb1hpOUtjaIThJHQlTBDKQX/2gD3GlXyqLDej7FKSCBW9NXv
I0bpsWqA+ioGNBkwmjH+ulv2dqpo2l0cp1kBiSXcEWy3RZjXGvG0TGC84xAkSgNsrn9ezwAgiyVS
a4yOSvNvbtSkze1jV8dCzDEYIdgKuM8Hx7wVVKMmZR/be1qavxrxjcXswxkdNW6E4wybMKIwFgaa
yyol+hyxi1VvG9zDYcBUAjTssr+q42dyP3E6hzT5lwzFhqIOvAmTa0LDMb7lVEzbV/kNMZDgVH4J
rsfx8mNnt9dEnJxxnLIhTqApdR3XUnEe0Q5HAmaDuxnk0hk+U9XRNsuf/1VbRjJXpE0Je+ARMhKG
9fabbXHu/wW4GXHw9ZZBLzUWqV1/4b6jtkuxHP997X1147PB/ERySrE6LMVqZo6v0WajXKBzUD5w
tjKcXqa1U8LcxaS0mZGRM8j6/EtOLp8BbLkq5zXxPkyyUorJV68F+F3UOXAi9IEEznm05GmQq3I/
4vqskWhEKVjgmiEufCSxdWSTYZhzkTDkPMiuA3do7zrQ5n1DvxxIyW5JIfWmnoCbtrewwDqBOHdl
bSIv6XLegVkN5X0k8r2UGk/77KqANurdbGWg8hmBJUea1pKoUXehwWV4xMt0z5BKnL/vrFrYPaU8
6HrOnzHjwrPmHy8SH8cU2lH2YOI8eIBUbG8gXLa3pN54inHgxA9cat0Sie86G9XYwArqEhY/cyzh
v8vCH+u2TDYmYnkk0cbvvLJBCixyc8PlUKQzMqbn8fco3m0uFjTCbZoUkaocUD2ijeP+E83+v33w
pZSWiECuTj72n4sBrcgfIhfIt5det42U7WKcjdG9vH5bU/rqh60RIWdLhmRCPUHfI5WQA8AId4Jp
MZGQbUUEgqGrOEVdMtC0ly9AF1IuG5kKJYYzEHKS9lRGoETiDYpjXXWOiYkZSSlkic4W2IM+B9yw
v+d3qWq3tC9F8BRpDaxtYAhQhLhlX4GY5sMmNNwHxljkqHnld4B7wl31MasZ1yT9WKZUbtp2qEzN
dOFsPrjs4JCWh5e446fv8qSM1lyoVvxxALkKlAwzE4uiucc2BGPz40tb5Okts+S5hME+6rLKIMZC
NXP5akRYEyrmO8jNEvikOuPG1Ov9LtvCnWt0eTnjCoXNGQHJkuqEE+QpQZLRtOTKTNp0+zVUffZY
7lzZ6BbRWWClPs5o9DwuVKPWansBRzKRzK+ll2itTD2VGNOT+IGHjxgtgKHbMAebZKpaCyEO/KBD
qHkM4EnTcIf9pi9pETQn6bL4s11j7aGiem+YYsMtuSVI5ove+/uLWzgYi+H0xUwF3Tt7Vwu51rDX
fqCV0gbsQwgjvyohf72rq4q+Z6YgKidBKof7ztnasjcYQjZH47hGNSjV3rm9cEBiQj4MX5umr6ki
/BNeqkVrKUE2kLy0bHb13PNhOWGBKWB09s1ZpCnUEEA1VuQmd3pew3UNfOFIvOelo17dvd3gUPG/
U6Un5L3gwYPccshncBDbtQ0YrRDlFGyqCv8kaashoXPY2OalBkxUjslQvaJCDduwcRGJrgKJ86sK
q1jW8UuY0qInEANINz1KR/bFiGhGKgV5YUMfFf+XAvBrVCQXOie9ylJMKtJW5F/0XZ0twGr9IPAD
IKca97IoEUu+b98VjBr6HK5t9nslvHtAcK1It2ELCPV2mbS18fo70HN1dtY6BYPZteTpjDqr5S2M
1gHcSORLw86SURt6ztfSQMpIR6chQEir85q56af/ZqQW6zjuA3Lavdo+FmragDOkWOE2CLfc5xoW
Q6dkmPyWCEXotthc5q66Gd+IWGbZ0IC0yuZ/4tSsKh1fYVLE6FkzSWeSBtgNigiO29brE0ExFBrQ
xmVQAUbOhkmns/sijdjxRMGnnCFajLrw1YGdfVeNisYkbkOnLDumnhL1exoBkK2ZeJBBqtc3uHKn
yhBTIHDKdHsU+tqHk/+K+Y7PGzcjkbP5WzUzzX13qRGp0MfN32Uy4Es1NT36RaSxNtdMb8pthJvK
XI7l5S2QHkAmHVHcJ+eC1hcFBkrMWIMvp23I2nFoGOdJwDZ4LvIdU5a3Tb+vwzz9ejwI72oHMoHg
Rbuz+mKtm1+jxx02ukU4rJ6cPhSZM7zq30nKIze/W2k4cgs4Vbu4BA0Eh4RUIsStvegSIUERsR4e
cXLGFd4+QsLOhYNHNIbOf6Lnd7lotq7JBKr1uNAgPoPduR5f0tpGik6P+q2nVXBJoK/edieDLjwN
wwZXC8JaftXao7TWr0AmGKFHAo8A/qsmaXNtHnrAu5G2A5oU/WI+FmCrpell6vM1lbYAnYhqYqOR
TVFWpsDDVjwpJiRspiNnSJjN1VdG+qgYdqZ8zOl0BBnyamk9crM1hTSTHTMnpQ1bXSZnYbfIHthA
hXxk1OfVA/EKY82cXILaCWFhfXhVj4MRMlZhFp3bF71Z9QBykixt0w/lgqCF40+ndRz/1wDZVqol
fMNQ3/X5REnsZAm9LzBFP55731MC/ebgj+43uPFbEqs6mguMD7q84XS9ztngi2QWWwUyUnw3wI0c
xhZhVe62d9/d13g18/xrQ9QcB3oE4LI1Uai3ytdVB9MwDanm4TdRBIlC7UCaiGg7wO65XAdhXeDy
dBuDciS/ru1ziM6Y5Y/iAqQsV95iHblaI/hqfVW5IUPtAYyFOf6FwKsm8scqbi55RFgWZDc07pRQ
hFlgDcV4V+zjI4JJqnbx3Fiu18MJzhXngc7AQnqIOStB1fx5p+UmHJCNNzS00FZaxWO/qGIGaGz4
Q5IRp7B4G88JbaJUlTNuvgnjABT3P5Dgkf/zvwhZvRvQeQvHhv5O10ye5VK1qmRxgycccL2RXAN8
EeUCmByzwME/sOJMkeQAsjFh5BOFtAYA7I54iqVv6Ba6YVCXNG0oSqi60cheg9CzJ2MboM8/r4Yt
UE3QwgEvN4RdAJ/M8EZyKDHd+mMue4TnxJ5H8ImdCjjyWDfFw+gMQO5LJctvcKlA7aROtxuXyhmv
AZgxlpYgGuTc0s1iVspzKbCgq49zKZLc5f/E8EbQhzbviJBw2/g6axqlcf/pYzQS7sefm8DK8bbh
doO5ZCcGCMp+4ehDQvGwBinO78z0xVNwu8+PHNknZh981WhguhQ+GDklKUX2boIlUZ36UMH0oYBk
OETmYaK5E9enzXJrE14nynhr2txcHIo4kJc4T3tBjdn114wk3yedpIWPKT2chgFTfoFrOz5etMHN
7cyrY7iNZi3koN+2gCD15BZcwiWoYZJc6Cra3W5xxmhzu3z3TWLMlDmb5JSox4ggRfDGOHhhhz0L
JyPu7lHAhHFDFd5ibu6cCU4xSDcuw2GXq6gqW77HoH+Gtv2HOPakvYDX6jt7LwGugzH57p5ft6/Z
RZhYZl9Rkmxpe9PrELO+yry/AcDSV08tVKqGgF5QJ4wtCU3rQACVM8TvCtyXelvuLUIcOirqhT4a
C8hq2jLwlIowQBwnEjFP2tYdaVEDRrQFiOaF437bWVbDgq5qjnfW7rLDGyqV3zedyoH5H/FdHINa
AA75Ljeymjzc1cipm26/VSRaIkZWoK1sf5Xpji2c0qdO0lydXwqGzW6yL4jg3+mWmTzcFekXEWyK
ub9LFEzMjcxq4xhrUxhjElmTL0RyCOKty+FMXaIBXxvi107NyWB/kHkkO1TtX49o6mI5i838iljO
hQ5b1ARsOBC+3uFE2Cg2mCzOo7reD0x/Q1jxweKK8zgCSPsUHmVLTSD9kVzBr4mlIq6cKTewScvp
nblFbv6FvfSj8c57V99CgOyzmenYqokz1baek/sFRyh6m3HKACBXMJxEax4l54NYpTfdcujHIKrt
eQX3rb8OXTEIAR/bEYVLIUU8glQHgVIZtSzF5TW3qtqVDSHwLjmUduE285nY4sqkJFDzEr/WbQkt
XU3hAcqJeaMt4B/UtXiPphXvlb4TrP2YF5QOhcmYbsl3aYpQwoSweHZZjfHeddzZrcFYY7/JpOdB
p6rYu9aUWXgwCOG/VEOlskx7qWvhxJQ+X0bvYqz+Lr9sJfAu8xlLFvEMrbkmGvpdBYRTYtDPS8X2
6lskfiwaZk1CsojL+UOkTqUWA7/AKtfJvEYJi55aF11slS+cIY9AgPujnnHvQH2+UEhvz9KsdCqm
ZRN69ulWFOOY5R01e3B+7mNBr0gsphdGEx4FEn4AjhfuCYUcxReA5H2Kqd5D4HAF48RNXnropj2G
Zo71iWD3qQLBIVyrPxzQuTaLs5ShHv9Cl/qtf6TXk0HC/oTLNF6s3ENwFG5Fu88QlaVPZEoj/YGw
SxBUwce3nqQ/drklmVsDCpID0Mfyahf04obbRIpCPPH959vCpDPFPgw0Ak+JaCRXQg/eh0av4vB8
ifXG140fa0E9E0hO/hv1SUF6kgLw2qWobbAwHthzh37uVvlRDqDTR1sbQXPsDwjLMeCaPho3o4YI
+YB8tOtUmowB7JcFhMMwQbCA8eMZyScY6jdLRTXnEf6p/AgRXgAO51bTPX4l+amYwo6HoOe/tcdM
T3k2gVNy0k8P4R1Z4gC3MZzc9yQWfHgmbf9d8dH49AwVYsVVY8WrAPcxZ6l3N0oowoPFFpYnaWAN
as+POPTZiclVyDFPDTpyrCYZQsjYJHu0CEY8axgpWaDuJjRrq8KShRTw/4VF/HqsA/TkbHX3b6+F
pYXkfXEBeB6Eo9ICK8HonwLFaCAgffMvBsASA1PvpJ2iSDWw6a9CaCh7rTu2FHGeH/SwO7VnBHRn
8Sq0BZCU+DPXVeDJrp15+DsQVXdvhMYEaBGdOTuXc72Of/HkJChLNEb2IdZGPZLNqtMB9x+onKpu
zpH2DtE0WErzm8ojVWBJZ66NX9tWGcJ+w+eo/YMKstBQe+i1R8fYHJJv7asgKqIc8X0r40ZnOtGp
6i2iDRxP3skXZxZc6d/mLlCRvLT5/58qzsi7V6eALSULnpvbgdZTTM+bMMxaCwbhUZkO08nr4IS1
EpEvY8X6/y+/3KHiTF+YK/qQKfFqtlxDDm5RuXQhGtvjexX3WXV9DcD8eF5sKIZxliQqQB/zVeNf
abauQ+5EXXJbdrMNKpefcMdfngcSt9taudC9+mpl4uBQ6PydI71yKKP0CfXWl1ZNwmtLg0JuSA8U
MHrqEtA4jVVLCu6c9PmbOwoaRSyXE1Mo0rbYSSCEVSsBypHsd9qxJWD+CQbM+QNJb3j2sfTGafJb
zvmKjiPkIRG0ZiBflmNhx6sUAgvhfYIdBd4y4HCXBpffQxsZ7hCFe52kO4jQCWzp2Hj4HKzk0cRi
vJatoLOxXaVMjimxsP9fHeemDRJ3AuSDobyJ0kC2eMt2Dw9KY3gfK8KEdm69Fz6CX0KFeIksrjso
BiD2z924RdyPthrHqZhObBSSA/lLhj+65aQVk9s1hn5CPCjncMi1g2uUTXibEnNvSbDjZMRKmaAw
lrG5TvGzwOp5kMc4aumBrUJHdeqEaS+PQMbmAWGui2asTquU/G2vG4EXcbzRtqRtGVk7wvJsQSZC
mWXPPQ8+G2rPlQKLagL3ggmsP/X3kCoS53lMFk0Gv9gR8b66uXR8mkWGo8b94NnO75JesMW24vN/
IIERzljbu7qEpqvP7omgq63VLwVb7zrWrIvHdsVrCmgH/EKPL948UEcQOTL3Tnx9KYyjCZ8YrXQP
dTIkxDGdWuohjZ7sBndxFJ0jF9BRgyTtXLTAM7mmgPR16GuazwztCeTcMDQJVjJF5hyVc9yWYn3Y
tDtn4AkkzTeUut80YUVxWm1EeX7s2+TVIGkXTiNwVcESY9d+D4Hh9T53DonV7nXN3VyWBUmhtJRO
u2dSt/d/kdQpRzEfAP1RziGOWmkyr0EBXmOa0QFOwkqXTABgNmyGmguVYm4lFZHZfHFyx7X+iaSj
zHoUKAFJSeF4DR6+qajn82Blc9/e85Z+j3X58NWvWFniJ9YYs4uOnP+fxOBHAH2NJb55j573IxaF
k86+fI0pGDtjqtXh83qlOTmOm2AfG8+BzvKcKNW3PoedWsWx/Z81MpVkpZr4GcYZJ4opLqvrR+yb
PDzXZFnDVrzIHq78fGQYKLPaN1SRBq8DBc4uAvmpS/nzK/q6LmKFZ8QJXIEN1TxCSbqM8GJAKWsz
GrcejZTTQinDP8Zh+ltGu/iuRHA1cJbb2z8/Szscvf69mMgUs0Pq4aOXJOYSbbIkIneydD/EqgLe
QQmVc5Sod9vnObIL++s3mGO6qwnq/lFgCNfyiUQCPwANVjMtd7dkn1BsfwRB16n4sN3lvgZRhnPn
imVgNWLs08FSJF/HUwwgGsXlsWuV7FKIF5qPgvE1fq4rcVikfsK9KfAFn1AFSkX2CjYmkU7fj0gZ
IjPr2sD1Fmmxd+LednPJWqV6r5SetkxL2eXN1R65D9HXm/DKGRqV1+Vw+mWjVVzlu/RqTTmGwBwJ
8hXgNrFWle0+ZrQXD9iCUI3SuAjPv1OR3GeQmnw7v4a4xmZhO3uEcAzP7C8aQ9fqxYDDFNH7Qpcj
vFh/z5anJMmaCG7xQHtwzcx0RolcjtVZZOBqE9VoY0rFeOywlYH1ES5BWh2/oneDM6eDp5UZyMUN
ujjKrQaBjtiEr0pYoxXegGUY2IthvuN02NyqT5i54d07PdugWscxbVtGKCAZwaCm8oqOBuMd1G4R
sSibDEA2JqtfwVgQL4+hCar5htPLV6PAKn7AmStDJC1vCVIaTovsHNEO9APmSiiucFCaEf4MB4lf
v13o+NmFU8hdA42xOq6rrSoXDkIgQy7aLDul9iOmiVuOvspaGoef4WATYa/94QqYiL1u2hjF86SQ
e+s1xSYNbV+O5GQs6jSVhr9iYT7Z6CfZMx3WWV8Ogn+gfYTjUYqHH1VwgU/xY430Fy062snbHkGe
EBTsXdZ/Dxgh3iRy806QMMck7pVsL1tHmNBcAe0CZ/4eLmYTFvZosJPZEj2C/cR7L09x5Dtvk+eM
pySDAf3GAdESAUEIxEXg9s0x/ATAYXDDEfBUK+diUow3DQU8SCjo3S7hmoTXKSGDhf/VnC2YTDZ1
wzaWh8Dj0w8HHcGxmUubknST8CsGU16QPQHKwmC+DVGQNDXoX0LR+8mEis3lSPtpVb3x/86PdWdI
pEPdUJGgE2nPfMoSnjhjUmqudG87EaVqDoT1WkaF1BhM/BzpaA+YU8yb38ZZ8tT2+v1ZQW8I8W56
ZYhlR0cHj9Hz4qSuIW0VIp0ibVgTXvbcjQuaFnSYxZXs1mTLtm7oHXHJ0b4I+SMuyPNLkH/Y3Sg9
KGa+Ttea5cPBPR/NBFTYQlNu9lk9bSVxYcElQ/SMytLGfEM6U8n9t+kqGEk+1glsEv3BVcNOZ6Ay
G/oZ9zExpaqOIWZgBnUxOgnPXe4QtJgDFXWuaqEHaeacD8PHx7xWfAmWSm9TfDGGaIJMbLXjCLtA
86tqtmQiTwZH//8loTH0uqXAuPKuBuhezLxKFEliPeOH7WLcwIkTCs4OUfjox0MP3AY+0OX3qPAU
t2gT9rPYbY69GYmmVxO5ttfS1W+DwPmzYkWeWe+5vE1JsooqoE6T2HXydHipchg02YNLJk8p9AJ9
4FILVUaIjfkTwiGbKpfeu/QNnefkZRiTEKIn9fIW8Sq8LEAIYyFyVk4307Mi/UZ3oNoxQBnPY23P
uDQ/pdWtEGiR4wKmA8310Df5e+l6/OLoDsyyTg28FPV+7Ch9mVfuEOHVCqLE+rUQKgdVBgOWfPPp
346lLJ2YqkNCyJCJhFOey64slJ/VqDAjkrRuMUpy9fkg8p0wNmn6m9gH1ku4ZVzNjDZsU2mfoZHa
DzUPe3TUMmHaNh0ZWU+xo/Gao980r5IVzoUyCsLiuoesdvNYobQox5GBDZ9Gql1FukUJFNLmEejq
IXSABCuV1o3UB4YZD6U/DR25hwLPxj+08NFXNXh6IRpJB+cTAx9e04/3gLw99lz/5Qg2jjCbluLM
Q1a4P0Xy1M6kND+m/Lo2kk1SWcwCFL87/WohIF0klItrTb/S3+TPM4c/RRYeDur13FtYtV+AAAs6
tqM53QCtXFaG3ikJ+eCqFJVYHrLIY7YeBwpLZHsVyrgmcE7iukqZfQrzMWCH7lC12zT6WoTMZ5HH
H7Sx8QtKny8oNcEqB0dgVYO6egwGRGd3bcaMID4RxZ/fZSw9htT6APhgfJ/gH4Pn29AKfHjyRyo1
ll3ESGelOSK9UuDPVKkzE4vcjCA60Pbbopn7dNGaEyTU6BQGJMvBSj9aMsSO5MemaEFg+DjerU1w
1brLi5QKoLEahNwu8Bl2xT0Q1fSr7+hbVmkEMQ+ZjTp7dHWbGNYotcSNmSJbyn8Cc9TNyajrpBv7
OIcK0jcVjaal1ZeWwuZ5aYhayW9INPU1gHB30q3/t47cQ6Pqtyx9jfdtHXn3In68A/f1vI1vvxCY
vWHhjCZPtDFBhJdYZ2yPf9mR8EMJM02Eep0MgdO5OiKCFr+XyU736CMBRT3ahgkGjBwIaT35F9av
v2ETVeanUH6Hn0AUNpHNtGfNzfa66gxWsmUDXfLMGXembsNgD52ihpKnWZLT2LHTiHsdw4LPpuFh
0DaQG6Px18vMPU0A0IPjH681g2lmLWqJvtCSqBHNd5LQLTHbM1ONpT4q+TvStLhSJ/+a26nWegfG
YTsaJ8ch+6wwfC6h4pfw7xOfjnb3fiDmuub4qodxSFySpNT/aRfW0PNRQVraHb1RwRVwMpkkNxzF
DLa2IZByK82XMpPD4m9DiYRFAX2HzNjoz0hgk6bV7RtWcQWanU9Sk1oo9wk/rqMfxtWg+pEtS7PT
+llghc8miQiTu0/JPL8EIL4kE6NpNRdJvEH21bxssfdewx7A+B2KDhpAxlKjXpHlXNkhuToJ/Pgk
qmfMtNwdZSUUPaBHX8AB+Av2NFJ4oJLPONYhgM9/2N4Pf+WJFfghDncKAfHmDu6D/FymkovoLUP9
KV0RlE/G1H/MGumOizOHBcAf6aTzf7Auc4CHkLX44sLWkwNFnf6JSPmboylAJ3q3c7mJvqE/kyU4
RyQQMQyhdGwm5KYrZnUwErSEGzACl1kmps0TzF1mtNoz2ddKhmb1NeoNFkS7yVIiwsF7MjGVybYG
FMrxSRYLutvmITlO+MPEOo08IAUZflq4v5ofo78iOzXd+9oHcY36W8iR4MOKOBxMz4uX7mmufAp2
hffMB1xqC5vv1KLVHaeWf/OecKERJpnrkLNeIexJmKFIhxJst44UDeKrDBLWhgGx3OhflUY0aASE
f7rjQ/A/DZ3mPVoA56BwKOq6qc5TZiZHeH8ZDYCigbfpTMcvEg5r/8OrPHC6M8qGmI2pkC69OFlu
gPfBuzfVQXM/4y6HoGJQbRIKC1F4VbZm85F+lS7slUSIeic+06hDPvsgmM4bCa6C9ke9+02qPYGa
RXq5ofLxf/S3FAyQzbCPwFdLuqHrv3AdeStA68JaOBxLALLJlTHeAJ17FmEsrWZzEzsdt4zsKDzu
XcaEaXjFtNqKVAbGqZwcsG/f5rpe/Vgwe9DXE8vdGPpTkgKpWXzOACe8Frtaj5IAHT+eHa2VyxYZ
xPVxskyyz3nzj8H8ghLJUSjP10swbfSSbJDJJYdViGrdEUU6ytIVkA8MpADJSm4QSjEdXdh9YKi5
m1Nj2GNyFrNFMOv5YumZsEQ1vu2SbNboURYGhZgFwXIO7VHpx1ij6qSMe3s/rlLjTBMvn5Qyt5DL
uPB5JzTIOTPAvkGhapHbEdsHDWwNfodeCIMWWKDQPtnO9TYVYfQOq3N/opcEItjE1DtNff7VvNcL
fHZCCFJC2AhfxWVU1u6mbxbe+BnbfSxDL76/7y4Y9FG8i4sDyGvLRBWmykdsRlmMve0Nu8bQYVdO
SuU057gjycFYG2IY0CfoSLr55iolYO8YEju++yXdcLuC/js/hzKpoy5RxPavk8ejyfpzVy5cOGgN
mPV1oGitRFpP04e1Ka3hvYCdWh9EfFRxGQYafjk94vHjDvS7eujNNKy8Nge8iJDAKDn/HcPmxXG0
2UBYc/3IWLCTxyOxZLg9wmLqvZJJht3fbTzMOxXrQJbGCeT2+NiA2Fg9Zi9yteV2cBQHKxxmrZMx
emaf1ISbyC+rQfzyIMMqjbmNK5VCWDlC4QfjMJwrKp91A2N4Ne6kZVSlEHaxyz2TnbEwNUUdc8mF
GhyCiLozWJQCNHBLoKZpcX8FF6GsjNB8jv+YqJW4NDzcMm10BTEry8GMiFbJdamM6Hw9F2j5UlF5
S3qnVAkj679UEhlCwBm0Q9ete+3HkoE+52Ws2VPQ1fHmvtYxnITrpR2okvmkgX7mdmwhSrQrJyi3
aCImXwBh4l3u20AKSeS5VyRYaSocWrRLB4JHotZIk/u8XE6LXiE1prwG5yBTWCoNBVzOWV5ghH8x
0vivtb+7zy3XNAS1Bblixun5NM+zvLwB01liV3F4kQk/pUXIcNfgT03nHR2Rj2MHtiNevZCZUOQW
M37zahq2TrndqfVYQPWwdBqFdl5t+6/iW5prr0IlWFq74M/4y74BlMEXlLkTDvkKz6UOeRRkMT8q
rfjLMtuxq1o/SzCAUQXofh9hMs4PNuVq9TdqMvc2603Ll71q1/jhfBEn8xiAeXiFi3x84XjSqBGg
sU/GIsZ+6UacALrmqsDXSsAM3SZKm0CyYCt17oWSK8F/yPw4pJfzB37uypo2+WM5oQbWU0hwG0bP
aca3KVqKTfbT4tqRg2hQODDW/6FwEPLONPhkar2DZWAiwdzzwg1OuNOTtZuihCrB0hfEaRVlqXt8
R3t6w/Xi1pCjIwkGHwtItl+xFykdY2oBchAtlXg7q0t59877G2Clx2ED3SHucQM0fEOZoGiKEuBV
osvFaQDb6SnNIWyzwe2+85hsDR+Bm2EcHiAFJgYuyQq0Rp8t3RhEc+v9a06X+YVtMY4ke3Tw1m7r
/lrwsJ6QpCDi+EksO67YcMgqhfhyO5PbYsOlbu8u7oKodVrK10ZqUxWrQJCsSryMPCLlkRV69g/w
0chCwimPJKZDzWsTrdcvqocEENhn9bG5ii5bgczeGetZfqWPTT41C4S3rwLDkIx8rZyS0jvrpZ8H
dVWcgTl+nk6RWBKvxg2B8e/hVRS0/TVFlQ4PhV4Ga2UNTXCLo12LUiIVoB/ZTttfWgDaRkizePxG
xoKHSvk+01P0vRBKjvVD4ugL8YNFcd0eETFnL0s/9FwJsAymF83xpZe9RZPse/Y2X7nY2v4KAbV9
8RN3WOTnrYBIkU9uhhG5Bp25ta5d3XOVngI5dlYOVI4DXCDH9tOShEIxjeW6UvYjXEqJPO4gBiuK
EGGrh0A+eHElcbmOfgxkgypXkC48zITMlBANpX/yQmfdKBItUjd0zKT4wVvvlQyX+3XtVT4YwaZi
TeBMOpC7da9TjZ+1ZwAXn6q3IH2RXSqKY10P0Pehk8R07Qs2672TllmriAqha8MHId32VzzTRBGl
SyjXEIGI+LPfknwp4BTJePHxoxSUDZvAG/TAlqf3jvozpI0p2lALlIrpARJdB+C8zGYYTAa2nRVM
V/lUd7EUIpbWTLlrFpZjKDD+7HYnDDa/EX51yLNlS08lQGl/Mgp3rGbN+6r95Z7ybPNNTfY3kOcD
HQJaCI95wX3HFR1FpTCqS7EMSUtUAlzvGz4cZPXlXBHfm3xoXjUQbQixyg218YMP30ufsRo83GIf
DuPQKrwczi71VAzN7TxHl73nAt3Cb4NDirszM+ElmMcUFqKnyJBtQNSIloAGVaLe4JUUGc1UM6Bq
NngZYZtxlC4FiVq1v1hE0JUiVZtSoFbpxoALBdYyNFrb6sF6Hrde8Pcbk224ixUD7gY92amdepTa
lPJj599DtkHDln2SxcPcZhTeARGtTcQuNB63E+qZjvmXa/d7/0kmo0vQ+sRcxJDT37T+wYL62ORM
bTr2cthBSJd2PZbpfORSijRWEs95I9zqCrO6MMQIAovFXzTOaoBLQhUS1FZUwOoNbHzVR9nOhT2o
XMPUntq7+G80PU6oDGLq1LQeSVYfLMumnFJ3zGTqFaaIfpFmLXe72/Vs5CnfLwfMBUAiFIbvI0HQ
r0buQwgWLrxZOSPo/UoD8hwo5NKn6IKSJg38EAJctK5Kghde+qj4d2erTCjxJkKC61+mLStHOsQU
FqxWREhwarNhItUG8wVXhRolElkzKZnjtNEXpEsMUiiR9CIZW6GeR4reRL/akLqnpMhgt3/qlOxD
tuKHrgN2cYmUcfJpTNbbVUZNe63BSQUsx/RdoiEvdihn+8u//XKiyDH7lj/df9b69sZHTXg5umiJ
ZujN5A/0V+4ATg68w3Un6eBK42BzH77w/DmdHVok6FoFw1iUnrxggpRA7RFGFM8ptqAnQHnUeuJu
yTq+AbM2Fm6ewTlddcCdNJxv8x+hA9YHoQnfbFJ7NXgxBDfQqbvXpFopDqUtlmIBsRsFMASS6P1S
+BQDbJnEQCipRSNGISp41zZDK6pDc0PM81ZHsiml+gzx5CbV0fknK2LX0ZzAnSx+hRezuGdtIqwK
lFQK5J79vKaOzgVO+mWrLqyTdSnzDKFFDfS+LlHQiR/nmk8MRQBaQ2BCGXKyL3KyWuLGClM6zvts
PJbUvOIh/oZp8VAikCgAImWtMMoE428japrCKmiB+jcwiqkDhoWgbeq9dyfTpTw1e6qgKctCBoqo
j5xFp9SjkxC9RfqfMZGgELVkZXqxutR9RMolvOok4RWafjn9ixBqQF7CLbKLGmhF6fSMFydKMeTT
jpJXKf5w8ql9Pjar/D+IwHkA406CqCvNuLpfL4DsZOD4xw8zDKC/UbYBnR/gAPs/21n6VvJPKJ6Z
/xUR2OvympJBIHGvLk+N9aLvcDySTZLwy62WIHCbluSM7j1enRIJofMnIHv5SzxiskUIWywqYSzO
xvwJ3/6ty89Dd4UkVtG99kszz5B/eK2qp1+2Q1+8WGWlDT+BIbwPKsOK4HylZHHSQPS27tpMqaKS
u+aqNdeGhLV3A5yodg4cPE5UEU51lsWAGnjU7/SCdHJNoW4LYeWbint8uE9t1Yx2oHfpqAQjlCy8
B1DZ3aswlEyMx8MZ9ORSNSg4DmZCfKSrNzGWIQOghOTc7/9c+LxPSIRY+rohlcY2UJFbb4x3lJzx
+yvVoT4UMEROdwww4PfjEtgMpNF7kZpSrClBTd8vlISm7cax9A7QL9ab1QLIGWQVxCtlAYwS3Pu/
y3fDaBnzJnNBRJePFWtYlG4csIVUKX4LHKx4bKTs4RDBFknLMCCZ0Fn0z89x2s4UCT6GCMk8ur93
Zq2cib21E+Sc6dR0WkhXEhceV2gQ9hHFSmtXgQhsZ2z5bzel2nEFsHMcbbQqlekYR/ByaoTKJ7Y1
/+ZueqVr6Lx9gE/JYTTa3upQFMM1Oxv9MTjShIB7gmVcCgr4uNWaYPt1ThImR3QsJ+WV9Yz/6Z81
C9s1EYunU4cxMJDOHYWiurHafYGr2ylpqZ2m97MsxYCO2RdBXJzykbBC7LC5sPNlAhc8zUI+lk9T
sQr/g2dw3ymL9nkYnTdxF+sk10W4TUr+oQ4AH6qnkL6yooob6ttpmECnd0L5DnM/D3RXZg2mp06i
Nok98iI+0pSQ6bPpcAtj6lwvEMUoYR8rYM5fjoOAQBFVbTp7qXkG6BbzeYgMWXfv4UupTh7aji6p
Ts/ikAvFY0j5o2AnNtpU28ms+yH3RSsNZDY+3C8CCuUDa20r1rH2AKSrHLpuNvDtVF73Vbh80Z7K
Qn+OE+9eQdaeEhimP6Z5UOROOJ3G9sI2HkaCqTpQXa4yJ1jVi3B9h5fKpNBurgIE2b4sTTDd5jrD
AeKRSwxQLsj7eRLTYDycJUWk6Xl5Zf/lw4mywLtyb3wfEvVqA2e1zpi79JPEIZTZjg9xWTs/Fe8l
j1qPP4UDqJkzIqLJaQ1/oxzd8khP8E06BJDmu6V3Mzl85gQYHH/hYKxwuWjGWyxRMx7hFGU6SuKf
s1C5BasnQ3acolL5cYrySjMa3g3Bi9FXr7bTqkfpdbjmZAtAM2QY5qihqNDSsaANC1EdBhcNL4U6
sDOCFZh7sEnEsbALv/aVZxlIhoAOnJKO7EUIVDbGnK5X5s93M7h4RcE8aIq3PJJTeeecO5+nZxVP
9824Eeudr4bhAjcq/mp0GHHrfuVtidYmOnYgShS1wwg9oLqkTzfQT9rJWtyqhpUuOP7u6NRKoOr4
6Pt5lXpeBF06pr3hSMuwP+JD0K/p+kbnqZtQY+IcRcvdVsd9SmtQoy+/FGNmSw5IzhDXCpfvGLod
RtJDW3eHF5i28YEqvKKehF7AQSy8KpPW2AV3wRAY4+KKiq7SANqe+VYdRoXlArPO7EKZwYssLHih
U99LADHiaqAYnsLhypy1N0+k6rv1pzcBMg8wsGHzJm6M5bJXo1E44wtPRxfjF76gVr8XHK3977Li
hD4VmHnvkyHW7H8dJKvDC+kR5mZLkRXNjJVpRP1h9H+d2DO3Hw1d0mBFxhMNK5lRgwRYMRP9gvNZ
bd5JPQzfI19b0kgzEIEbjlKxWAEK9oc+kcI1L4+7SN2eD/7C+cVuapdz9Xv/9kE+LZObb0vrQZbE
EAIh2HdtCa5LJ7wnKFzU8kYHm0gARdAj6PLVzgGU+jayfEMwJbn7pEHr5HoNCF1Hf8Yr+bXhjD4N
u5oq74GRIQ3EdUFzCACwTVaz7+9gEZZp7sHQWx+XQBIjfg0G92+B8Mx3yFveGH+XNerf7SFP23nv
PvWSMaqx7qO7OTEhJrVLwFrWNmQ0D53mGCkutoSS3Pt7UPiq2j6Wv1ZxpRxIJDG8asaN7j2AvNzq
4U2jSeqFfwOFUu6wyZvmCEI07gYL9x7j0+jxPtZV0aMo8gjui4wu3sj97J7M+tflp/l0MdWgvX9Q
Pu8+CmV9dUKL7ZiGjJqBMRakIPWN3AtfmsrX1ZhDqwa5TRIusqJetYnIfjSKkxzXdgwKg23cDVDM
n9RhTlvRfCnmeo55r5ZFpfdJrw1JPvpmgzt7TbY765rswFFMfWx1mPOH/0qf5b7jze4EPsPCRZEr
kYFDPweeQ2hgoJ4m4Si/Qk3kn6L5JtkEqvGEtcHLvqHueVUNZwGMMrqeSWs6JdgtPIL5MLOcvhVQ
/+nfGurr/1WCPtFUA3702iICEDe+rIEUqWxhKm/t4y6EaqNKGGUXSrXbe6Jy7c+LGSITjWnPaThC
e6Q0/UOg8y8We+4Red2BIVZGmB3dIlIKurvMTBAzUAZ2wyyANS9PZioMcnBxKN/5lTL1RLti1Qy6
y1yVHwGYGMW/Yr3mkAw1oRQyyw8NYju1hbDltFo8ze8/zlsmppLEaXNdK3xiOvFJnzW4/14HOSBo
wfrtBzI3RLopdfgun/u2Z6UGlTX1L8kBsmTO877ct6DBVOk1daHsp6OXvPM2tKxSfAZo71Jvs+gS
9wO5hRVb1O85yFtXXH6nJAv+fFBirrxN1xyw5rQ2roHAfuTmnKGiq4qFo8B0nOUe6J1BCsSF1TOU
9v5625sJTw2p68zADBX/UPhV0IS+vbVqd67zd1shQZNEFLvSxDb22ID2GlJKnPvNCJ3d7gKq8TmR
SLYeV5G8ig2k3K53+PPNXS9nk822k/xCi4y5zTnQcHtTLIkDwGE9xbo38cX5AwKJTYK8dMiMNxtS
6ecCqD6PeeLh2SsFVX1Mayt9s+2Um8VYcQZDqTytA1qzMmbFtcrJDr0h0huiJi91Fh0GNrGq5zO/
uvZ+e5AkYiGN0cVtl2D/Q4SvegvN9R6+UVE9+UkfJObk50b2qBW84XNZmRcanLjRisFPFTXIJqL2
IaxCv9/pidDXT+UtKi2S5Wv2bNLOquL53qRs7dvSxLRLNlAuR/2qGBii2evGJ1aKVg+BZ5+TmV8Y
Iq55+cv5Gqsof/fmLBoU7ebIVhmBirT0eH2Z9sqwbELxyTD9pDNcqmpZFOvfoGFNon65L7pwOHQj
kDpQMpSHoMIxRFrWc8s1K8fyQtSKhgF92JRMl5InmhKOabGBcMuLlnl93vaqkaxx++DxuTngImAe
wCYiA9tV5l4ThsQyxzsWz5XsCGbapDnqs4yS8kp1tzjeARKaHt2I/xFnUBb53CtMzSGk4UBUlPfn
VYGU75U/F2NZA/XtfeWi+FT8ezXMgfsMfIbgCt+p1fXHQIKxGuUZWezY6Km50TBMu8ACwXJuri/n
5VTpl/Q5HC27D7LcsgpcX0jHEmG2Wu4I9cCrNOrBuDdjQ3eKwHlBMCx6v5K70BLpZZG+xFonLWQY
UtIE/3WFhoXWbVo/ofwzanWcwrEpfGoP6g1TONonVHcz8LmVbg8mGlavzhIDtJEzSl0LSaisJmQT
+JIUwWLc1Y/oPCxLqUw57pOaxyYER74w6F0xKdQN3Cvv0NQlHRUXvxagn1oVJlFba6W3yGFsw2Xb
HvlRTALBlKV+UAJkctp2KASno0Fr74HAMGurOGIEKytYPOqw1LSdzg/9r56mBOWzjl+wDBUVJ6uh
nC5BWqaeRu9mqIqtXqrGchLsBhZp3Ms8/OLpUsoD+gPy4UgmDThIudpaAQzo1yZVS5e1KfZViCwe
HLFtZNiXiho6FniLdJ8ksNiMxrRgRL60fCLswH+QWfJK4mLbOiFeTAUeR7JTF4GIbphggbei/rbq
Wt37fVwzKhFKMnwrxc3HdmXqVqHIrD8gwTe7rSJWkwNCMiRLdRVLuITOWIgZFDDDTnq52ghKLXro
8Obo5WojLBRxYxd6vz5fc4DpUOdTQlBUZ2yMC7HTAJ7S0sDdKPkMI/Cc1EqhVtobNC6Vl1TyOD3E
XOAw8KvMkVwVu7cxlnr7lHdnSjOxHfoRttiX4mzaOIhZw6P7PBMu7Qin6iH4BD5/zPN/9YUSB8Ky
knHqFCwrU300lmD9X/mVS4EOKMFMzrrZKZ+owuVB6tNBP5zgqu1dRobG8q2MlWeHMrc3QIWxohJE
O4DJQ1aMC1mwYlPGznVED+42U/g1D0OUg0udQwkFuZICPEK6JY4dT+ucaSh/aeYBdAihoCo8s+6/
0DWz+LFr0C4dAZNg76OAJgMeREv4KfFIPo073qIZNnbkf9pb13c2AydGmTAuHWEigTP3QYuKqVDa
va7GiRWMogpSYnNdjopmLrKiK+nkiFPoJiyxqKR/7XW6KkWmqQrWsz1MAcoZZC/6zx23O4RKH8zi
MyJFt7lV9ARSE7TX4s8OqQ7FejhsZaUQ2xPTeam7kftWurhrh2OSzO2XLro2nQCqi1sMiK3dTarh
RgGEB11wlnuZLqEXHJ+E5wTaA5RhLeMk5YFI45+lHLP0DB+xvR/eDuqG21nZcuS5J60uYvDhie7c
YsWkhRlBykx5FsBjZOIHhj5UoqktUTvXnF3oBDncyfvzAXfCYrAaDDQ8CvWtPTTaOiK2wHqaBM7f
AK/HRJUH4zhsWDfke1Gb6Kcqq+lFUF/PpMVUIObw6eUrgnOyl2O404mGdIFwl1QoFuwhYTYAHSAI
I2XmDFxUdMDi+qzWGoo/wM/bt1PeGSxEudxbqcq7NAoxkVngnIQnPcCpHII3LyiXR5EwdIRIwkO+
PppLH3Dpp9Ex8H3ltVBWRJJYBN3tSiknyDZNZ3eGTtebopn071RukxNXqD7eVTdmgLM1L306aYML
pUWfQjLNUlhd+rPn6xv1moTKxahdZz00v76ytbNiCPPb1N+CTaeOAnG8Ruoo8hnjKGLzr0p/IhEu
IdmsG8nQ6/zHVIF1sdtJmtF6bxaGVQbIbvLYN0GKQ76TzPCweYTN979UG9LmvKGk5VHDldlGQpeX
H0/NEY0TDaYzLindB62hkgB6g/rB1th0WjPIU6UqtQZ9kgoxSlYtmeuWq3cfuHbsJ/up5B+5Im48
bFhOaoWdDLYkJqFs/lbyu56SRcHrqOB0YF15Y0nM6q6pEzYxAU2Q+Kv9eyi3cZ7AEZHkatqdciN4
C3m2F6i3X1H9YKcoBSn9v2iw2QZnviPpz3QeXaTxzN1Y84HvHVcofwTJubJFxs7XbyR3xZ2DmQiM
Kx7uJcFSFWkorjHABhPy/eFVjmer8l3js6n5RlkV6vele/TEr5N0jM9LuR47oVX89XVyjJK8Uce3
xz59EhAx5BN4RRBVHcP0iQZAdPFgBAee53tCtZiWcExZO3ksdibkUMN4QojLXysQatKcX1dk6qN3
TN8SFKclYE4YtpVn6Fr8Okl+vfS1aMVVJP96BmpuMufAg5ZqIrCU3T98rpP2nwbyZfPYIlrKNecH
zZkQhNAQhvIJxoGY9qmPyLhW0Z8X49799ltg+9kjsFVF70Y516MG32avqVfEss22VYeOcvZ2O5DU
s/HXavppRnVDQI7JPyMYXQ6XfEnFuY1ZRzAE/o/eKNlvKRTnpKP1ggwPDjO4sjcznNnhEF8iL4z9
1FeFhEZgwMZ4VcuYtcK2i9wel/W9v0vccq8tdl/5rhTimfqPX+TwZ1SYRia2UNhBAw/sCb6ujVyx
pU1tSo5t7tBC5uwKyoOw8qpxD9a/TkYwA8mUdycVWhZi1A4E/goq3noYr9SiFa8vYBOx5MkHiAJe
vFRehkkXSU8CUzwJrq5ty6c6z3bpJnwSIb+XPP9U6WMPFmsvXc6BEMMqKF0b6gPckTSY7o7MQ3cR
BIOpKI+RLMju5xuH+UGAUn4qXJhB+Jqt6dIyZK/lnCweBFSkLRmmLMJ+SlK28mXauFRrgDSMbou+
UuOimL6y0pYuvXganIAHU7/zUU6LqQS4/WQYMfMZoruqbFUl96CeZYxo3l3m4+ZmxUPMxdobLAud
RMfxXgj76vvxk5tPnQh8jsJyubze4btdx7AEza4x+W+QjR/i5X12khF4PQ/z6780Vi4RQthXsPmc
8e6ei4GyRafwUiRCt50fbz7lMsIjc7PlAETuiKN3BeqLEQtBoX5McFLpQ8E3YdzL43wxdi9tbVJt
Di+g6N0VFN/r6ZfzuFvg6JkFgaOeFTyRfVPe2tDKS+H09ZwYWj+ZYk8M0phAQiNz2/RDOepNU9zz
euEpptjpNFQ1iq5a/HMGAyLkS3QbfJWAOrrVhExi53hkRqrX7UYgFeMbRs0fGuTHFT91cQism4uO
aoT99m1doG3877tChlTtdR2x0Es1WuAGGVeb7B5PdgiFSc2eyHK4sw20pSZJ70pRtkdS6eySeb5n
nxrP/BeYpNNgWdLFRYf/F8V3hC+5/r9sPlqnnEt8DIOZF9j88qJYABls8D+jmtfq/dvOIEHRE2xF
xTUBX7kqZ00rANFuceOTuMv3IfcBSg5TXEOUtPp09e+BqIjCN9/6Jnw61FD63MjMgzQ6moEYHEww
OwXBpuX1pRGN+CWYLBVQyGimfBXwoGNHSijiWOaKXBAe51ekRGnPIinAgIsGpeoUnC6gS1AES9OW
/DUdjMTm1AMEFUtCrt4NyzEMLFCVOL20zqiEwr7KOESdVlUz7XWl8VxLbZwob9NMrNSkOBfWAMmG
u40Hs73g9JoztR5v9NY2VDbRjBdShY6UhPj2+3Bo1zM32bvPit2ZaPkONtpo9wySH92xj8dHh5Mr
tGf4JIaJYBaTTaMFKhBOXG24w9oHMXBSn8/91+bhcqmzrYD7UuhuFYZ0UlIXjdRPBerdK2S1zyR7
tXsnkw1VMzfV1v5PyFp6CBp7gRvjiw+l2YeOlFy/qq5ojP0Gg7NUNqFVwh/oQ+RXijjROim25/UJ
N8X0EybI+ZGov7ZyZXr7ecxYbPOLwnA92th/Od5fobxqA+0X6ykoGmtFeg6kzeKs/ZE6+GRFmyFN
kyjMNhWiaC2yliBkEIRkM3hKrfxkN4Ri6QMho0b0MExqiHAbZXT5Qm6vMe7B4iInExcM4uKIOZFw
3ls2jJzQu2oBwM6jyLfFYBg2iwIOyYmybZoanL9YfR5Djz2PVN+r94yp4QtDr9hwEkX6tZd9bGy8
on2ayZJ33hddLKS8yLJq+xVZKzx/iFEfmIzba6sm821RrWT+vQ4VEKQtJ5pQKuOhLfeS39PuEIEK
6cWK6XDpW0FUqO9VbsrD9cAqZYqKBdk+kzrG1QmQZCYZr7UufcxqTP9ckasXZw76LTOHHhtXIj6q
2/nx5Cgk1uROuQWubfvKACJUmXROqcEKs5B88J6NOOyBGtsxZfWkZBezRZmwHW9EbYAlAP+nxhxQ
/ImC7pdsnAJ7+4lm+Umw77V4LUl/RLjaKxBxwMPihUvt12b5X3ddGto3/yQWbsOU9407XN0X7Vv1
tY1w6otVJUW8k6SdSp1f8TnHp2Fq9LBYgJ8bwxcTIvkkX/8Q6+faA491NSUCDTPl2gokKcc6Ei8J
oPRuQ8k4+qHCo1x5NkrekgdBbUugLCc0oPM173rXD43HyMmrC6B4DX/qz94ll7J7MGAANUMLe67t
ZyuWRJBpRpZ0iMHBMxqA3EQzJJRpkcFbEUXmgCJjqtGMJ/UdzflV/WPRPIYZGfvdf/S6YWPapcs2
exmPvpOmFVOLrQJ6jrY1ykgHhOQJDu8+kSzhEgTz3ETxbpQzAwJe00DpqK1wA5UOxRLc4RTdp3tm
hsd7EQWGIM3rPJ7zMgOU/iEjIJcU1k4+dI4M3RHDip6xTaNJW0Rb4pf2U7xa4mtxjcEUfWWoFtPC
4OepssEGD8sldjfnyt8DlrLjc9kQ/VcI7L5LZI+AS1x+Z5ENLtqcaWz9rVENsj+iYZHLjotAmquW
is10O237Hcnd4ThPQA840uVlubalqCuAHeGhuJWKm4Db0WoO/25X9XeBmtdpa6kSfYv45pUq8Zdz
bttg9pIXFkCJlmFrdQi7BmHN4cDMYTQ85rgcXUyeYheCbQkxXcGszcQqdCOYlr10oJbqT5XuuzjN
Z1AqDSj8f8ZnelT3s/QVuFynZXE1ZXxQ5SXZVXmLMNSx8DDacNTmovFcgdahx1VxYO95A6Z2oppt
WDTjDZDGcmDCB4XfP5D5MYXmmjsTf/LbnwdPoyONaRY8mMxR6T5TAa57jJm8EMhu7Xv/eE4cD7Q1
V6qW2vzCFTrIp+8Vvz05jkJtXEyBhohK5tI9b1Hja1uzvcsjvsdNgC2K6h0nb6QR/VxBvDRAHH9/
ZkKIgXgAKFuIL486ktXIoVl5BF8am/U8SGKDy3dP2F5mUioBF28Ytsjf8AQhDBsBrJh93FhtnLTd
KwxmX0PJk70h0FvwhzmThnANj0PVT0wDkOrK7ClKyfdEKfwVBKn5iW1FWo/M9ec5Zkbs78N9vPEN
xqkcOPUdakqjwjjz3bXkoi67v4zqW3GXBAp6Z4pz08LqR9dFFzpZjleXXXYCV2qOXDecpNYXixwf
IWmFSstTIDy0pJy3qt/mY7Yt/jSfA9VbY058L1ZyRT+uPjuuUZtsvfiOCcAas1rV2JnNp0wPXMqz
QmiDbG1LzKrrWnJjycBbvjnt083l1QW6dv9iZDM2fHqN6rZIWQM+mStnsVyKdRdZKnGf7CY15aYr
yK2K7rkyA/u1jkJnTDuLFU6djsL0WJ98FLBIwqBka1MwkCYYKOvfCWXwzHmMGe55+UXZwbf4uyGt
0QTBS4dKDGkISNMgvXD5Oj5AfADyEhJv73Owhl2ZU+Y/g+5YGzSvbwqr8NqDOEdEwwtMOuUvtgdR
imYy/eLoUsGbVK+gX6d354iVi0WGHbWLVmnMTnL4LU0iOJWaOCYE3nReYzYRV5jtBKXFAYp/HlRk
mqhXNWCedRZJgiErJWHQG/WPCmfuf8gLE905tOqXrIzGGKaSXMExEk8UwbQVPBMMqTwG8CV8b9yX
JK97JTe+b9yevLrBD2a4MQY6fS2F4ioeadtPPT2PUmlNpCdrsP1Mhq83Y+YI+8qXqVAOFBP/bWFt
0hCStlgJC9JUwQIlnYxYIaI1rbK4kDAYlOPMSW1BcxetBR5bd9Pil0VeK28ViR870J/IiBGn9oPO
AFXNObI7lvWTiOVW6jnNTbiI8Gie0AsujWq2ZC23IIU84Q21eTVhm7QveYLsoa9qglqUvEocZN3/
LVYd7G4AfJ2+j3pZsjrFwNaI7VpnMRwqGz4RTS+1QPJmZk4rTDIefMl0e0v93Rbn5Ii67xbpmEA5
DNS4XGVKtalr7CTr6yQGNuzS+w5UUiXB4cZcjIFR40IH7d0z03XyCUhHrarSjjM5+oeGew9hQEWR
pMMvIM1nuNuP9sx3N6qg9TEBK/vi7Kgj1KTtST++AvKhTm4yuYcIpGETZkPv9rR0TUjUvLip5jDt
rMwG4003xYjUChXHY3NPo2AUAhQlz5CouIIk20GI9SIsGueoY0ywgE4CDHBKu1pWBIFPbdNO78aX
Ts7ZRfuYxtA9uxMUYFEXLYd6EVEzE9Oz3YT1wLjW1gqxrDMB7qUy3WSbpbshUaKRY7YBaEeSO5By
wScnZ5Nc0/dK8iuE9L/9grvM/642ru0oYqTJOnLy4dSn4DFZJRSwN5osaCoVTiZpz905/DHdzuK9
8ISyjwUbCfUpMpfHIk2HoLR/Szf0ygy7Aw1P+2MlVjUFCfdx1nsknay5P9tUfF3QAfG7S45UnzEZ
GBv3f+EXZ5P5tenBoQQCGl5lchmwRmZk2V1ZkYLlzvVvtk9C1ySRgAM3I4/oDkIB2cdmWbuQvf6A
urb8LCosGo2aDiMo6flY1q4y75F0Cu++EAci5Ec4DveD+gdYfnGLFxuCpT4xmM/j+qB1/t1tPJGW
R57TH/hIznlHrUtj2DId7VXN51D/YLgbzgn8nSHJOM376zoVFEynJOhdmu0VBYcsAu/xnc/i0YvU
rv2ygaagmRPw6bZ10C1uBY6gVOi7uSKpCA3i/uTMc3v88uty3R67OppHXr3dVFsTZ8YhRGFC5wXq
NrteeGG64BNJ5nhrD/xsGYQsn++2GkXFb8CmmdKzu5eTjIEQmv4HFDflnnIyp/0cJfhfAXMMnQFY
KEfaGD5rD03fie99vIlxMPXG7NjVqMcRDe6jXGv6iOcg6X3JxqkxNv0tHu0V4/fIh2F8gDRZT+Qx
vFysqKRQUxb9skioLwz6zDtt5Ir5Tvd9nGSUMyJ8Ooc7KVJbxrOWYz0xqP4Nnm8aZOq9ZgFCESn9
YzTUuWjcTxUz9T/J7cG2yhgPKfbp8voZtwmR6EfWMkhFO3/zMZjVYFtghj2bWPr8tMmerY0EaYVY
gOJDOvSktoeuH5srnia0cIN+tOze9T03Z8tahXL7Oy/d9dkc3vASDBZ0GG4uuYAG+NHzQQz/8auT
zXETMBvbCTAhu02uUxvrwZdfGGV1YBD8iSpJ11yLTfiXNns8ivzDyjeV6EK5Nka5xOGijkXmpOoS
Q3tKyBexXD6H7g8K4mZ4k3TXKcUu+H+ZhLsG+0nbvw4FDJnORdcsy/x9ZMA5Y7cmBKeBPzJchbmF
tb/XVIyQtKcEGbUMPB0Q8w4SXUvwl7cSIjfjCPIujI3410nnr57sHNA6nJqtfOLMRlDKgifwpm93
Zwraa/JpUf/+gTnNRGJgc6ih+Kk+g92xXuw3bG+XXGLMoSLcMWK8eXDiQCzAEuJwKhH0PNcWTJR6
PruNPqNNfKNJLthBQOWdzlPEpDoag8/lu6uNr9Ws3u4qMkfiahh/N+FpYPEY8mA2L0vEitEcSiLz
3ISNLM4bQhxmNPxkRfY5tSsAJeNCVf065KoNtc3kCchjn02bCjOOxIE7e0GnG5ZMZuVbityx+hgD
vk7LnrUTf9LawCvU2I6ufnuU76TUv0ngkOwRvSa27uhsW09F0O8yrwHAUvl13OV0C5LEtFZ+cX9O
m1ZwXdBR8ihllfxroLsrIFqG7baiNcz1KRvKL1C92xVQcV0qz9t5OkNB15yrDJpRYvWmnGRGakUw
hzGEGJ1n3KBp71r8wLpnPVyxb1ZeBLdvPLtwPEh1yNiUFB6WsjpQSslMD0zuN6U/64oIMHwbaLj0
xGTq/dcy8K1/GzBSrhXZu8YfSgWsaL2MKbEeXFEd5WxTF1SfoHe+Pf16LHaF+OoOqd9y6jkPRY3j
CZDWsrDeTpcGqG1jJcXGQG1kJc7vpsqyYJunNEWbzGxCxyd1k1bOnUGwwo7hKD6Rc96uGotV31Lb
MxrpD6uHPl3O9Fqz1Xz8m/8IYCkWLE4ElWldIEQ04Erl47ibV3BJ8H22SOu4r7NKfj7/ijirY9iL
aJWfnSdrGOcsDIoQbBjORYPPChGLu0vRXKt6UIF8v/IXPBst+c0mIbIh/DDUh1qsOJrksc7Sx1SR
PkZgoOYwK59G+PemHOfd/yFLnpwoLsUx5B8eWM2rQYDvMYz+m4XCux6OPRyomRKwaQgIA8W6lmz0
Wd2wpG4WY6SV5lMkrGBg7zWvGH7dX4lN19CF1puJ6Faw90IJptAVuTMhPUyTt4RL8tm/8cFuJXk7
tSetklm8G+787se9NmLGRTGCMI6ttgoCCk0RXK9/5PFFI6FSxzr+VIBV7xSNeymqVDm2Zin/3WPc
NHyA2FJn+MI3g8ZnETKVqISo+iYqSC/PxW1RHAQRbkxdP1vsDXBqa4COHXt8o04yLeJdtB3DhQiZ
1J1wiD8prNH680QyQgcJ74BHo3JllGQGgpVkV2C9yNbpueg7SG6mWsIWy/Rfva5zWSUFLdpHmrXc
d+SU4mwByL87NEDEgmveflhllLJo5sN3mcQlgxrIot3EyW6WNKUtgNpovQMmWNZigxtPbT8Kl6DO
jWAw1B8jSQxWu59mCOXeHAjS6FAma7w8p6gAbPgALor3JJGW3grYgdfNjFKOid2k6+Yl87AlOC9u
RN3KeR5dqCyUM10temdy3czLxKtSzykGsc9/PMc3glwPvg69AXmx72w/43LQC5zUkvqqjj3ONmog
evbSF2IC+tUczzW0XouVy48D72seoD/+Gfyj03nzu/3SzsFv/To+zt2yQ4KCkumbsUVP3paClhWp
9yv/V8I6YaUqvLxjQTm1Sv+Je4jaaxMx6xR9+OaF94GVNNJEEM5anqsx9COHPe0e50Z2DFE+kdwK
j/cw1O1gp7P97RY81+3PLcHhRHAU4jbcMgd69YctUes569QVkvdk5gTtNLd4mkWQPoIWXlRgX7r0
PpU81WwLGRPlV3YWxlhJ2V9gjd7SGn05PWgBMOHrzl1rDfHiqumt46kGh4sgrezg7EDjZcPVR+FR
3rdYDR9KvUDcD8RExpLxXJyvuAmjmgGfv4moM1o/ccwDIcp7EJUbZDMl1z55fXbihjOLCyb3HcIs
Pg9zPugff84AWbvC1jsJiDPE+pZ239Ngwxw+zlmhQPNj8Sqblzsf/0qm6vdzEPkrzb0NT/s71Lxp
BQupvurHva1K7jeU0UoKvkhMhdVOU4cf9UosK0S55QFg6rAONeK5UAQAGrUu6pwyppgsOwD1xxY+
VlhIyLgFbKIfSkx9ih5/FyzybaBD7v34Yso5Nk2ivosV1efupt/FBbysYeGnOPzk7xr0TaOSCXv2
9tQJd90a3sai6tyRyX186nc7bKReYUAF88geysOwYCeWY8pLbumF3qu2Gatg3m6QKNlQRlBn9pJr
y2+xKCDFANcaE+HS9uwGJAmdy1KYopFJ3/v4SLZkClqFkH40yLGBiCXCcWOFAJRTjqJzoyfuFgD4
ghY/xzpy2xbLxapJjAVJJCeTJQOGEbel0ThPf7dDuRoHRKKZfNU2G+vTLb74iych5Aha6OJZECqH
7YkD4I8zITPNCxYKeig7gBlr06rmwbf3xNJdiBHO/+y9zGRJqpDZ0WPR/86p+mRjhwLQASpRww1L
RiXdWmw0+b96m8yXTG5oSwzUqsCJt9VuVgSaXWxwQJl+d4yoyiF+7qlGpBriQdmXBiTd9P1KbqGK
9CsWgGYMg8oXpy7nqE9jHxTp9jadmqIvBCueSl0Nub9LRY+aafUzgoAiMgHqn8UqcoSt+mU65AjP
UloIxPGsXGw3yYZf/PMbFQrrMg7HDdK6U0aRcDMQvJ9x7FMRrba1jYMELTlRnDncygZxalPCFfto
nFkus6h4UULBpi9y8BwxB5Y61N9bNab1/dhXkmEleMt4qyZprCicCxNAB/9EHvvGwYNHO/bLZg53
OvsE2oGn82msJniGEz1JFIyY6Te8r+ok/WrQDteHzIHhHUrhbrYjsxHufUlroO9q1sqmL9o+IWdU
YTCLSZ3uFIYMn7jmuaNpGYcyNx8hmAbYClUUVitphbhMhMIWAv8gs2QhLYIO6MI+Ud5g8Wm/4PON
veDPlSVNg/CtQ5Lnh7601vcHzsJvApO/12E0ofg7eH5iWz1B9GZF/+d6ysyi0gkJxfzEf+ApE2p/
anN3VeKI5deTBq/jhPtPkKbdd3B6YezzwYtTdGyey1UnC7Bu6StDDUJew6wAdDpFOgLtra5vUlkg
yKPWlc/a8TiRwTfE7po3dzisInaVYUoQGLch+PYcdn6HsicOsyBsT8sBPp+bW2CU7WknmSBn/nGn
U2C4W2I2gl+JgljLw7XM25Lx00LQRnRBD0MoTY2pMU8+qk2XDIiYleta0rKkjiVHZmi1EJ3wZiSS
FYT3Hm0PNwKCc8yhnPzbwRuqXcyGkziqqukP8mIgdIIJNQnwOCFcj6opZOJagNplObq7/kkrXPJ2
eKSCb9Op01N3y52za84KLWPq5jh2T2gUD53pDclEXqVLmyURTMhcUFn7vRyBgxbb/NxUDifjIFJj
fGNZ9DNugWNLH8tyJRL0I2ncZxmdZHG0+a9YUUUhibqr3LVTXRsoRzexo2trW7dV9i/8Qhd0j6H0
VVotmTl3ohg+M+UFViNCBhePid9tKMkh4fakLCr7PIeuN6wYLV4FTxY6wYKfKC9xgsFNDN8T7w6Z
1EIo1IJRk5iWmVKc8lPbrZr3Dcbqssdp1VV19MZ3C3PYojFCV/4r6ZHMGdFCtZS+5FVYjAlo3NI2
j4eXR9G54LogI/8VUExzYNSBWWmEVX5K3XQMCbeE2eXP56MzP9ENkfcYgbn78BHHZUOJS7lMCGUC
TBKlElgDzDcZNMf7lX4TD0XYclsBXfGDYCKyeCJckuZpLRHvtRVVSAYFSkSOxtF/XijLMkrwmfWc
LSzgaYnMtYfjQnPBViIpfjoswKPKsVENCsooNyD91iwwnMvFB1MdRKkOtR24SEnTJSQOltruY/MO
TiW2JG7igYzRGnvZlGdlwB0f8dFQ349q6x7oxQYVD46taX9V29lH/txHR/aLEngROnXblthfPvq9
+utLCgLkiVKoBlGDHvac11jRQ73QFjcJ739k1udUp5QKWxRpb5wICkn/P1Vw2Ueq9Wajyptf5tZ0
XRGdP4XllAT33ER5jycRKV8DLqIrGWlklwI0tsbv9Wx4XkAwn0R+hFnvt5joCPpeMwlNahFJkSY8
S7795LEU+JY+3g+i8Cz6ZHaks8w+CueIZUDV+EydJgDuFWuoIsWApkCpfCnM/38bcxFfiFeIfLBh
3a8PlC28GGCFA+sXykeF4xF3dTaGwmE1GHD0I1KtljPCwreSHfISmrnnDM8gR1P+xVY0EL++oQA2
Iprptlr+1lVgr6F6h8oG/V8Kto8Ozgl6kew2XZA5LlUYHPvW0LTTWA+U+wAI7on8KJCzuomXz/Y6
4z34rGeO/VgWi63gncGWDvNA2rbqU8dx0+jYGPfbh1wvQScIDzLEMaDAyCpJ0PEr/i9E6MD2A+M6
KcWoyKOZEeoQNAqcShCZLuOvv+cm+6qrbicq6Qr5XPBk55CgGgMpXOkIO1UslevGL/go3CoHCC8L
nIVEaBUucRBKeyLoiMJL63G3t4B5mQkFRiesl03d+rDU6nPMbKYW+pP6oZ2dJMFVq0dS8a8QOF/d
gkxokOT7lRLKd37+qeR7nDqWNs22ITIQA3zi3YnTG+GwKK+w5Y/sa2T8mLcBgrFIUxjDvW3frokA
wp67Fu27hA6hojD+CnzBVrH3SNPpwFkYcSvwai+ZvqM6PTC8DqUZrvsuk6y6Duul0dkluCa0MH3f
FNmy3tzbWAaVbRuFmGGV2RWzU2GJXpI8aYhgNtiEfS0R9+g1qbiAr4Y1BUbM19JECT4CVXUCz1UH
QSAzdJv9JZ9TaCHjAO5/yDq93FFU2e56cHJ3KjACimzHap/2FelUvtaHQGHxtblmlN8BWSxm7IFK
1sy1viuaFEZjQ3QbPHMYRp+9UGRrKs38K0/C1P7T9rWFz5c5ZBZXoNLzvKScTgIoxhs9BYM4TzQ4
0DSNTjbjHwGTQZDSAPXqu8/7Tzr1deOeTMriRYgJFoOpHLapoi+f4A+m+VnT/jIBuwSSqiPG5dc6
JCEkhhHPb3sY2OiEXYIaHBJ9ofuLk8QJfGYk1fbMaQMMy0dAtarmWC2EoJiqOqL49B5zhuOvUwxt
2nrK4gEbTKQYGsFfjc6x1R1s9GcxZFxLqvtq6ALUMvggkbgY1euFquyjEWCByVQNbO9rcv6vFdaM
pY8/vbQL1x9JNN1melpWmjEOQIJ8fA31NiKIeLOVfXLIHwEjnRwlzillSrPxc8xtR3/XtIWCsFFy
KI3RbJt8J1IoUNZvYkrtNS9XJlw7kDGlZ1cA3frgWaLGM41kh7n7LP3PsjPX4VDhukqPvsUHxrlp
5dR8C8oAS/5WBSKUGNCPVK8luqkKiu1AXYOlZN7VYAxMUTd3CZPsmkQCvhFVff29lZosfLUrqsq6
gdgLoUQ8y9lP2GG4rsXuL5xvdiTY51MwbCa+Ep7x+HIjJQpIz+oCK1Z83uD139HbbprNtr/M0iCu
GpgqPUcc4VtzlH/0g5w0Uvot50YjQnuHfaZhtQepbFu83Az6OuQM+584uuioBm4Iiqhg81a0PllK
vCFpbPp0+uBBbLjCCe6UEo3IZns3Oe2N/pFBg45ub576o5jn3nOfm50x7DCzgRVqCY7NdacYrsgl
QclQ/hjGMXlwY5UkIO6gsNo29yEE7PjuUebuxmhnIlvAJcL2u+wHHrBqIEmMIm115lrFdvQV4HeM
eKHeFPP3yH/9qv00lQSJw/zEkL/2xmGw9t6G4UJBwu6344BVAMmKBZYaH7niAska7MX7AnXYpt2j
COjzlicc1zLuCRXfQuGd2PS3TffIj+ODEJYZkxQTSo/DwK9t6mBI7J71IkClh3XTVQ8fzmsmHCQq
z74u4l6IvSt5Cq3ySh3nEUH0aqA+pVzbf90DmkAV4j1flh/aZanONB8+7wyqyJ+8xizmSvOXULyl
30OmQHY+W5DskFWi2VA/boEqv48zGpbdeUl0VvIK1iwplBjV5HZ2d7uMagqbQUdDV/0mLy4zerHa
ZOHmzPzdxc+UypCr8wdFjH5Enc5i3AGgsIDS62xyzzBFIMrVO3IdpXM3V6X8zF70gSsiUJCV+qnM
MaixBBtm22C59ib+Wv34JxWWqcaCcV/rOF+ABXH2MmEVpkXjszxRsOaShOb53zj/yfyHtT1ZPg+F
NEu0aYVA3cvHqITVT2+7BqdSwGh5LlohdobJH9yGwYROXTEA5Ua/FeWTK4pOosKJE0CVQhZVJAYF
YA3ZbSU3hfXwZkZpWDjCR1uewAd7IQtpu3KkNN4JcaQGA5UOODYja+WjGACyfDuQ83o18AG46+TR
u/JKIUJtjKBCGtUVHc55J6a2GmRqBwZfnFSrXb8CCdB2wDrF8ZxHoUNMEkMXqFMN7exTuHXzAbGg
QIXpjVLrvlhMDk47EetA7qk4C7PG0wObasznzTlALiGEaKhZGt6S/O3S1VyA71o1VIM3ggGWoSxp
whB+oDxuzi7PjGC4K+MkRs6xI/WCPzN3ZzLn9lkOYqI4u80OAsgnRGXpp+fTFxM0j2AZ4L8iTsaq
hRbzh1jPjF3QUNbULF95UKHTOskpVo47SgKifKvSekRWjSIR2c7vgqaoFs+ICslfM8BNp8d8JndA
JrBrr4yNQtDDTO2uD8LcEFUp6Tcm2QuQMjdtFZfO9O0kvdUw+8SnJOSCkhzsKFa0NhcdSgFPVZ2/
NgldszfO3rkEGH614z1dIR0ExALY2x8xQcESjBjZrJZfAOwPipxAsqjD5+iQcsEI1VbAUhYZm3z+
8fUlB0Fk7t5DBY7Tj8gJumIq5/jBVwKPz18Pbar4XzZJdOjDo74fsvzQy3ki2mX7JOtREZGc9uJM
wMCFcwHDYjZzppv1S/u+cMLuhe7nzxNvG8gBWmJZ/RzrzD5u545YvA6vXUPxGM46PIShwO6VljAy
vKZC8Kkd3t+kgmjuCl7vjqI4MEL3YiF+K80yxvvKJLxvkfz4gK+NCUc6x6SVl9qsDPVoaJiHgM/H
WbfmRntkJ/R7mqrIBpXKbVK8g6P2M39F3HoWY38sVx9IzV8kXKW/qBREMVFpuktFNKrzpN9gbtCl
X0dYueKCVajcTYT2lGME1AL3y+Uwf3Dg7b3PXASl91Mc+Uq8S0GmHkU79GsHz91Ci7clAVoopnGw
TgijAjnpsR3yett/hifJHpGD/RiGDgzZlwpwfrYC6UWBQPRjcNz/wYEvWknClBPjkHsvslXoSvd9
ZZXns+GHjYwl4dHXBwWoq9hCjjYw52MEYlYUUNakyCgjnebLrpv+gJkF2s2F7lsrG0c6jtmytpyj
T8tlxDBU9UwAYfMue6UhYJmjB4rRe9BTRpHCqeX/+tXx1uyJw0oDPeYIQn3hOc21v84ZaDaCjfmN
vLxvGMjJSFp86DbJmHn0FIPdVE9cOFwgMn6c6K4Ryd8jCzQIMPqqRCKZ4DtuUxI/9T9oo4jO1YRX
j22O9DE3ff2xWnP1Qkl/iJH8MKK9rG/3TLXuHM4RvPtRPPKDKpMatUfnGoJ12lXdQm4N2eoCTmMa
PYRiOlVwdAxMrSELtbZhk5TacIvUojjXWwy0lZuFJX/pkOMQhQ4NdTYzwzw5QyKDupGood+H16zD
u3RCWePs7U0ho2kJOW0rS4zzhX18u8H1RfXR4llLGxsu2SnaMmziqtGDL5FBpSPPeHWk+3DESI3I
faXBm/BykLimkqLTFHuwLlsrzOtyetgw6AtQAt75VjamoT9o1NINDHNgUtBx21THWVRyZsxJj5iK
F7T28qG1OiewvFr14ZRoiFDH56oEZ8qNPjf2c9o44k598L1B1Z8+LN6UjGrzV/5KQpof5aV3TIoT
fMLjdaq+1EGteZR9sdj/kCiBvFwrym99f90bzR6SiLuBpL0wsOE9Pw2N8UECHpyEVUtfP/brALb6
+SXtNhzJ0rER4Kx7AvKVqGOsWSGAOezcXSOyzMgFK2xM9m/3mYjTEeenRbahz/081UEAmv6vXPI3
6hgu4tW0uvm0bLKqurqF778Vy02wAHFbN2LpT0MDDPkLb1oXRC4DlJPoc0US6yc1clQPAXoN2ZUI
pB0BOZJ192zR7zi8Geo0K54LQhCircg0mi0mBlItHfTgBF4XieBwpElS58SIENb6RYjK2nA7OHUo
aXmBfFygD+IcT/qSBEa2dmSVpiWIi51Zsm09ftXe7h8EUpyRdSyfnUXz+CjJeeThgLFQa2KluYpy
VdPFQFFy0HtKBlytUrcjGYSCwXTEkKxb7ZlBYNwcq6FdhW4k37fOuvsDUd/Brs7GafXXl/GlHDFF
3vXIrNcpnPPwSji1JtAzTiiWI4CpndDDjvVPf+bEjG5r1Ln3DegFqjEYbTtKubn2HJSAHOT5B7nX
IpyUUxBmFu5LRVsYWominzXNXA8piIBiA6QffPbvlMxV47AdKLome1bIA3j8C7c/izqayfLYOk2j
VaeGgDcvY/Lc+B6586wn8r09051RROFi19rTvub81iRE+76uiMxYR5r1LxdlpEbMgnvz8x8wNTaW
7XOgJfvJvOagQCTqeBY1XO2LUR2vfpwmWVD4eLesyr+GOnz/hq95sYNNDEDXBtGK7ShcwoyOjibN
yxfCwbQ59PSRaQEnagH9pOTfXVJOUR1dUeuCwVTKAU7G69swAwF/tC2rlfwu4IFWVVAt2uucNS4c
maNqbkz9vE2f3oIDQeDud6PW1fsDqtfm/hL+mwHeMoXJE9VqAE96KcwMpIP2b9Q+Og6G/tXKB98z
ZIDVKN83+HOP1/BtD7zQUZe0fy7I3l6I95rY8QFboQ+Lpc14McB7BGquPSz41+OwGuwegpD9WkIo
OTPFL1POM4bkR+t7kWS7FLhGqHrxXOEeDViBMy2m17WN152dnZwShRJUKJyNlBAZZEXJFd0e8xL6
FtXmiApoo4eaOw8dL58wP+8vk8+KIzrGfzr+m/N+nffGRUQV92/iN6W0inf23+IHgZlTWIDznNIC
BMrwdMSEUyimHvw0pJiAzP5AWbQUuS5cgPcjcy+I+dLlfzweAC5xKnThasBoWqbwm9HjOpcdqM8A
DHXVwwlCLX/j5C17UneKvhdlQiWBK7W9ftHYJsva7o8YigfdguFeQ5lZIJWdS0l/OyRK8g9UC6Yr
Oe/6H5kP37g2Q0WqgSaLd/w27Y4C2hEyLntArOU6gzIaZt1C3K2lD5JwVveFlHeYWqEmJpm5Dkso
0Xn7bpRtT9Y7pdw/q0SHxazOS506anVM1S0GbZrmbYvVL220o7V05K0+4ijwB7NCYN2AaKpwiMFp
3iKWA0pcbENZ1siEHJr3VPLvhd2H7AaH8L7g2Ztb6waU3zELi4mIm6AV4z1B2jgtP4vx/rmP7V5i
WmNCHLlbKZRAHIq9zxpiq5V+rq5bgl4336tUTmgCvfw4ocDnMZCsEP4Mb9pxo2q5LtEIuihvcfPG
vZxSJfLEy2A0CTCPhe+2Mb0cStYqNrAnCmUdqAYRHyqX0mFT1qd1oZfTWHYiteXpv6VGU+cVl8yp
G0GCHJ8Cbw1XhrP/vFiejwhbSyzOSvmE1XuOWtChjjAZvZm1PDneNCMhNWGP5pvv1WZlJ0vM38yP
nxMWOBffDIYwGj/tJhY9TZ+KmQvsmxUaHuYL+WV88uimm3617q7NMq2aqFaR4Kc7gugARZtA11md
IxsGbYpBdUOw/w07+LjeF6aMTWHy/WjVmXD9nelNqGXSX3IrHz47W2tmHIIQRlIGqEWQVs/LaQs2
mAZs2/5+qbs57z/y+IrWpnjFUK+H2zkAaXo444NkENWiYwxUqs0lAJea70iIhAcAaaU7VDpM98do
ZtxRoxmt79PcrvM1Xk03npMvS0gKKfsZHzJdQ3/C6l+8ldMTEfN/6DDUVAVgOhxXd8/lCaJMj5AD
RnNePy3M38LNHnP2lV9OGK3EJB1ZU3qozmYJDbtq1WrhEBFybKOh3J9tw4o2arjdjux2oZ23Ek2x
TwKu9rq40KiaItshE9xK7BAnMwDvS4bCaAXeZQG1uhY7lU9wlAhzLJjkTEhy1C9HVpIxJgexQ3i2
vTKxs25GYyC3Z/sp8X6sDyyMOI3x0JaosiyyX+kGsCnMP1K0PzWOS/sePxO4eM2jQSRDB76r69hX
5gPS4fxFrj1AJCoKaQGm1/P0jwv/S7z3Nzm3FaEXI7A4H+L4Zu+LveZmUx2CFybZZHIZEBuP3OBI
iuguFNASYbRUm+rR75TYpPf/rM3YMeSe7JCU+kReQ67GNNJJHMnZD3wbD30Xs0lvP1ErOz6Kl2iu
jkJ2b21ScUfDmTWJ6da4vS0v6Doxf+5n8JlLg+EQhlrQZuedVrai6cRhBRUfWMX13LZ7/NPPTNRL
0q3O8d3jZDAJwWiLn2k5/nB2QNgk3ADVf7psv8FYRqOx2w0EY1Sd4KTenIQaYe3lkeQZjMT4SaMy
QltgLfz0k3lz+FanBg5qn5LEu/eLgQA8+AH8NrAeSls5aiJQDK+gFVYFpcbBzxbLcWhhtSbQ7I0H
Cbwpz1LmUOAbLLygf2D8GiwEYdbV1mg3SBIwokO88UA6FPPOxH1rUzUbWhVOUd6prjcjVur4zE0h
XkT06IdanPVuppX8mntzBbtkVMXS3oPEFub417pEdeHTFJS8idyEW/i0iqfCnIOae1PgsvbczCsz
8u0KPTar1MYHJ7XYbYCeIKP2ADsnLLa+LxlQVa6zDqX4CX6Elp9huoWbI/r5Chf0/+pXxxiY7dv1
6PhMk5b4Yj+VSjJBYufmyYdPSYMg9jXWXrIYTv73gUrrOVk+t9a1nX85/RBWrQtGu4yYkTtW6RHS
YcPlbfKxqY3dCG8nwe7S+DTU2yXkBBHw+/wnb7f3jgGmlr5uoC8MxjZ8MSnyFjgEU+RGbG+vtnEG
OxaSMk+99izzhKRF4iSNRn7c5j/oUz/hZLUmrSJaCUVU+fnBN98lYEwD5j7JHU1RyWwPngKEjmZl
bvfVGs7u2oqudVnQpFLVAOJag2NWHaX9uaCfOrr6YcYSTXyZCahg/YO7O5+cbVEENbXHs2x5gige
8Kg/PaSjsGExdo7zZs+spsnAluu1tbcoENsSdjhiSBfC3eCXO8TL5ztE20VaoeBd75Jgg0G1XJEi
TTJQ9GihJm2cBQu/kCmcAjr9sPWhM9DWq1W6/hYfcUqOVDoKsHMJD7O22Ay2CabEgEdFKQR4xBd1
rFWvOtdlgvioQZy7Fe7hSzI5fDgyJ5xd3ePpob0hXIleGQO9o+AjBelKZCJUHhMb5heHXSalNr1D
hCMQVgR5vAAtfRN/lLoInY3veAkqTgoAcuVAu1s9pc3+NLK98Jo904o0v+YlLHQZ5LA0otO/zrkV
1S0JFPAXGdjQlxmC9XlDJpNCry6P5ExL98aOinzEA8L2MEbcnsD+2DKS3HXC2kmuxbtniPKp/ZUq
bQB2/FOlzCFtYZm2xwDgezzqqHZdtx+jCi8pbNHe8IuPPJS/PfiZ2MkCvVxzKmExhDokEYyZ2t48
zZKeeymbT4hRV5lnivdjZOSlChCRWpWkueFwXGSLM9sjFwgUaN5YpDaIvbVSC4M+EulB7Tq2Kh6q
QizDu3j4kjmM9S+fLVZ3oDsqKqLmmd+EacSlS3b59XvzDYBdAlNbTMXB32onh5VFx84WcIllVlpB
5Y0plHEjOaEvitytCiKAxj9sNQTVjIP+5EI6cRaltyGaRBq+ctcgW0lqSJUKT+NdoE6h1g5MbRZ+
Ef3wAWs1aZTkebCkDpnpP36iqQdKnKyRu1RB4MfTLokV5Sy5UzUvncDujAn9GS3A2CWxc5hxwRCw
tp7yh6/zR4VqusQWDqS8OIGA0aYX+GVDNv5Y8NQJjc6Z7qPmdvw2vb7jFqD2xb5qv+P9kjJRve/w
y3pRPa4Zmfpcf3F1CLqwTpPH5gb13W/fA4RqHjYkFtJgWO3EfHg4hS8E/q28xx+UpvuRC3cLxKCv
z9vkYXTBZpY7ftIeSSDOofiWxdJgtzvRLmNo6SHsuZHppvZpZPObclh+gWhBxPAXRnB+knOGARsl
iUt6su7fhV+zyvKuZY49TZN6wYeeHx1VSCkknrxXdyOzcjqw1HfzFLYUWtFYBualJdeQZKIiLEYo
HZKLGIdhfYD6o0C53x0Pq/fAoiMukXuI4u+GwU+e3MVyK/Z2b6idZg420cOi4oATv+W31e1KAAm+
GFTO9rHG7N1IypP5LXGbi/7eKgC7g6arM49Hdhb8YqTktK6K7NdXujqa5fismvZ0waemCntWtbyV
yaamMliSFWD2UBUb8wXvBN1FGaEIIwoz/6DTC7ZK1aqiSruRoZ+kxJfkMvl8SWdt5JkOLut9ne9h
1rSQrqK6VgO8p0mnitSunGt4K8iViHr4+I7T3KzStaUqo72x4n3ByPk1IiPQw/1gc9yqDiCH0Sgo
ACQE1CwqKaNFtmq6lUeYWbpucpFgTmgayl0XqOXd3nIe2amv6rhpapnJ9Lpp/8UcqXGj/I0+hOqQ
A1bA8HNEzbgpdHvQuRqBxqkOXZwUfVa/8aQ3fcFcm5WrYilMYGvHJRIpo+E0S5TU+Rr4w9Pc/rci
aOkcFk2X7RqvyWvONamE6L0HLZ7dYbdRQABeAYUzHCsHgBjnzpFf5Sb2IRr7qZD00ZAcf4zBFpvY
h8TjNxh0PjhC2Kxs1FqmAC//AEx1RlQkQBYEk6b9viKt5AQc78NGt4y1d/L7G5jqOFVLa+Z0B78r
tFyvRlZEIYQlcSs5j22wLxQdAaeRxFqP0onO+U/7nDiMPOi7FGD5FOPVltPd/XhkboBVc4fg/fWY
5YVH2FWHW8HlDN944gxbkQ1Qny5PWt7+95LXEcLcRpPMxX67w+Ni6Qvlg+o/vGcd0dEl0EB0FkO/
MBRBcT7VrHDsGqiLwlvKpO0Acnzmt8svVtRMdE3nxiscWd/GNqyh7PHq9nq0jXy2Wo/O33Akf4IS
NfCSpxec/McRKEINbGlZdBHM2J+CSaca/G/4vKrUDZe9o+zCdrm/31IYtJki+r+eY8KvrOzedcdm
FktPIt/D6HujcL9WwaTIvrFsRQ5PgooGJ2/oRtVl2d/YyQR+IYWQ0mSSOitftJkuKpaYX3hz6Ds7
IAXeFJnRKLKf3zZrITyWlvoNRQ8cZc7wD6KG7m0nSl5bAaBdRixC0D5STAuPKevK+vnKqLLGBOH9
8nSTyJttYO8VmDY/x/oeHp84Kv5xB/VB7t+k2WxxnhHcwT+15GxzZ8/D45xbj61afPpRNyL1EZG/
ywmPoGd+mW+JJ4xnlLfd2uzFy5WSgOf2wg2ItxNCgqQN4HXS3bjFsdDntAbdnjyIT6/CDVY42H8i
7hckFoRKf4Su7Ciwl/oFPli2eRdzI3gFFgzr0GiB6MFGP3ZNODLBndpbPTFxpIW90v+JsPpfz5+6
iv1s14wYCkScVG7HUSIsVeBeHIANyQgBE1EAJlvUFotLguBqV0L6/EI3sDKMWZ7IzS94KX8dJAKG
3iD+/BFxz0MrMvwlNzcArYy69i80NEdiFlA2+/AKPe9CKLdU6kh4on9X7GfFM9psYb2BoQkcCiOi
reqAGlI0HP3n2PhVBAzBgS6ki9IFHPkmLsRM6F0hkJJY4SRmp237xWHAvWuJ5EyD8Cqhsnvu2j0o
eZAgTh4mMgtO+MJBn9rd68JMUClJXR1nH9m3ULKJ6cFHTquC6vL2Ko8nkpRmY7P59mCa7oozyMbQ
qTaMzTp0ljmkLMUgWJ14COpuLiQjM6u+3KQNMgvKesdVI5rfu1C1GrVPeW5lChL5Kyg03ld81lWe
NxNOwWeuqekZXfcOJFxfUNpAwaKUhbxduh9ORsWTx/scf6qCpRSXUO/dP/ThlUZNhS/B51GWTznd
BxoVtA9IUXU1FYpHYx9IvxKkN7n/XfbA+oRLANYZc/wTekLbwhgKsCfveGIzULaAX91kWlK99dG/
Hz7/5JwYZdLl9TP0JhFxcSvFiWCyQoBkukh8MekuTgzY+kRSfKVUgzSwWGAZuLQzbeUcozvr2G1p
an+gvOiRT6np1Re3QMULuT7nXhS2wX6ffHsdJ3ESJsebXskWYy499/SISmT5VY3mH8vKunwOGr/7
1hPPmUkjXNKhsonI/x9bhl3+uIOTSSqc+K5BzUkPf++PO3/pD0cyM1u0BzMgWxYJNXfOiZBipg5J
KHuibB/v6JbX+UzYfbReyd9Lsr82VTekrzEoWgMy60jQkwxLK4oHwo+XoyvLp7K0qrGiVATCFguv
x/rMEk8Hc2NR6YEQs9a3rwt/sYjYKyhQPaNSHHQf/OfWHOSG9SAQzV6Th+zki9E3kxTdps0yUtOe
CYZaAGUoZylBSskUl8cCthrkEdDTAjD2TPB1Cw2zgD2n+Mct37ZK5IeLPDKSXWswEWNnlI1HtQjO
A+oiPU3B4QgDw6/f/wVURVWXmEvld+df8NmoZ3d4yeHe2VFe5whhLQwFKKDsW4jtqX7s+vwoDDVA
NGAIK+Fj6BGCvav7xkNeN8NCqeGy1tpY2MhEtjVxOuB908tC0lChnIr0LPLLiT00gC5oVhxz3vpG
wQ9PQ/pCculb5hTlyBdSoYtYhgJ3crZ1Rpc2x/UnxREkKUS3PmniylHOZvaieQFbiQYxU6+S4qfa
Y2C+/G+RmF8tzIU1hxtpP6m/ckJfZPEKVjIJVaql761BEqju+ZR324oWhNs2Ack6YcWxLuz0gAtT
M83WJhIfbMpLjVfJqe3CvFad4REEnHEllchofxX7ngTYpid6AoaNtnFzKJN3o3c3Zm/W124cEkeK
YekWXenZmEA7WX6k3QmYgMKedimQRprsWpGL10DplWxVSJpkM3JurOZh+6zqm9MCFk6KJDUIhpt2
Sz3D8izNBrrS6XBG7ed9Xaitk8FjR1S+u2321V7c5rBv2XMLdp4s+zI+NKwW2G6A96VrErXWTJjW
eecHkHmjTwIzZx7AGEv8JttbbHkcNNJYFk4SWtabHWL7gLgp0cu9VzdHhFSLQF6XgeN1FDZg4TwG
TpUyWLWCnSl27DQK4SRP0Ct1PINThPHnaRs8u+f6hEHv70ynlp8ZYgiqaPSkZVxKjZa8KfNQ+dWS
dJ+QnGf3IYnq2IE6hm3Yd8jTD9bWUXXNvHLxdZl/xHYrnMdDMRO9WZpdFWqF637PZXfXhriPJ+wK
cTW8P3MhmQERoynLO4ZSzBgVRl7irp4lz/VaNK73hJO/pyITqVa80kMXOdPQJyI/6L4oqRukfQAL
cHQlik5Wjeqz4eekOsIIrHwmI6ihVVeNRu6tYrB/F91FwW87o5wCMALNvn4UASTs0bqHQwdc2XUi
s6UCHjoHlr8K/GU+Kp5Tc6mlVT0pSzZ4EZTfu6+yQFDnod1LEXhhcXdt/iCjvuHn6ZWOyHEKIvHF
bwKBrwpC3VnXEV3rAGzYEFAnCAIQeJjxoHG4Yi+ADJPgMv5uZqycQygJ5bh8DtfV4EhIKY/LIoDQ
ybDsAK6qFJ5UvoshrPCh0fepoielhCb21CXsVBddZJWT/Y0SiKBo9zokrunlcZGLn5ne/XoNWwGH
ajBQWFlLrlnwNr9uBeHUr1n6NfozthRiNyWTvnbxCRAPmMVsXlhQqS7B5R73MapwMYBKE33wjDR/
hnXl1m6e7Vk3J33+Z7zKPUgTZDHe2YoN/2eOQnC11zCpiWZV4mTRbawTrFUwNy1j5yZ5tH50DmVL
gIv0OoZ8ChdZgYRubpAfVoYFF6nDz7eFRVq5aOTeS9BcJCtejcAaeU1wu5TXLD/n21Yi+FJHSQNu
HxDaK215X/91+itA++6MMNDJr+/YV3rmh3Xe90hQDd5qgOFqSudpIsyYiUxmYzRrZLYfOz4WwfNg
/C1StzmjY7ryCsEih2Fcd+Oy4Bf2yPcfj0RxbOntG6Bt+RPBDbGcJ0VwqDarGOuvX0SiIrsLHkip
mfC1xigB7xwzwLxqICNnClHlomRbZ85X7cR4uFL+iRnubMn4sH+wnIS1Gy1w1XE6c3TxpSgmm4Kc
dcFe6ansd8/DILt2BlUAfYIY2dcTVFqXutSLF55Fpin9s0xUUf4iJh2k/V9sYhhdjw9XFVMQD+P5
hXzf9lPxa7mgK/1RtMX5t1bkq0SzNWhqRnhM6TxwSgZbjuUTI9Q0Rie5QMgPB6YMosRHCjgJHIqy
TaYzlUSEeT4JMm7iWfZrbGuwEgnZPpiKUmtUbuBlOkrHEi5tyu22wVV+FkCVB0I9AdJl3tJVXR7x
JWbMm0b5rLv2VXt6Sg4boMjmcwgDdH+z/ebGwOa4xUR+EgiCx5b+aT0zxgO6mSC8w8yya8fAw78s
lFXGhjwgI+x9nwdAuJxlAwg4Z0kzNd6hw3MfnUB9yL9MdvdaKdYrz8K3SB9ssw1d760CkOxNp2ST
7anKyerN/Oz9I2Bd81GTrw2GWtuZpr83loYVJCeR6NnKoXUug7IW/UAHsETekQkzbpSIWsdUkWhc
FW2aIDorE9LOtyH77qQaFDe1VXogEfUU7F3oYZ8/6riO8Q7nC2gkEL5CsNNpkdYAa7RGuiVsdnoD
qrCqLhYgrKz+vDIBDdLfkWX/6YPBes0L+2tlya6z4bxCnqrezQFX+jV9ToGZ+bCSbRjJvq57TAd3
CDU3Q2hec/aF7C9LcbQasGGCLqkhBs+t5x8sGzLYTvCVmzWyLYCDTisNuNOWvDbIys4q/Iktc5il
aSfdWTtJCCIbQPI12Vk/A2Z1kvUjliEi1PtZj76AHMeTumVI7Q/AKK8zs19QjOmwC4jpJTOCRejM
/sX0gsZ/SQameV1fOWPzmLPjJKfNL43qgbBXaDgsY2vtTyAayXNTgE5VUVKe4IEQBjK3DbJqmQaC
LkwRj9PAGyKeusku0GBeiIerI+w8ZlLEjXne3KsfSm+xPD+Fyd16NbaLqhPjwZvdt148640RlJD8
Xb1FSzl5ILW/RNSMJx8KVLMbVv8dhEsH6EbTuqTtDNqiOfN7weUsoUg3dFneot666BX86wo3RGTk
zB3pOVg3nrh0LVSl8a2du8zcaOHL1bvAmOJRvFDBvPCEcN/hZn5TnPUDCrHOaQK80VEoWcLdvt5V
81liWWzaw54Rrltd7q3xxbyGbuuflKF5+6rd+ACgbns7LN/yOLAUz7+xxteQdlpGuqp+3wV8hJha
BnwsLjwyZb4fNHgaswpnribGmMwai9JHM0sLiVG6OuqXl3rTdgiyf6+ntf2F4HcXzK+Hd830Iz6b
wGImBRnQP8MqGi6S5Llw368BG8+ZZJYSB6Ma5h0SKUlZ06ssd14Oc9il0VMkaBL4qrUmRTbHxwd8
weBZlFRjz6OO2ikpSHe/HHPl5pNjKQiJnPP1otQSK4VqlcaljSE9JgcmgvtQpz2LUirskL/SiQEn
gzD1mjafChTiigcwOcjdfavxUmeQ/hHwhFwGUldP+5uP2j5gzADpUJ1lQthrXLIbpewzgR1JY849
i4GIyVcJrMNeBiDZhXUP2J6wRsi7JmWxLcXNFY5k/Vsls/hPIYnHhuVjhsQ0awljTQYKXlO5hp2y
tI2Dj/yFx9TAXvZzz0xNpMB2r3+7AOLFsetgLlcrAmTmX3OkSbdc/t45cV6Tk/zqr4F2mpFgOwcA
Iqyqup+ul/ce81whf+iYgdj5NNgEKKzQO0IN2CWtJClh2DCqr5sGPVYCxVhD2d2HAx8q8AiawUT6
/V9LQiU1yTNgne6mbssMDyDAbX10mg2ffRJFhubHwZjRlYNDGzg0fS66OVKsanoTjaj7F9L+PRJi
cMFZcdSF1eLicCZPU6Y8kMRi3CqrQX3iroALWuEbinwOyHAHqNEZjLpfzSDBJHPXsY+8d6dgD8//
z48/2eD0SbMXEV5sC4Dv0tHDi7ohjp7a9H5U7n7G913FxdSipD0x/JciQN2oRHRNqyjjyVzHaZrN
MQuJ1hh8VWsLFfKf9a9V0QYEqQR1pLjOn8n0lAc0//NCJd4TqMlxPd+whBIhrPaLUwMFHBzLAeKw
p2+/eBYgvVD5Rj1v+LahjbLrdpNvFkVfPoZXVXlSGQPMXC0Keszjbeu2+vuJJmvixyHTVWczYC32
UX/QsOIr60SqYhMdDaKWmXAaoMjH2vc0JHd9GoetpZv5j23E7C/HhO8Cu4eNSEldXmK0VADVwlDv
/osPiYwFRjCGpg9xUJlSJ8xZGjVDWZuBOkjvqDJ4J8ITK2i3cPAvJcxDFD61MFNlwGjzqFejWOOJ
odsvuWsmRnPf3XqmwTIHY4+IFBj25YhLKjZkDYnUWpvAs3zms0FDC72dt/Ab7RkWXyrSp+vQ8p3B
Z4y/lW5wkl7rO6T+NzPqzdYRiI6vMt8gy1HaODJEzaUzE9yuRq7MaeFvWDxNNFiV8ElCsMsbE+Oe
gAJm2d5pjhmr0qQl1w03NVdn+CWzgKT2qrdqYBgYHwWDjODQOeN2m/i30ZMywgwKO0BRrNPIxP9s
zKF46sAWJf5sNTn/vqZfUP43JhA0QzHcTqVxZEJlpPuUZpsAhHkRYrx5+Ugcwfop+U0Lr5xDz/Io
cNkNNGJXw2FCJSnCbSH2TfpPqUMod/RtFCpG8fJz4Q4IE0RNtwsEXztwCp7svSXKgsEYjsHNDIRE
HK+DsRwir3Jyt/FMOyZuyniHaY+M4M9DBFMLdhIbRQjjuekAArPV0FaJcrUJfMIUUIcuecX2TrjD
SuNxAeO0IUg0LYDDKtNKsqDbCzv7WedbVr59iJDKbzsoyqAg+/8WS26BpysOde6gk82JxmO/y91B
89K3C5MRn+BCVjQvZISBIh/yV+f06+kA5417JZ5q9M5Bjs1swy8N4TIgln5pteP8FzgcRGPxuvgY
4CVWs+0vEZc1fxNlwqGBjikM5WnC42UB0gMvWEHCs3WQUtV5rluZzK4ZBcKhxwWOMrLemV23Seqs
prqN0MrK1i7ARzg/Q9jAhWhZwinVARRGYwEvJ6xe87AhirqMhpl774xsCiKpPSuQeEi6Jnh/hGJO
jet9X055CJXN/3swKL03dmLjfApUg2FKlCjZNirFcF9eeHufJhA24PVL0PU1uGHX3BIiL1bH5FPe
NwX3Vcqm0wlZ4YrTNH96f2ckAtw8GiThxIyW96xGY4q35wym3ZOiuyrjfchLV2qN1zv/SADbaYwD
LC+7/g5boIgx/p2xNWuY6nc5uGY4cb27WILvDiuD0tQfuU6UFqUDd+wXyS0HPpGIUpDEp5UxD8NO
7jTi2bLYB2yYHjn6lesD+Xzep24jXmwaxwP7V8Q6pPoqv2l8ClQOrEoZ2+4FY8Re+scs/OmVnSFS
86HBcmFc0uGzQPW5l/4oHUFeEBcdymnXa4KkypIc6bQL1H+al39ZWoGMHV2kHkoixm/avifJ5dt8
zEbBso4bILjAx7CWOam2dj1/hofyK26/ssWjNVS7jAxUxbmUzISaNN/DMqLF7qoQ7KAkM6ek326q
8tBuRw5inEuDmoLYojpxCXI+zmtwokK3+o/AdTeYZ4o/Rx7qHa9XoYj6XLVvim2TleHQE4sSQg00
DgpBhqT/+pCNAGRXfXs6WWcTZOA0OSSUrVevUp7Y0NV8k8mI70nBXdK7/an2JLSYkdZCJiVBAey3
Qv9c5bAFASthQuISBwAZP3cDfpms1v3yB5+ao+b9JgY+RdpgAVV2Il4H0jTHghTsB++bXfOLmz+g
5twq9/VuaAl9ojwi0XT2nmRwUV7EhXqxJjeG+Z7bZj09YfpHGALnuz7PJFzlNVcVoKNMIx/noAOv
vwnCZ+orPpAuNDytpPHbS/3NLOXs6VzxOrNAFKEhFn73bbnHNbTbqxAOOIw3idYsITr6fArOIfdP
V74OEgxXK3CKPO4qjtVXCESPuQHeRCNj+DCXkZAWjsqUflmc0dhxC3s+7D664SiZ7wecW+ipiO4l
da0NNBQ2DZCgQXB8F4P7vaKRwemOTnK503x3nSrlFDed9u8+zDGZ0UAuVspRpo43tBqZI9CUWJ5T
4SFMBQXwUNDLd5t4I1LNfLatB4T/9ONkHDsFNteR7Wy8HrJMnksnmO41cC8prTzAiyLGRiJZRId/
huvBwlrG8CSfhksCNjjr0bSARS6ndpAOuRhCavK+V0Fb9h3o4+gHzrNKO8WIhgmBvtzurZUf4ikZ
QWrr8XtJKMj/VZyvQ/wUMly6tJ4xdoAbM4zH3W1AXj4+s+VHQN5EU9Lm21G9E52oVK7+qRwZFoXH
b4xmbTsGY9yZMoqOZQ0loksEY+IdlDzyUIZMobwMOzixxGmcWpuwdTDP9UoyPvkciGkoNjCaDXM5
sj4/hxzBVhmLOT1GbNr5pNtZNSXc2HU8ThpUL3/Yw6Zs0/X7bBw1iRFsWh8QaKyD857dijO3qhyq
li+98myc8OK/PNmEd8JY400WoBVOxrZ3Jfh8oXMw5SwmcyBvBSB2nZzJp40s1bX4dXQsqFaSbd8W
f2qI4zdtqsnbWQVHYczwUROYztGG/ptLtmaIGyTrLdrGA7LzdTXLjrP+zb/OrwrJbOOrWuwPH+Di
uw3N93LxtQ3Zmvy7eo2ptLVRnniB8L6iLnjRDGlmmD4rG6hV//Sp/31NcBH7WsXWyZnlBc08a8Va
KSixMhLObapP9QtotPuYDWHy1KWUrC3K5XhoIKHx7LDpIFHj7EyBqWXXL3gSSjhSAM5JXVl4BS64
B63rZoJ4vJKQfShPSbbDquCIDFFheYU14FIPGsM3l42a/vkFJ+3vXtx/f/qxlwp8uKPXyFvMGGAr
5Wiy+kLS+4sFfpMhBosoRLIWUeDuSnDy3DYl0BC/UjWlDKT/RIj3gbCUNPW/HYjKIWNuiBaP5xot
gonQattMlvopJugxXYhn++fswaNA9uAjN3p2IPFir2ktOAr8LHU9dhAZwme++nvIJzZhdTtLtb3m
Bpad/Jm+IPmp4aeleuA/GXQqu2Wlk++B6UxMBpadHImPFEkONMXqD2lBfrVnh/og0clrn/3sLTc6
y3tfKvqz3nc0LFmz1xT0EzGtc3k303jDJCCeoeFfNbgCPJlxZwLYwRq25Jd79rxKcVXYeF/CwYTG
7nTeo3rPwhMigW/Up6wXR/wCLFBiyLwtV+VKtDGKysHx7JQwHWuz2PPrEtRrwwO+idInnTkHZ7Zf
FVSDFuWDkxIqO45zA7z6o3UsUrukHdnANdxyNWyDmtq/PEOi5ob6hsmYU/vECqEh9F2KaVvI8k2/
f24PBHuQCaLqARYeDYNcwb+0tDc3mD+AOPRUjfgSPiC5xsZk15FbojI3LVB0jDNBDqjtegdFAAb2
RaQ3VHwsDGEp03ILTxyAw8HL7OnjiipKpbFs/mwpp0udbY7nBIwp++BEmam2lP0m/WRXaugttStw
pL0zX9eJfDfuJaqZCVgz6ai6SsLA2zKwbwEaxjNy6FrKdS3JI1UyXbWG/5yeuiPyoMS9acDFpZmJ
XTB3DYcQi1FHpORQt1eTxXZ0L2HOLP69oSJeYnFUqcT192LHhMkmYKk0xK4WmELiEdOHDp/ted4r
gBRVy+BF7lTa/pnrQJcbtwIRkisIZgz5jfvBrRo2GOMS2X3gCcTD3l5MjG5ya5VKv2M/iZiPy/RQ
9PHViBpTuYF2V7W6VEhN6OMxDmPl1NNon2XXwvK/rm08dXzoe2MBdyFWAYthYy1wjVwi02xsFV7e
matfEuxyl8/IR0e/IIMBnB0JcoRu1Yo8aphRQAPV9c8LhK1ZvqQq2Zvy+WEWY5QdEGsht/0Lb+1h
xjMCiLE197cstGmQwSb8BzMIGQ8Gj1xgTgjRNZeWF9e+B9KR9m742GQcsyCwY+8G2+35j55DM6GB
qt3hQ9yDR+Ifmtwyp0CI+/WGHjQFEpljbI9w0HiwOCwH9xVgfnkwYQuQIj6JTpGcPdh3mQvm6clh
/PcQofFzxPrN4BZAaCvmoA739jzT9d/JRo6zDqOzTtH2mrfv71PKfbPi29nzPDQyzUj3faOOpKj3
HZNvDryIWnA8rxNlDJKDxD0zEynnecLMrmBKZqoogq4Yzi5AjpzSB/qVEqKq4g5ljp0j3lJiy+5f
tKgarwFSVBYttav6JVFFQ41C79UUhOlU1tCnNPT56yDps6ZelII0owvfC/lbm/PIQsH+m+5BANJ2
NF2s3/oHm4F+6Ml9+oRGHgZXuWOs1/kLZn3SroKaEqyg6wkT2pqYenR5D4eFx04/0kGT8a0CHxCB
zqu+VJbsfGCTfygtloUMJ58Vj+BCBLIOyjv1SC4r+fDUk1g1ARzYXWm6fUQmOHMt5p0K58qEuk+a
BMomZ+LZDwxSJeNHXBy/dsKlK3w01Uh79tqBNdyaYBFDTkDnbH+rgt340KC0Q2w8O55eDEk2Qj4h
j8xKCl8MNOdGssljK6ltBLQwrLFi22KxhYIydO3i5lkhDi//GfcvJKDnI8NRor1bmVqPneRDOpZn
BekMH7j2eUTQUGTVYCu7eReJXBxHUUoSUEAI3IrPeoEvhe/TlmE0zyFqNLHo71/YaLgbxWsHIbUw
YPGvZlZmrGNIVHJGzlXbcGRldhLyIrVh82s8TZVLVdD81idd7K8oF9AUHE2qxbGgNM3nvWGTjopy
UxDuAylJjAPanPblTR0swTPd7ptELxhX9JnVsxigOvctE//UoHOb+zESyznbymCMo50kBH9G970U
Vx+zkRTR8/EZofR9PFTyuEkNxq9OaJ/oDZmKkKs/OpEc4JXKS+9VmZ7VaadRjNOuTKfpoe/zE22m
8F9erZyLKLIdJpoxpcDz5u9zH8Au4ZPexUkkM0V0jb45d78sFQ39FZs/2HaWl9Ayu5vt5ArzUOBM
fUnuVMDG4TWXU5ZjPOiUCYVLY7kaqf737xwcxTjEoLxIN3kKtW52GxNryB5fmPx+euZBTJ9sNs2O
MLjshPQqXBNOT9z1LtGfvpvIDbFNIae151bteaZOs1Pl3pirI1Fy7lOodha0MSHTiYwpD5xMA1HV
34aATM4UAJ4O+BTLOAhCfYC20oDgBttytwhHIdp3xwBoLvbq2RPyITQa/cfR40GT+yRQ9uVKCclj
ZlOekg5HVzaW6JKMv1woyOJ2S8BQzMUWjc7eoWhg5tk5gfgCwfweSwTYc2uNYcruJ16cJJmZEkdP
W6sVBTp8JsYiry5y7Rk/RN3vHu7GVKrlu9y61VkX+QuaWg9PcIpKsSaId+sxBLteAY7RiF+MLWBP
ykAVtxFz4Knhx5Y2qGCFktfHSO5o7heJNDo+ASWu9CSEV8P7aeTV0h8UqHoP+728rtY2OmUK/ZGJ
KQwHbSkVuvsZBR63fXEhkemo1/92gyYLWyxOG+O68a2FU5ELLyihqz7SgvclE2DVqlSYWpS/1erh
jDHi87Pe0c8AkOetyDPgZAmJvtJX3S2BtjjhuZOEjJRkHaTWQ9b7mAksxX3Ftz9lvPF5OoPeWuNZ
T39NV32sxNhfv5NJvj/mwQkoLAgAxwVV7+NHyKpUWRWgQU6FsefOWJqVxYPjxI02XB0wWYTyO+11
ovHMqjdC9zvQjxoE5sWGtPTUi1XG7Ucu6OVKj31HLLHESksmz4Vy/xuam9OEBWCE43MRTq07l4ng
6qk4VVCC165XgZ06Upjls1c55d/acyuyUGZnpPacWom0Fz+/DQMg1w/VqQlHbC+mWJ2t3gDPwEaU
5E7NvwNEcLmKk7oLxRAq0uhnBQIH12uwM0q5ZOJhqE2BY+uvk1kNa9N0t7BNrmc6KCsdpZtwqt4s
fpap+3t1iiw0s1w9b67MdSjm7gMTJ/SXxYBHYFzXNgDvyh6798hDmFW0JDQHdcvtw+AHxbW14aTU
Qou9EaKQPs6Mm/QPqGTTrcWpTdGlkiAbQU9oWyrWgIYEXkCJpOcQ3wFItjNG3ZGjJj94qr0UssqF
KXhR+Z6GFi8eAN6jlpWI1rysU2fmpaHhzxxBrWaRx09zQtwmczloGAcxtIWAMRQt+PFvb9DVvK/T
PyH9yo/Yh/fL/MXw5RZEtTDxjJAvvk0FhnvMTNVogC88jEOO/nK9wMmgDFjFEKBeaY3Piw4I8TR6
7vBiNa4c3r0qJfn1Z1DuaTsig3i98XsOVqDL+/DO/gIa8lOZUUcK9C3chKxKUEGcHPqVLnjwl6CT
tm+XF1Xbk34gtpZwa18b9MOY5/xReueOU2ZzaV65g2W1dKqqlydIiV1tco5+xsma5P+zZ9EikpRw
JL2LCE8R0vy0vcPQlvvBHsKrWeUTGHU/3g6HJFbBvsjKhL+P7CvQ5XTnbxazYahdGPAYBzdMrZkw
8OMcFb0wLVce0cQJj5dT5ZVkryHRg4Rswz5kyYZRNxHUT013SmHqx60PR5VX7QvNHfbiHgp7vjej
IB9LQlq45T/XIiUEbe36ZwWwY2T5p6wAloRee4PxuihHlO/5kC/u4AbT37sR4+V0F1w6rHytUwJC
fJ2PTmCyCThmCoxIdqdJlEW84/VsWtUwuPQyUqwuXdc/Ki7y2C7jnVS4YucYLWXszvwQh4lPq7vM
PHer7ol309kU7EDgIzhszV9GK3qkyzxl/4ySeUc6YkSecPn13lHoPGCuoQkCaq4b08v1i6goZY9Q
yKx5dXQvhKuc++CVbnKztxcXF0TIt0TwN44+Z7bc6iUx7i13DPlqx+gqjpCR+VLmrK+XsOr1Yo+Z
C9IA+he28Y311mwScKSGiiMICS6rH76LJBiRMd9/vEluMHYZD7+WW7euVnOH2q1b3yMEa6JVFh8v
JRdmYaH5eeLwc2KXg2grYZ9Bmn1XP7IO469YQo1Hc1RUP9amyOL803jFYI+lH3zU0NgTv4qFlwNb
7/MTq9przV0RXEsm0meU8wDLoYSftTBVe35C6d4RY7uTABNp94YiPE9zrRdQ4onvUuNa8sR4a88G
Bu97l/HiHE1iW722PnKtez/486HTog4E8BNGN62KIISzZKpAEFWYMsixmGZGo4xgbgfZOWvMy5n0
v6HpwaQZ3FuKjPt52NC2Evr58u7UEIH+38rR53NmxtCLXwozO0O8b3AtWryYer7Bjc8Y8SPmckzq
6NgPaBmoVg6UrKmeNPqnPetHQgpjs+tjwwGW3m1LiW1bwtJWDoMnV0Rtt1kNOjTbGwGhtjiY3hcP
dTHXQlNZuHIsZ6JyoBa+E3SpO4J+IvZyOm0Z/SDQNejz1AeT9INZqsG0it8dYS48ALbNu5vxR6/i
Jv/XemkEHI6HVd4fxmuBRXK0rMHjqUfQmfAgajGxPLnjLwKow8mIRrh4zmOLrRjwT/AU0hwS7HJE
7j9VS8+9MtkgHkoUPf2QwECdp4uteDiR3GNSuAgk3zfMU0dLi9qvbmmgkMvHI0SvX1i0QPwWBczP
MKaw9ji6nPTLo0FCeZ4O/bmU+Dqa0zf7SC0WxocrzCTMZ8jfWw5j7oK3xBRKA6omTqPva3c/Ueet
VzIaQ0kE/R2BYjgx1LZMI6ESw9En5c+w4Oif+I+/IrQNI/HqtsnXudX5dfEm96c0Ayw+pTr4SzRD
GG7Wr3l5cwFYCDwYGQ0mDX70dWZXN43cebI9msjxLnoWtqrfJYdEA0kV1ATFrd/235CuODXi49e2
lqXmKjPOmlB/A/pvwsFgyORNJPNPqG6T4vDHwt4pnDRAVs2tT7YgNBj9eaQFI38EEcCnPC89i6fM
lwn6nPIZNI16q/ZOVdXkTSgQmGYXEnmTzTN6TAewhQ40wv5mDqyvPMlqgspyYcQuwm5K3AH/WqUT
9Aoq10Ed1y9adZH+HLRAL/iwM0OPIH7miQB67rXxZy1ESnKXKOzMtfiLP/VRckY4BsT9CLqlwQB5
0nWFHIyokfejWjbkvfVqKcK51b4qmfP6EJknpOJ2MndIaiR6CGI8gTTz1sNnNANmdhj3QXFyPAly
FTfPywmqQXqCSwZFOBrRvaQZFQidxfKsXXYtyrpxuEQXsZlckOhoySircUSretEPgyI+h+VNMOrt
xtIB/DTTeyChk0efEO3BIew/vkd9gRFMcWFl/Bp3FEbafau6HU/KBu3DMgdI2etaFAQIrF1VhFLX
lLGLD+Jwb/dZ5nmkET3bJIhkyRcuMoCle6WtIHjdIha78ebDSMdQobPUk8+0GZpZn7ElEAe43qD5
O6ruQmY1RcmIllhkGVJ0SDFmBY6vwCjU6T5CIFQw169MVHwYBLP2QsT7+pqJ7EQ3gZXKWZnQg9XE
ObEwqXLM3MXBaPI9B65Q6M4/nJH5VJrWTf8vjLqpwAd6p198qBylpvpM73yAwpJ7vIwcjc6s1tez
ubotAEHt/2sag9ybNlTtIURhISf/DagnB0B7SrK3qc5aHWwEFI5cNyDCz5abPqsET5KnZCBwhmSr
PlAqDUzJgW/5yLjAeVNY7VK72VJVKEUCCjmnQii/QvSMfCGlSdyrXJwmb5de5qmYh8c3EYQYNhlk
d78tNEt9csz5a62PfKQGjGD1aU+rs2DE7NqpNsip0caP4eKkQdsoxZE/d/imPBM5xPoNms/AHE3u
Wr72LlWsYH2bwmQ3zPSydrgFEGaifyAhI2JSFwmmiUfHsYd1wkSaZbYhm7kfWRZMml6gVKo80FT/
49vQdMGk7Ts3KrtwYLkVyMGW5znYUmoxKuZkMnyW4IxJtH0hHFUL80XnkSnXbevKB1uYHMiT55r1
VOAQg34Bl4zErXlQgM5PIM0664mAbOkRjH8rFspH0qtm8wkXzSEXc1SNJkjwDIgSYAmMEXBJtN9j
Xylii45+3m0g5CVKvP3IAcJkY2WuL1qTfBvQTWjPFBo/r7mvIaLZwAhdO5RBk7yPsSf18eHci22s
sciBa+7YHGdeJjuy3N5t8NlcWcy2M9QSdbODGLCtlFLup+UhXshWb1tWJMNrJCxKv8z+p3Tqjwv9
cnNgcLu73lBbm0hzuIBhziUNpk8qWWEM8w/62/DnVWTUijpOKRLCAFBLWupo227KPacv5/C+uEcB
NfOWjxDNZUPqS/EW6bzZ+3IyAHUlWYe13EcssqHKv9AkHCJs0b4pfpF4fu1aRq6cLh+dLr6aplT6
SDpPzOIZ+Ju/YPQ6O1FnemQEfbrVFtzmAgXAadOC+xIv5d92EuGS60VxyTg076+q+eFlxyyN/pf5
O1USHdPTmcqTvsAeWOSkFycKiqCx7c8qn5Aqy0IKDHcY3c6x7p42N8CAoTJB5KMEq7Xo+38id2Wl
GexD453hvUM5GzdrgCI2L7qBSec8owSK4iJNpbCVKsJqc96/2FIV7ofphhXAfnNiG1HDU98Uio+c
mqNd2iIpUSE7d2dGxUr6bldmtb7eobpRed/apZvFzmct7dza8Q/J2446fCEiNCtt7KWx2q15W+kP
N0qvUDypePon3y4rXT+gYX013bvg8K7pzPqmEuhd4P6igF8JK2Ti4UcHWD7aAcCGJC54dIm+0TZk
jjiEEU41xle9moOMRqUjrvyA5ieuYG+Pn36+G+WNGIOlJpQ9yGQr2/xapd7P0NSdaUWUKi7ELzqR
AO2Ou3tFmYmiUAuZU5G/ADgI5U/hzpiKD7+wx1aUBEFzGEg03IZwPgJj7AVxEwnm6ef+axc5vO/t
Sa6sd8sFh/VE6fEHtuOT539SFGMA700PLQiy2WPKd8pVTgiOw38ITGm3B9ITwdlPGcaglIrtsiWp
nPLl+U3JlWTDdKaMLZDYtyl8prr3KJQfnaH/PeYTO7LEOAtWAGKTdgEmJ52eECuA5gYRVcvgNqzj
dhgrthA8Rt51M5v/TMvpu8ATBAj7s/6HTUi5BvXqcPqxSo6vm+dF+cBlXa4b2TD/wKc05lISEO5d
/PZZLXrM8DpD/PzE1uzLifa9ZcJ+D6lplgIdmZRuLok4zud01qTJIJc4YUpbOJ9P2nrrLcXdJPgT
dFWPb9qWCeYtaa8g2fDMty+Fw4r0GPUCfJjsiPmNiD9TQELQ9Wfh9sj/1CPmObNz/hgewgrCa+/M
jhjpqYwODY25wA49xheWZpvImNOYP+CfCV6KmIBZv/9O2OG5VTMmtaX6zlEbKg/3OXO9/mdeq/8q
/hlkzXxzboR/xboMY3jAY2YYVNH8+0X1JWllXorXJyWzwgD/sBZPrr2HqfHFX5T5Uight0AlaX0E
gkpj7FZjdxHC50CmYAApItPxSxK/PcAiSN2RjTNoymniMwpxkcaIOwleoHg8EaS5h6GGfrbpzYrX
1R6TDB3BPir1Tbr3xJZ0zoOFwozR/o2ZfurZK07MMCBRPE8EWfj5mewd09p7/x1TVmoVzg8Y0HjT
mo/4f4Q0LtPjvsKs71lhUTqnsMVLip8Vj2QSS0GVq/MN0msrE4crqNa9T72UzHheTIN/YqAW+sIQ
gzDSTvgS6uzAjzba433uoYGuHBGHwuBJ+lf2PeSFGvfiBd5YwkUrPzBwdqht91q4Yo1ma4Xbtxul
mPThPszN6vFaHa4gPdnxkohydhzpohxXBPLt/RDfhtUv7YHHMqnjT5oJJ0ypx2fGxn9VmcHiUD2F
/Zp/P5mZJFakV47LUyW/zn3PHgvBtPq2rv8LP3/NG1YF9tPwWGHmi2+0cpo4IssO0V1T8l86F9qj
SDxvHIoIZaXmu8/c9n5aHUKniR+ZqYVmM+10SE3wtrsLxWbg3hrtHuIirrHF0H77E2UwmIYFA3S3
Nbc4MXHym3hrJRBMkw9bJWrbpgPBIo4u0obvDKqBtaWom3jqoRenBhkIHQgx1sKSQvGH2FhrMLJz
M/OgXTJgePuo0fLlywUD8pQy35BFDaxijaq0WtC/nxeeOt9oJ8G0uGhchNpQtXwTCWurDAj5/DnS
M7g0Xm0TcuUINZgnq9DBeI5rdj4IlHVWYb9aszBzHNxOyDa2qjqCsQkDyF25wYW66Pna1c0e3qnp
hy1gRxYEqwnP1eMovAc79Up/ufCR8rf8FcHIJob69oqnwVI9a4KbmE9q2lJuWQThY0oOYLJYzfmh
CL0vcSmPT2Cjo71PjhPttZo1odt1tt6op/nVDljZ9WJFL8+3dancHTZWkYq0g4rN7hXwmbfDigSu
mR0nvcMIgFMgDuWFI15dNASrfUdaoonJyr1n8CmE9PYdSC/U5sMJMoZaJw+V7Ck1Mg0ylE2g8LRX
SUNFTfGrsDR5vgK5oPcTokSMoBxHBYZmuE6kvRkTkjbZB740Wc1sDcQSJOont2xjQD+VKjCGdbso
ruNByVZtbpcQPf8eRqFsYqrjIjOXo0v4AAOE7Zoz8N+pZpW1K7Q4E0o4SH34e+gra5Byl7oMsnTz
uV5YlJN61xjWd2hbCfdHGpeGpWvld0gRGdjPbVumuF88Amb1G4je24tZ+0XSkIZSp65UyDqWUnl0
KNzHKosxsgoTelv3YZ3P3pV0t+vnzzlhCz4llHLx4kWsD0i6IzAQTZ9b8rogV+gK12aO6B3dQw1C
1JmxkvIiMW0UfSxK0LE183FUwVW63sV+cFKkVuSKT+MRnUjrByXc823PPbtj2TKyopdXp5S2o+Wq
BNxISlRN3Dh2XR2benrBShvfNk27rfUuPgZMIr/aH24l5gVLS72j02c4DHZnAW4B/MiKUd0mbC5S
EhPMerhlRcAM7HD1I40dUzTZjtdkIFmAGML3OBTMn7PAdZIfsprKwgAuvxVcrWpBuJz6IBijnXU/
+p+jt8CCqopj+K76J/Swf0X68IW8yu8PzIwQFMlF8ah+cuk7YJBfOEpeIu0/AY6r3P2OjNIb4NNF
09UOcXR+VxFwXJm8GvOTHtwCnApWRETG/7bfBFeSz0JkdWGzoxy+m6kEd9fh0OYxQtoD4hbxu9FV
x8NDdosN61sAdn8wAcrDvtgEX/9U80o8CNfK6dr1uMAqsTKGO+OgBDmWSSuA8Qgdb0BJUj+mB/Ql
vyz+izI5unvScQGywjsEYXLSX1ESmxvnCt4ROuOaPTnm0BfagV43yxoXdmRhnM/hT5HINO9X046C
Y3p8fC3bIZmd4WDZdK/M8jS9iNtl5DLI+klrpdp0WAkV/4hA0Q8tc9uKSwfLLY/4s1V+q4tP2UwP
i8eqEixDU70af1TEf7ZsJb0PpPywGgyCBlrGm+tHrjaBLomBM6Zxotg7QlT+u+oMlKA01dfak/bW
EnYKSA1RhNogur/wUQVdFeTeKo8X2hmLlD645XLlAUlWlBULvqwMmLdSwkVFSXnqjUsWv9iZcN0K
kpJbLN0vlaWXiGm8mqsXDdfkWvTRZ1hTt90rW2NiLVQAdRYvOSXuh/h3brNsFjrjeEidzQFTslu3
YdX3JcvJa4rjUZKsNDYDoQPb/MIhGJsHz/m0HwZoJT57NqtWqF6/FFQV2rET+3JWyzy1Z4CWfDsO
WDiGD84dX9H2xYmFJi8JAKZfZy0WXYfzdg4I1oLr7iR+NIvGtef7Kv7eoh8TT5JCbKYrXGqEkp6r
zmOrodnRKlBM1V61Uj+qtsoYOTuknq1CL68Y7KMb64Us9f0F0X/mXPPuG+wyoV/4PcEvfVCCJU/2
hLwa14O54vgFstzyk1fVkUNsqwMp/pZ8yKp4nZNsbJjxnd15GehSzljIK/Wx6qsOWEDceOFBMRpC
6ZqQ9Ly6jLwYn9t34M1PmhfKgXHCgeCMFdXm2rLomINB8fsULqP4mduJfT7Wg2y6i2lMjgqU4C9W
WfN7OoZEhaQt6NLdxJa8SV08wc4BfiJq5DZQmZ8PYcuTZwdcibifrG0aSbRl/jf8syNtvZdPY4kv
SqundWXstLQz3AeDMZGuER+6PaGXA8+snw31jtZJDFS8qgEWbh7saUX+0Sn54nG0GpaykrkMfY/D
LBWjxkX35y+6S+sHczPYkrGkkgMPZbDmqTKsP9IG2k6JOQ1DmnBgqu7brRAI6B937Qtyy31Z4LWt
qR6pQa0Nw2aAmSrLld56XggAVXmwfmQxFeBZ/kOa5D1YoEO3aF43XrozRtBdgNOtIjvuEV9tk4nz
fu0IPPHmDGUbWDilNSYLgyCLwhMVX1GMLaPtlsqJCWvv25DnC90LLqKSPTqdQSklJU8ET+/Nae1E
a8fhthPyU6PQ1k0oSblhzU9bMZwxPjDEo09RD8xifEk4r4o73ltE8HL+trBfMT4nPJu+lOirR2hJ
0DCHXVyJQIN/1xBxcGnInS6PJSYM6r5GASX6T+HSRbWSieHQy5rk6nTOglhUK8kAQYk1ZIJ6dPhx
ou6SeA26wNwsT1ecrwNyXu5u6eQLF+alBG+mEA5UhMrnIK0E7fwP7vVSSIOh7neLgGs5YqJuobdV
7JA0GoLMwBD9FO0Mfbmr//2/Zur9RM2Wc/60pcb736FUdqXcMaZ1D22VaPsTinpAd78YSN5iRMNR
M+WaNQtiCz3Y9ga0PdnI+Uo51rqOgRPO66+XqPjFSiy5GvEpoaolphcDwmSsTpZpf0kxT+OzphaE
F66yVgDLzPvfYH8yg35qZM657kZgMN38vy1nn5aDjddtXod4Kiz815OCMS4PcJ36AajXcrgv7nFu
VhPf4IXRD9BvE61cEu4LqumV52JiZqBLRc5yTw08iaKddh6GamTc3OUfufCzrStEUnJgivRrPFSQ
uY92tljtGfhdhmjfiyLnveMIDj/8u3dBiBwR0DahgnsYvn/YcavoXC6vNf7Ti7U64HI656/D3UHp
/dfCtvbPsnCyZ2eLYf6cmbI/XMBw2S7hUIiTirmwduO20RBjhFkmtdWNZvnGuSzlcBanxG2ghaj1
YgIy4VCzGwWtYkC2jKBbflc0b3v5uHOV1rph/wQoazVsQxFIVuKzb0bif8/wI/RbOAqwCFTmiPcv
IDiWJ0OPO+Hn0DZvOgzlWRFjI4z8+hJNi7dejZsrHG2x9AXcvnxlWY0YIlKy0wgBZQTUFuVXxp6C
upSO842oSz0c6O1/8phVzbCzKNhziTeP4Y9eLxAuwIjwbKK+GXAS4igKBnYHX1lxBgQSYb5cCbIG
I2gY6sqt9CDQemshiDlaONpYD+hsCZQKY5iiIrzXHaA99k3eX/TGq91NMp6M8+qN0bB8a+ZA/MgN
QgScoKFtHv33mwhuJXhL6a5P4nqMso3RH+oGgAUumpXxFpKCpbdOUg0j53mLucPrF0mDeyD+QGJr
Md41ZtyiBgdXKrcdE48awS70rhQCTT7HD7IklXFYaxkDeo7MMDgQzErNNA210nMlZ3aTAt8uTgx6
VcfwZ3M8jx/hgs5PeGDt5nrSV2Br4bYhkQouqPDYmgKJo4DyXELSU7zSMwfNMT5w+4c5i8smq2YO
fhYf5iRFecPtO08ZE+REhMTqOrCqZZutrko8sb3Egr7idULtXHZFqrMesMDTMDGWvle5UoWB3rda
RksdYf8499zJWFD5/YwkqBmZad9MCV9UCL4J1DSbJrKH2Un7CS4nsjZ4FkmO/edGHi4hzlyfCjM/
YNoeoopdI55IgzsbWkS1iRZJq4l2CaraXSgI4iQqNmGobsBBrpbg06tSMlHvQpZbzQR0xaiClJYp
0jBtcbXYl2gU3P0+MwvoomivRCo9YPzvVEKuxmAW4zd0tR+2rAmYr4GacOwEm64+IZ8UvAdqJ/ik
h71ZLqoFFzTTf+WR+l+RklHQ6gpku3OlPbYzUqcLH3fmf5P19R8ZuK9Gy+i5aRhb5TxfmUE7Qb69
l8vZJw538yvVuRpup3UZijj5v6EfrielvDGIII/0klhutGS9SIXkFlFHb6U620uAYdQ+NNJR1Pu+
p8ykw2RjjS1bUAY0T6D/FP9lSp/o7MFeoPCxSfkK14WTf/tDZPegMj31EtyOFXdQ8u90pSFLsfFG
WEShyJUH224fqlMSlXNxqBCtA37JGqgEkR2WJcG2pRkbMXL217NNQ59cEtAl3msF9dsbrJcb5uDD
UA5G46KKcP04jL6lvP+7g2kKHnWgMPDrFxoxJJuMuGQeRlRCfalOIT7a2UzNaPy7TLjsxXnA8z0u
tSAuSpF19tvv//K2fOD7Mm9mAsRGcVe64ANM9mdIX360inPk3lMs194o3nrpf4wyR5NjfTlgHsy+
bwGOU9orau+PemDNa+FEiB+f/zc15+enuCZsPw1jeEeCgeshNN4cbZMgMzOviIvW15UCNi80xkFh
PZCriBbmYwtVm7w9Ea/Tn5Ib0JrYjV2gHTldqPHpI2AFpLIoNRGyjur8gigPtXy4DHsKqs714M1v
Jl31gGfN0zyrlQEY3ou6o0RSfPk6nhKbOesvtkpkubLcSWJCQSlE2hTgfHWsdTDG6bT8kujk6lUd
OVKIIVHNzK9l5+K2fOHclsIiUwLX48HDi+sl9iyqHNXFceP4Y12lEcA3K50A2wBPC2uUnqLfQq2X
o2pgSZC/BVLegNL6rAyBKCWppuPx4GGD1z9Yg4TPr8SvLpn5VU74pcdpS8MJS4NuLtjHi7KwAoNZ
oVuEwgKiIIS46l1qlLhsLcWliKhdTy1meIy21t+MSAXXMEeRfEiuTMkpbDhUgl5yQzyXc1pdIfpM
jK9A9Btjx7mw1KHuLviHH6QebkKs95FJs50zfC8H9HSbre5+xa4sAAGPk5ZB6jotDs6TufbRu08P
gzbCtOBbR5iU1Fsh+pzEdthLIPMWnKNzbIschYhavdHJoEMyRti5Zt8//OhZLkk0EbUVKNJBvY1d
82u2ngVV8wBLdbCa0LD0NxR1GshAW7YITtn2ZTZWEhQPhxK1torOJxc9l5pt3Rel3G6wDrKBx0z1
oMqbseBcPc7+KCw/yH7be984/B2D5hEbIqwfarXVyWOZ9/tfqRoA4qSDzIvPB5qQrOAoDqY88Iuv
PHERTyUtdbObBG6kotZtBgHMzu0EtIG44C+DlOSowoWV4jAn1QXFSoQtpALZy3CLRc1g4NGfPbZL
O2gdeWlHoZ3urARL9tWjW6UFExAplMgcFmI8lYpLbPU+7Wu8ON9oc4lSsldugKQiElmiV4r7fV0T
JhFWXmKe8oiN6wV4nz5LqwJPwCBiNhXKjKRs/iLZMHYdDaEaDyQD2Blu9yiFHjiTIRSYClryzvvp
AGnIi6ym2T+HR/19hG16k90Sqb+mu96hfBxaCDcYkDywjMmIB9DTBsSwtrUPWLvytpG2Z4llzZCJ
CuACZQkfnv5pH7IzmyjFnxS1cbgViyHPXiYTbqaqrvp0iD8YXxnQzNXciR07n8SW040XNXDh21qn
cMIBjIe8RISenC3JB99EBgWRr/ySrLHK8fBkMPoFNDZiBv3Sr7DIg0OSpe6AlRQ2BpKYTUU+GgYv
517Q/s91nCn2a+LTaRE5JISoXNVED0qABx3F6dTkVHsbH0s4PlYKBWFO0XZhMWg5BVnm2hj11qTp
kHUNT4DowYvjEW5YYItgTuP6lxwEyeMd40Fo2sb2QjADwoQ+q/L3RHHaHNhTL72+LA6whyFTpEVI
ZajDkCOmZwoQzqtvfRoAv9H4/MmWZJghbx421l7Q5gbFe0q4Fsb923LO3FJiscZXHBqAmSqB9E2m
x+9owSkHSrGmlGqGt5P3DDY+6QsNPnIsuku1zbxeIkrI4HU841SGV62tl4nuovuK4IbH08F4lwMc
BPUzcSuD6htjw9Ybs4DYRWBZ8uw3fv244TiIbXjpF7n9/N+vCgDV0MO1HzhuhfmiaIgu8YNFMeF4
/xU13N9Csff97tLKu6V0QkBazZ23ZTgwPmiMUyjEz87CbwTFSpeckFFZGZ0+VSbbeXgYil17Mi6E
JTOiPCkER0/iS5WFFNM1aslQ/l7MGLC7MbJuDp6s0+8P+TRTNzMBKZrpcQ2UKcfr1cuD8/z74UX6
YP91CRwq1tH8zeWtQyKBa+JDhRgPI+npL6XcJM/lzix0Hwo2Ykhy/QATStOCEHOyhpvZke5dXkeC
k6dcKlIPcRajN67E4fel6TjwNrxN+glFc3+QXaKb/GYFlEhN5ldtJnzm24QXj78CrXUXLb4Doxyy
/Qod5e4+s5llZsYTA/XTkDoYoi8It9L+GnnQ9HecLmZjuDZUlqFBUS3aswO6uuewTGrRvVFoHWse
MnUU6aoc2PRcFyLlp8tOM4LHJ+D9yCb6t35hz0PoQ/P4D9V1NJloguAaMoPCMUI5uCuBSYFve31D
2LmYTGl+kSXT4q0uLZ4PizMU1KShstfzS/3N8zQBwWnVd99wzs7b8lNfrB0N4lvZ5vG+ETEnrkHh
ZcX6bvx52Q7etxEbpgtTitHAkom0NbyJc+uB+qRR4trSVSrUfhRkbGVJpJfl8LWljZQxK5NBOpbp
TUjdErv/dm6oolTdQdl9wzwPHMBJCiTd9AwBK/3tndHIqQnQ3/nDfs1D1gqDikUTsGRo5WgUTsQs
3BufibR3g7MYy6GMmgP9+ncMtmTGAYMyu6j3RGK/2PTmJz2UwFiGLdgJbRpLN5XS9d5yWAzzEFfw
nlJFgPkj3Lt4EsV6H5X4mkNl5EwudP3AbquQoCx0kdU5JnKtvEjrB03mbNMYOM97OzZy344v/MHM
WljWFbk0ILtpt81RtEo0gQzf6YEVXqcpoaOwn6lNR1OFQB3iJUiHqfQcjVs52PhwQhcIRPUAU3AJ
d8svNJJQTxKCgLkxrdNrQlgCPJreB4AUisO+TKuT+x0BvorXndU7fbno3dmWaiT8HQ7Q8zz30Zuf
6gIKeBDThzsq+vdGKt9ouES6UQgSYNBW3HgspseufBeC2xfUM3QXKDxt2978eWA0eVrHqiue/bYr
Py+NuNDbzNGZycjP27WDxZKwKo2VHrqowSW3mMOL0+E/yOX8xQXbpCjqx3pNDzIEC8xJJSzIFwa0
ClLZ1d6/ScsNv306KegPl7xX8b/UyzIZMUNG679eF4zn84s5klpTcKIpmKQe29QzNmBSDcvVnu1v
QqReV8io6UfjyS4wnGDwxqpTgxqQcUdue8B9DGeC5OWvtkMBHvi53/RBJnfp/ZpIVTH/zeds/F22
KbnV55BT4l8jwAB6DYfPcy8CZTL4lImyMIfqGkU6UqA1wnYzX4fMl7tiH1ruL/K+U72r1ZBxf3kO
LpR4JjK/8nRWRiuIYUJ6w5G5tss44QIAfu3N1zkxLqhg97lZaHlAjm7s0FrnlgLlMNiP2AIsPUmJ
W9KCe76/QihHOyM8BPEd9rcjN/30ObDoH0X+L9Rx6nPvRrb9MLA6QBEdzDVrfjE6CJz4HpN7mx3Z
w4qVmqvyoeXFC6tmXeQQv9xRTKoybxU63xYxrlvlvg1QPkwmO8syo/bC9rV6LXUW/NTjPTngr3MB
+IlsonyMIMF2esEWrSSqOJQZgr5OYGtR896W0H5gwN2bgqVGrp1MrXxoZ3wtaB97fK6BlsB6oSZO
Q6h9Lm9Qq2pB0PwuPM1OXcyueXS4GrgAE/4Pft3pZm2fwFpUzanxsmO7QeuXIxDTm8w1lq9P1fvV
LQU4MUAM0H56PGG5yoAVXyP94r161ylxxNr+F7+uhMJHlL/7y0JVD5VOGlc1kVei0siMnJi8lXGU
otgya+cpEn3IvFSI/temj+AbIwCbbDcO46qedBXVBzgctxxGGKkMBcKDkGdoTOpVI47P3zGNyGIC
8antSftYZM5yObHR9L6NwXGDIH2aDFzZVWPgqK8CZlMi47WmZZ+I1XbQD7X3fjfudBlnOr7Y1N66
sngZHsmf62l3kRWC/M468/Gey5InYueLUrkoO4aWaQoU/aKF25iwU+OmGRMQC0cjXMwGI1p55jqC
+vLYGst1A0g78m4udZ/pYs/HoCEqRIkR9+3tRbrz4JcqEnYcl+KLt2HmXozaftloT0Kz8DKoudNL
DxsM5u2JM7mjkRqJ6LCHCPsHLCogLQl8pFhrE2hkoxnNePU0txBi5J09VmzX4rBLECYlqnk4ivXh
6yoQAqt/V+zgPb2FaMfn7pYuYFr9X0c0JSQW1XnrBwFlnRDYhpOX2ke5VL6f60z5s2N+QNDFaKnT
Ua1kb9cMbDOZ22YRxP9GAoC7sG0/iVzmbwV8zmdATsDWscXaBR8tNHQJydp1M01eAkIOzMzLsTxx
GKNnOWN/UA5QRpIGhBVqiqCnSG37AHPrFasvw09fB1iPNid283dcMMeKambjPhqfTRzgy0YmGzgF
ZC8YGrNQ9k/AEYZPgPyB3zWz4VvKBYRNAGveDR3mF9AMT0xZ0F6yH12d6JE1J+Tt3qi7GDa656Tr
WmXkkzPv9QxXMBfew/F5PTdt1ottOgjHTHQ4WXTJud1znejZ6fHrBx2p1eHLdPZUmrKWrWAUy7cP
CqQMVCb4N8QZRJTNX2YfVQGlXIM5DSOl4sx4D2sMY3obMA5vT+1L3B6Cg+/SnzGwJwseXYOVkkWd
nTTlIVSLdfQdBhs1KLxvn90MeAYzzRdt2/d47hLl7UWI8/SG2ZiyIFYDl8WdZ9E7mL6cp2qSWgHp
HoqDm89zymAt9W8+c1o/3QNZ5A+NrV/WIZFFnC7jRZ8GnU0B1X4ja9fDlbOOTGJ1L0CttXWubRIz
N/CuJ1I7yFJO6mTybWVawNeYSZRJTjgSw/hvCB0eHrITrH4KfvM65S9HxDhrRuf9Z6XXry2gNL9w
nBiQqxg9UPaMXOG/DUraRCBgEJueFeXhP/HgzkoXeUCLGkkcGHgB+scomI0vp64bA2ZHiTF1yPpH
eXGVchI0bLVQ/Ug9iMBfmOKSQLR8i7JOw8nEY5vn8HMLqsKlR+3bzg5yOMViU/yl4IG4r2r1sgBv
EVTkiZY96+K+Mf445YJAZquIl1qQpbjygYWTuGGfzlFkFhL59E+P4HVHhFck90XaPYDCm1XzN9ag
a5bvgXdsPuEoy6bpNDx92fQr2HLV6QFXq7+vsktfNOTFiJk39IwfcgXIsSHwtaeQZmcnHYRiBZxI
hHwLmBnbTMTCuhsAvi2TSjPaz0v+Vieis/CZVy302i7HW+f8Tx/+NcOk1hLmBLhWZgu9uhmJ+kpi
jD43seVEvswq5So4Kat/i1OrpTQ9mnM8nhvdpxAS/bFb3WKyKdRynFK8q3eizrNmTqMx+CZSC94B
oe1AK32fGmTfIpDZR95z+VYyrYSI8iESxKY3n1ine1SF889Mr4ha+JWCRcP/IOfP9n+pqSq9maQV
RwYZR2fajtIOJM3KSHl9C4+HXcoiszx7b9le5x93PqNwmir/Fd4Koso0C08UPvy149HXr9XSKeCv
cfNhf2yzU3I216cdO1WiG8clOIDDq5X+5sMjXhhsnA/fcNVTYxSGiAKUdIlUwphtxhKpk0AFl4IU
mVNj0wPSGnMLwDYy6AspwQ06pFMmK+5NMrN7SpjDFZBiv0/oMe94P2E6amw/6AuTbZXTLIycM5WG
Wo2hHwcH+2kDRKnsUtJUruwArMHmZs48yhL9zvrF3sjVidFFOJy1vYg56IIMeY4MIIXXY6m59tyu
8X6lm2L21Bf3G4raVhefyMRwnM8wVvUY1/wrtpGhae8+w7aDm9WMRdWIygKxI+c+ISFw/K3Fh2t7
sORKNEfSSm1qua5ym/ZletEg0/m7D06aTJh5R8YNgWYGisMBggopwmVsLf5XC392ylcp5ll+2Vco
ul+BoQYngr0xzLN/iq83D9q7NDxaWG4MIms8iBcBrGxfUA8b0g5i6clRzJ/Zadyi8Qm8oXeqftqt
+lE6vbBnt8nZP4Q8RrkuFSJ9sBH3IVGp5v/6XWDGwIi30piV+4z+C1WrsDgF6flchm5MhI10pJ83
In8NRbbzF/8A0W1TMaWOVN+quOd+XLnSPBgsMYVrUz7LcHeMeOcJmrH/iksKV5lHuac4RH4BV12e
JCt6smJqaffVi+d7i77xU6hMwThF8rFnNLgAu/u1LMkcikMURVPuDa3ejU01o/n1tpe65XfvzGDa
94ModhF1luXnZQUm3EFs0IkSmwKewTrJtE+b9lfeK34XVFgI0iApjDlBhnT+t9wFpNHT3xBTYc6w
roSc87j4WzEyzGUr9/9hjaQ10Q+ziUeCHe0Ww+Ye4yroj42/QNkB1Ssoegra7t+zm9OzOMEoV2qr
uugdyFi4jzZccXA6pCtNocvH3t/ARo+499daUEI4v+rwmo2RmtNGczyHQcvlqqpvXgXCbExG4yWm
a8m91aoK0TYWFIx3fY0zYxbzxrqWfq+TCHTGgRXuEn2E314i1KxgEEeD4PRUrEUFLZg5a501BiO3
xh8HpFaf4fKXg2/Flhs7DY34FtvUOsD0lknfIa7DWpjsoQ+yydKMoF/JfwngQ+NeGp+uM8A7hc9m
WOM8uI2K+X7B1o73ec5V/4r2yLIjll5e49r2LDpqv7Wb995jLEZ9781Vugsk1sLy2r21qtohix87
NQavcUKfH+cH+LXW6Ls9R/lqN0YnIAq1cU1naVyNMCUo6xSYxBK8Zaov5DA0ulh/J+IoE4+MoCxC
2E6Wg9+ImHQNxh2COJJOeQvfhjw9uZPeNrMMIZQ4xRyRAGa25ugKurqt/c3/imAaHoPa/xzyWnB5
gHR0H6K/zl2sDBlxcPVsUiX/EKVNzhlYrtJnLZcbIB//pn6LsTYKFcr0qgCVyVWtr4f7Nm2LgBsp
m1nhkpzcMbErqgKsHYt4SJ+eRyxV3mcWhtf/k1AXTTstmXZRWD80c+FxLY79s/RhRfFFwMYwJS/h
gS7ypM8RnLv8Mx/iXv3/Qo+4SkOvE0pSZ0UHgwQypL9Y5Cbp8BIltgDB9LeGroIe5f/zqo/Eqico
+JsinBM/e2M4dsSV4AWyDunU8iYOVPKrCWnlL7Z3ZKVi25YV7vWYjO48YcgLA9Wms6+AGx1ixmhC
18dx3WWKRq7BKN6quQE2qjD5kS6EuNxFJS4B6IUHLA8adoVeoRfL39woWbQTMzTBP/5hJ0yYeXJl
tZlloXQ9oIUlgd1RSRQs+TQQgusyU/kgnfDxpo5zWbc8Z5CKOQweUo+sj7ee17cDy/objFUXj6eN
2c4UIZYlB4nyn21h4bLAb/Ij34KGx8Yzm4D3pYrFLrtZ4/s6vSdAbKFi/cBVOt+aeZnqc/kjxwiV
Jnerga8oyNYiSXYX92lHYElv8rssjNSIOVd4oxABCvhzGDU7oMcP2wzp+fTqUT/XSUxaAGwP2Z7z
7zaqmQ+QTuXFk036BO45tm+F5vyLMb2Xkn9SuG/9ZtfHX4hCSFbqREL7NWjFaugGdRkWfBAt9bnC
dIC1RU7OA9cquFmxiOLidhPdRHXuAcTNoHLFf+xaeV+dh9/C2z68CLGYMXW3zcli0DMXBX6Ib2ct
sWkuC5Bo00kmUrSx0B8mFFdSsm1FIViE/AiUyf7Xb02Oun5IDr+DUniUh8HsGOWPST5pI17eEdgA
idsajq32+u/sweua1Ixoe1VoFyLsUt0vlF8F5O0u5HW+qqw+wA0K31e2I5xUp5TJviALdneJkYSP
Lc6uP3wRNYpRN9nqhdJzvYGJ7aIQaH1P+/HSEx1SdMSMieJ83lbYpAkkMTBAveB/n3jBYxwtXpIb
uhlqH++4Fc0MuyI36BmAf3+EKP9z1sAO1+IBSbckHUIOy3LzBlhZ9GCcBsjn2+4DUI6T67VkYFgx
FddvomVXyz6RSJv73IgIGYmFcUzC3ZBCMauU1IXt7XsTOcup6EqH/ccsUQLtE5cdIz5UYXMyX4tr
GlzvKRnI4pDXqrX/lV5DoNyVKH1lHAJ4Zynrqzci7CUdZOADAnLztUbCP9J+WxptjUqPq6izE5cl
Mexf5Ee+Z9SuPzbRS6L1SlcNYmDnm8+cTfP/PQGHyLIlsfA6tJOqFXPhbJKHnOopadq/UdzMpcj0
4pd3lKHGfLm+9paOTXdC1r3B71Z5UmgXsO1ERxSFoCJPPhBSCfWi9eE4nV4LO0167QdfTsk/SGww
3nqpF2dny5zKs19VEQyWhN50sA9lFAjO/esAH4qmtZFdlUkRYwl+hqxuAWb6C0EJFHNvo8peAVWX
WB1Z2Dc5IZsLurg2avAVSEgUmm2kuXWCiXJfH1/KCJkMdxnZF1wo5ZS101r2TjklmGgjA0dzHUer
lKpDiFutCJFwWauAp9dEKBmsleuzsVDdAWAue0UnsvOVK4Lj0NIWhetXIVEoCcDFxqmpjI9Cl8Ak
j3Z8XlKj7QWkWMh+heGqnarIDTjjs2PQeKI/CUACV25njCTh18QlvXQ01VdHK4gvREPMeGnhLf5Y
ndJfizVPuZCT8b5oRIhHeIQzIUtyJtuM3qXyqLnecu3fUIIpiffwHc9tAJsghgUeWhqlNk+ZZT6V
dzGn4ZqDZoBJLGlE72jDdXKOSZHJHOsC+ftsXwZFTiVzDRxWfWVqhCLaDkxQbZwgRvRhIbXstPZB
/TlHnx4ZE/ttl/Is4tviY5PXu+SanZovFuHOGEjsPGtOnBMsc5b290QXmds0U1zjAJKqn92N6vSF
pezWOUdtzktI7Htu/4zXvJnvqZkAJV1SVXNAvA0wpOcrXwGSoG/zVUooM6MdF8J60wWVE9DSA7xa
XIl4AlhomFVdBU6iWaDC/A5l05BGFHAvtSkJtdaA9KI+kyHO0ZkzLQEqXs7zFETSBdm4w/WsmXVN
y3gnyXuTVqksc/GTvlzOxJh+0NxM3YViu+01ivwqceuEERzyXl3N74wyAppixJYTzvw6CkxYm+Hn
u5KTYAm710MyFChXgqYqFG4cm3Nf4Dp3rH/1aHCkVzBeZWe+RInx1wfEnAbFyjSjWvfwKnkYrDCT
9KsQP6F9r8TBWXrU/j0cAOzUBL0o9H2kbQZX1AO7O3ofOFrGg5MefeN041pX1ikH/Y+arZ6JQK7I
+6bAlPWIUssFpQHxY6zicSow5cwBYl1PMSM9znhIhRTKBvfF7QkYGClgzbAJI3Sh5T1b6olLlx6V
uHrS3u/NiROdXd5givlVjrG+fGrGQevabPzxYue8ztqynpYqpaRZGc+Thb0PU8nVeqw9BYTNDTlu
vnUyPp9fd0UBtOSy5sokCjgE3wGfK4Zmz/F4IkLM2mol5Ucn8fo/X38La00hDNPeD2HbXIKuvpAe
XwsJ/mrBrauy0eEJiJ13lYufMTpDfTihprsdvobTnPbqRwa2x9Dlrazhm6m7PgqjCTsDhAWGIR2G
490+hQcfpcbiC9HicpMS1FBQWRQce/VCMl2kYPbY74tDPAGEsKsuLNGLBZjYqmwl+Mg77mctzQKB
UlslMm4qkM+S31otN+iDXaaXMu8SmzzfLYg/yLMk+WXfy0dWAm8nWts4y8jb0Q478YoXf3ft7o/p
2ZhNUSyO/Nlc5i2/PAl2S8Am7L3tU9N4Mp2vHkmOJ5HAyOgQSe9LW+5sATDm1vXXyzj3ao9eTQQI
2bEZ7LDGgBNsr/YC6EwachWlpg3vgqAM5B3pwR6xIuWEeQBBy9QQC0tAPkVh436F9iOLFoS2xXpN
30h9acxzJf+C+m42zO9Kw1jlmvSqG5rnBjrWtQEfkZ07TCYxE9zLtL0oGYblsWRb5508kw+VvKKP
089L2oZWTUZznPMyCYBF3SOlr1RMPRFZ10Vu6CsB1xMHfra8DsyDTx86YFgR7JeHyJ/A0wfgkjEx
3VwDciqtFOKDCaMbIQMvpBr/igNvyIP4N3L8sbPu5J/6qiG7YIDEIMHdDoZTU9IZwrOaivkWEY5O
OFLgh3VxakC5JX89OOWd7s5ZJvqviu/GdnnU4hdmQOyy11EXl3liz4vXznr2q8HZyQ3VIikITsZ9
4BTX8ygNlXwRRT9QL8X9KcR63jaDAagHWYk+8ITlnMVdGU+mtDaY22hY+X90xl8Hnu570Ql4ntrM
2LXSqHvvbSLRTnCzok389BoC55zgVvcnunvqlf2bmq0VwWS0WOrkgTtf2zumkHj6idPTQbgcYZHY
Wm2UvKbyy7RASdV4wtJ4kLulJ3NYmYLFh+Hp9z93+Py6V47wxOrYoLKaCxpwPV4dHYM9Ic0B4g0/
lPIPaEKDisusNX+f4eFr/7fOeUlzs0Up5d81N8NthRkT6aiAXlC3vDNSXTX7FsWSJqIAmDx96dqP
QuGjtQT8zFK2EoOwhI26ecFEI3LkLlYNeanEXCaShVHq9PeivndiT90jt/xnvdOJiEGJDbiHQvLe
Qj6zadpe0FC1JzrWDY9lbwsE4rSwD3/uWH36AhTxmYLsJTvj7tdLfkBIXnxOky7kEKOYIDYrseGa
frzEuELlgar/It7jJP/VhqKqFQo2m2x0nU80zo7GafrcMdxWgz15VHiLjf74PcHsg5ACZcMW+ug6
UZ0xBW5IwW0qGZ0vkAbcWeloJs+380+qFGEB3r3pYY/bJuxXhOXR9vLILeS8qrd2N5tXJ5QoWdoo
q0ioG/JAw8jyyS0dr3e8MsaGKAk7DdjaG2wYWrfqPikjIIzXLvdsoSU2apTCRydOHO8x0JaQ/Nqh
S2B7t0sW694KB4NO+SKVOsTJg3yXCIUD7QSHDRHk71nOKoMtNBBZmrVaxxksGtYgO1v2CtyW5wcA
OhZwj7swynHKPoGviTJEsw09dQ6C1niH7+FoZRE5hNXb1UHsEtWNslopuLmzqdgiBMAz2jUDukjQ
VjeqG0r5UNj2cFX815SC3+8wITmY9OiNVxqej9GVTrbAF7m2jhL3CDapIOJersJBtgu5GmI5uR8K
M1D07jLBahZAe0We2kwJi63wOiyfz0noHbKelC0ERlugINFVMRg6Jn1WN/U/hx+3Do4yAhgDr2hM
Z5EA2IHBsUeTzeBO8cmE7mw6r4Jalw1xD5e0rFY8lKGhWWaZLuHz9LjPi0qFnhuC8CQXxnKh1T5m
tviqgBv8MOCqmFNdCPz3gb5Z2yP/crdotHxoGJAN06Vpl5bewcJg4zLK3YYHULxe/FTM3qBDMJjG
jWY96BhudB/7HA7yBxYo8yR9t7bN/ZpjHA0utII7NEnx4OhzkpwEbrkSqEzZQCEVKTYnz2VM2iwq
eIKyckq4fpSpD75FyRli67coeP8b2xCVlz6jn7GwOd966y0R8RXdgIcti/Vf6O1Cc5xuaODy3UHX
MSuambsmKK1nPH7oEPl2eDcF2mgVKuoxuoqg9rqpOpiQtsKAbON/OhZ9IPHJcfEyMPrTblPgFYkp
yDu0zM/sFGMaE57w3VBGKE6d2jbmMJA/h6Ele59SXqRImXFaUehda3lU4fXr7UZXWrk82tSYa71l
1hxpyDNTRVI57/oEreusdNXoWwv2zLQJaDnYCKzIe+oxACuWro1DCEqhM20bGGAZqxqr/9+A/wD7
wSpbh9eMz8glIT9Raz7PUabLC4QgUPN6ASkEQ5DJswfbaO83x28yyw531taYy+mFSQFrWOnASTtq
nxvprq/DcHfq1uCiWOs3WhhA3BONqDDvpDMSFvwyOo/+G2wmhaYJATnqTbgExFiMaOH19BC13nYT
kOWPExHg+F8CJGnkbzn1kwQHxadY0R7Jy/p3vBKTBtrFg06UX8SBV6JziX7ULrV93CaofXGI8uOa
1VbCUFl35nQMZMvAuIvM30lORnOx+h14X6e/sqFExGJdVuF5PwYMaBsb3drrZIBCRW3pF6vI1C8I
RSUk1Co+kW8y421AqjZW18GgwK2bmqeOppUrMZhCjBYaS6BbNKfsnf3E9lJ53xLQ/VgJ/NHPJ9ck
c+27J4GhIuUaKMb7XEnVzWUP2H7QvGrMlqAD8YIG3G/8SOfGG1pzof4h9s7L35hfT/ox3JW/oB/8
JE25wZvzb7AiTt2HFdSjGkbOAQacG8dv9q8cHVPu6VLkVynLTnpAZNW6LbL/ZmjKQA6OAGmdCZdy
jeyIcAqShMjFIRc5YEPhXDroq+K17hvhYAoj+zvGgUreYsN+/uV3lRJLo4W44swy7sf9rvdreQwu
OZ5nzXfWxAT5iM/e04D2syZtN7Dz3gAT7vrJ7892PXHffHjdo2yiJ+7jvEbSg3QrPmuX6fDk/FkE
eq8WcgKg4fh4RErj8/0oaFhsWVA8jA8ZVS8sE17yl+kme2lZnpHTNLGmBaw2CIbjawfWJ9pBQ1Wd
kIXApckDdSUUBYQmLDjn7al4AC2jq89KLOvd2iyj3BCYEM6pzJYguWxbI+gi33Xhy5buCaAzoiD2
7rJQ9EwVEN5gqhczV/aNx7xEvfhaLYBT2l18OWF9sulN2V+3IavQcBPhXETpSVuwvLJjj0GQrMwV
w/ip39+k3TGgTuXPHuafVnrnm0RWL9QntFsiqxAlMVzrNfMarhkQ3hFF1ACbxGJ6QCn+QC/yILhO
Alqt95autt3q7mECNIOu2Bd/zGTRRS8C/HNq9g72zcZMRmf6WT5Q5quxlhUEMr3xwpkV9eIM9m15
jch7fpv20xQSsMRw9b+625dyHkGCY/gnCD32JdT5TI3Lcyxo1tOPMOyd88JWsMh82ldZlAHyYrGv
wb4tdco1s4Xu+oD6ph8RkqLtAuvr5DYvHGFZiXxVBBNRKaXLL9iadQeqoP68bc5hF5vycjkzjGFr
tBXm/ZCUtfpkkYIXnyzby4+xHlUft5sJ28dPO2XzeuOC2pP+IbE6blJCvP79CRpU+uaGzAiDEtbK
dzCeiIouI9NUyKCOzTGx3gDpaYmDTIWv+Y+d530S7TzeXtYCgufuwlnkdIzmTQsXixTI8XniiIL7
CDXEHuB/fRrh0SX+YMP7LHMuIq1L008ZlrbnRyck4lH2Vf0cEhURYGulPAUcvi6sPnV0FwGM19l1
FJvyKBV0aVnrwvNZqqKRJfgY2qnUNiMtCPYwU4qrb9TZSixcQiqElK3cD/8sI6Qz9i3UarlqHhDK
XtsFK+yL88QBNKYNPzrgt7hnUikTxNZdzcm/Ro//Bx0IQaBZ8GdO/rTzHGbUydypLTfFL/IIs5O0
96y1DoYXXX5s3YNwiDArYg1GWgQ4Ua93od8zyTylGD0hxzQaMRtOXRsPs3nVcq4/5xgswJpq68d/
FFyMhoSZ8/uTbb+KDDcbci30o7MZvApk+VMkP1yXjKGlcStyQES+HJkp5BPanNXMOa5mtnPSb60t
iF8v1eMkBPAq9BBIVkfVth4wwH8W8ni06RJ6qIqYcTE24ry4uoKy0xgnhIH6liR8MS4vKZFIaQCI
OiLsbJ0gGpE+esQ2OjQUdJ/RGMTnycZkXZxM8RctE+FOJQRC4KZZAUCvDydxJWT+YuCiQjLayCwH
L3tGVY+UKALSi4kxIVYY8tHuvYkB6G2ygH/GoFHE7J6FoaWw1BQf50fpCJzBgMlTEZyoWseYK1NE
lgOtpLD04G3GZUa01UdOLhj4Zd+6PP5EA0P1cHjUjXfKjzg0TLeLT8e6ETLuOOscSqPeWFM5eshq
/5ONXcCOnx6xOnXfmgMcEDOKQEQQx7CugO/+SE75nYeDBMkf0jjSuTdwg6JMQ2pNCKyIvWElbLrU
oCw83jabTdE+m6MfFpM2598RyPGpzz22GL+Usm2FGYeHHMVaCOfifwILhn2jnkjNlwow7HPq2QO6
nkr/nRJieDLYVCDqP6ugwtVmeh7XuzXHmStaHAzC6MW0KhcpU9/RgosZ7egupxNM8q//BsfeFR8s
vg/jZCzHs3fuQEkCm9Hu5TCW8wa0G+WQTEeQVwTK81+Jw+rij/b5xUYEVT3qcAKPRVop8cWd2uAs
+IxL1kdgeyoyHRLr5X2MetHWXOMlGt+uJdCtfSd2jfue+8WJNbkyJm/3/KX5/2MrMIktblu6JX4T
47ag4pyS2WD5TFjVQcf/fyqMEYqhc9q05VK25GTHZapQAa8G5SvQYoZjOnjm0vV5a4ItlJ/YWrQp
4qo/JcnWGtRGDMpBhBMQEfuDARdxxLHXTHJZ7S0Vfy632sF7/JBJx6oBxpobMGlJeolj0S0Uo+w6
HZ+bnc3Z/hhSOFwt2Rk4GObIjq80oxWf7Ha2cndZ8OCGuN2wl2QXlq6rwRLI2CuMD459zDHQdr8P
48HX8zZtrc5XC9bt8I/9NpfM2f/5XxBEduqHjJaGBXlc8NdElKY5ygvjup2yOk1MP3XVLQNMjBBa
KKwj0QEwmSZVnJxAYHx+skDnw9fZU6Man58Q5gmHq4SbbdPLx6H22aJ9w/MEP/1k/jFuqxtbaN6q
Csw5IQTimRmHVyRRUYyFApAzyHZqyr5RrW1IWmpqeUJHkjPXXM87+yxtBHwe2HkWyJf+DFCSgHhI
ay1vHnC2TK71xyXJKJpSr0sluVY1wnu/H1CiRokosT++XoLSTOEf+wkyqNJn0t1xqKdbhLoqsv/w
ykbnJRkMgpqnSK9Z7uPHPKwEOgxOXGtRmU6NKAgvya7ADoy40yrRqzqUYUPhImfo4UFi3jmYTXeI
vD/JtlEiwNcbCRJ7cBzAQnM+SaOT0FONqUbaV0kPXLv9PZCkOTfmFcnuLKUF8JaY/H3bEBr3+gtq
BtsrjtjSR/ucO/6Nageljt1gL/7HGxVES4WcfjCH2bN6vtp4zQwoTewUy/0F9YiNEbOksn2iLrqg
wOfpjw85WuEX1AwvV15KN2Q53U3uCbV5X5cKWVXmTvAHIuQPxhismJWh6qBF2dJKQHbh/dcEQ5Ck
PykiNLSV3kCe/Tq8HUDncsVDITBx9NeBhHOXdSojwczZBqIVQT42Z1eU8u1x3GLD8V1eYjTejtaf
EHzys41PqsUYUYUQU9fRrNgGth/m2gN4ejcvrUvSDxqW6Vd7JSY2mJxapZ/iFbj5h6WocZFGkava
vNyGSbPWndRSfR5kvWkGH8aA6qKxjL7Sqtbh9gmeY4q9H41ZW9YCaTyAHIGMsrlHz/tn+/W4PG4Q
MUKVnZU8+spBQNdB61UJFYNZHvavKAaS+RmAm9zn/Wl4C7+uaFHx9/R5HaeIj9T1RjYBQzpHkmBm
bdafeW//2PBQb+UwLY6EaGuPBVxV1QqOKX062mYaOrnZq5qh/DBc9h0GIHhWBDpRbJLtsrv0CqDt
+OKaotXYMvFjSPp8+z6+Ku7OTZrvQk/KMt4fFMlsMgoS8bfGkfG0d7OBFkw9q0YxBGBtPd1NYllQ
WrWdIjRHQEOsXKu8YOBhdNSgaV63gStIBwOPeA/lcKzZ+iuwOJpWznlpqIT1qgmD1xTeHD5JgAXe
BKjGMjWeNWwVdPdALGxs2h9wH8TlhN+6VoG4RZ03oxpF9oKbOS4N3nc9xbiaP40u/aeaPgtzVLRH
QLs83C424TfRT+AInmABSqhxlfzDGa1KclzoMCCITFFyqDQCKMOr60dzlwr1xjoqomI/bSkZn/Wf
X3n5YiogoKsqDn1BSrMDPRNWCXosnLrZxLyUDeEfmrdUHyST0BMG+N17XqQAMuLOSHWFCOJzoQv2
GrXx85r/i1vAMgobCm1ANjLdqbWphZcIgCezdtDgVaVcYZ0sE5ixL/EMkO17sSfTwn4JvGsLZ9wu
8LN0Ikj8tOAALo7IXmYPs6SsAwXBqeWHPlaxvG6yGqmdT9PeaTRe7hGnmhO1aNKadFfKzbKuzyb7
DmF623Czzgw4S9cf65LGPzMyTaj1exUSU4De75V6pSRSTjpSoF6Givs11p7wc5DML/w7VCH+w9LI
7AlKF24EJNF61T7Gc5zl9+SM19AK4xb4XpZAZgoGt6wNm5zzX8aFfVp40FRuxBVtC4pF66I11TXB
5MUsDhCD7jJO0EBMC1u/HWj2Cvv1Nx5nDtEhkMLKJF6ecKXbUwsAi4w2yEkf5eTP/KLVfPhc22Gx
XlC2jSX4nILZpXiMzI/0kImckLX6jmjCnVS/WwK1XJL4IeoDdR7lMVDZNAqlsXEryOipDqnRv8oJ
ftHO+YFGq+h5f8knD01SoaS/JX16ukuauDsWBpaG64QjGb4Y/jABTjJ1jNvQtylokOKxVdbF6FT8
M2F1/uu2b93UnQyPJlN2lJoX0m2QQEVcUgheE2yULIK4v97LD9o9iGfef4h9eETcKxloWmmCIAVB
lQzLyHsqP+TU6ugohKUm4cDLl5XXE6g3eypG5w/QixvtvfuVK5ulz95YW/3Q6nwfr6Y6vX1jsRBh
Vg689A8q614K/uqUZbUA9v0hy3Knn/WcyCXHHXYESfxrFW2XKjxYC50OfChEQDrXLEGPhJ2TPXG/
+IrtXst3hZE2yFVDU0MZJTqA7Mwq0M0VMx4yIVYTiwT/OgRtrJFKweSJ2XBFhoZZ82Do5hknTFlP
YJVbufwXRuv9Mokm/MnWL/vwePl0vkSticUg+pJGOQzrJOMWbyMMNnxSEBYIELUoXL3oeMpTLUIs
BblSbTAZBOZCYSZr/XKFkEGVsUBN2jPppV5GxHwkWgAmMJhsa6LO6QHAciMwTJ5R9NZ9RJahMCps
gpzl3/vAABMO4yyqGMqQSqqnaFBfZAHJbGqVSaYdM21ra/+q6R8YJvsGIAi37CTclfV6Eu6OlMFu
jytstM3DNT9n7DNEMPTLRdp0OYedTD2Q1PnZWapLc9tdMBWcMtr/wbaRCG3CkbMBGFuTaNs7MPfl
BvdxZJCNil8X8fMkOJOCZPBdG84oytGIFhvW6YHQ/aHuvLS1wEAPVIMyNdi6M+R8tT0JAYkfbIhH
KtjO/0eNDX0AlxB0NI3+qmf3VLQ5Y1qvf4QcRXDj9Pbx7FtXoUl+vDh5oW7K5qFl9ol7K7Xubq7i
fNQWSOSXzmFlwum5QFyd/pnptxP0J/Bj/O7bzwtV/+sN0h6xqh5aaCW6mu6L8nVWgdrn6g1OTkpi
BhMpuKezr2jgAPZlTRnIKWP9/uqlIK3Sdqx251r3o3H11fSpSE1tq6RJoNfjoIqV0kRr/+toHYeC
ZFYG3XfoY3GryR3jsKGYscuvgaeLYUjtUbo3c3zSLCTTwzDIRNX/Vg1yHr76ETNK1Ynn1pVY3Gox
4jdxWaJrWMZlVYiu/x919o0AcxMrUwFHy9do5PiZw9JtElUYthB5jxO6kg/WktqLpY4OotIGVhya
XdF7LTt42efNXotoN5ZLUg7FBonUMaGe5mg/Kd3k+1dl3XWsa6INL/T+P1lEjTUK2rZMfxRhYlqM
oFt6UjiAIdAiqeOdOQ8UD9yAywVatvRvn0cyXV1yllhIsJ3ujWvHfOimiZ0krqE8oO+r0vSbziyY
dK0Z8jtEee2iOb3lmei4wv4yP4BoZmhAMCVI4UNkGHF+kXgemoZIG/XQ2SsJleZ9RHOPrVoDajTb
V/lz4NJaK/JqPJiOe4HefK+adVNReFXihiepTKO14dgAhbRC8WnELdXy48Uc25fq4tc4/4pdp4pT
IR++6mWqhRoh8jR45f/00WYtJC1wHkVaWBnIkESoXdyfGNhBW1wHInK5Ul4P0tXpCZ44FGOu0lIG
JgDIbqWDlZKs7ff9HTyGsS7PRzxL8hhwWf/syZraX+vGmN/GmJ4em8bht6D8oaippRw7g8FdCcTz
0i0HKfu59SgOSiu28ZlIfXRpqudEiJ6w/jeqwFGz+zTLEFKmmCI3iktODub7TI3QY7kn0R8ISm3I
B2flNR1SDb37S5RSH04imgYPz/lN6eb8cNReiNfJx4/IvZfd7sxazu63kKfYMCGXgc5JpaZ59a6t
2nWumUn9+JWg8qpG9UB/kqJ95uNJwUdKrnBunSDHGoD9XY2bBl4Bxda45qMdbPf5uEdfiANQwSIw
isEhKbk9SIO6nGWm2iJMzPJ07zdfrc9m7qL/q2pqoLn2osGxhXD5mHzk9Az3Zo/joZN7end9DB7m
kUtVZXjlVzt50e5cGlKu86celB8ufYQ3XNimJahAYj90mI9ovGnU+6s1a2luW2upvd3Im4W5MIbP
ZbL5sgCntwrn6parY1KzIFBrWfBz0EsQeMtu9WBwdRNF2CBAX9m7FW5rkgaYb19nQFbrN15fxfAo
vWm0k5Uf9XwmVMxLsXNvAIWFxzkJfltspuW8xrpGliBMXES0eCB5fsC0qfX+YbTuC0D0tC7SW5Mk
fBwcFTfsbKLYqtiFWrt35SHauwe82yMiddnAe1Lb71a0iGN6v5BVZheP26W3PreKK0/0V0rEtn1p
TCjBKaFMhexnapdfdTJhMr10eVuHbMBlnpjjlLXEkDIL7OuAn4H1rDdB+zOPr66slgx+fuFrqWUu
gBbWCC2jJ7VD8kvTbAi4VIdLQvjGg6nF7FXRVMGEFk2k0UBDvhssowkJau7cSinu90zH3nU8Xnbv
zjqKdiEpby0sWIM5wtzTyXnp51TjQMSi/GevhBbd0TJlG0AFfqYX2+QvceednQpD1t0uWAef+T4g
KC2wY3KtO0ARK9mEpdlBK4Bgwn7hcqcrNK749wiXiBTO3v2sp8yvOxV6GYtO2kXoP7g2rEwKWp0k
nouAKWrz3xw1hEWsMeu9pvyB8/WlnDoh9Eeyj4ha2Y8j1o2KVgA+Fxp8uxrFg1nAZ2XoMZCmnEA8
6LNGlJ+JGtNUtTWAMvxhS5coWV2CHkMo6xpAiZ+V56xPqAuYSXlkjdniegLkJofvqWe9cse2dwR1
6x/Lu7rc2pdn/bkcihCT+ZbBkV+FubSgkdbRuyhpU0c+l7Nid8VILsf2IN5k+Zo+ac26l3iF06GD
VOXx63EdIYKsxymyABQ+qItIAXCIz+NiT8RMrFpUFwj3eq60JWZTyOzXX47Tw8yGPX4t9rJkFfIe
VAYvvL6t8CRcgi6ghSSjasK/yc/tUai50G4FbCAvsFlGu14cNTL2dTwEDubOPgzGwq1jJA+mic3L
Wkt6MHJnqqv9E78GBtXw6d+smie4Ob6up94yZEd42azNn2kvDQP8PG8k5dPdmDWBsfVQXgVsKDCs
3u9yLo1KHH51M1pfHGl7vqsP1HRZN9BC5uHrlUdkTE54TOVKX72ssPmPkhqFriACvSkJX4hTrfo5
yORjj0lLfzRf4+RfhndUheVSOaZcN2X+W0xNsoezn2fo1SYyGcPiAvOIq989pod6pDhsPmymO1M8
XZOyeSbhG26eMfUaJchofILH6UTKnMq0S6PapxDciGZyGEVITakb9X9tzwazd7fRRVROivRIS2x4
CncON6QjLogkjrtNngH8UI49+S4HFrHPh03ixmUZqywmHlgJ11N4+mGzPyLv1N7g0qd2RrxB99Uf
hr/wNkZqq0CCDqeoEP5nhmvhD58BEgevs2voRlmNvkxouRGaJ6GnkyHdrW3nS93tLRzuwMI50jyX
4Ms0HzB+3mGsAjgWy43aakmedmj3/2DsR4EQRPwmzv2LtE+QOSIlhuIjgZOiJzwf/saYoacyvbIS
wFvwfRfKZMYruOoTK3dEVHprGhpzO5SFZ+ykIM59nO9sCu6nDTD+uYA6F0gqWVn1OAIwKawBO6Cy
3KRTlLot081ocQ5Am7J6mszcrVcX3FnSzJWjjIjYsfwurjAE7KwohGf74Xnqm7MNryJjK0n2BRHu
9lfaAMiqHQQPbfPSKmD2ny3aJicBdPA5jXyfdqyZVfvvkuTG4s2SbRQGsfNkb6ZwwMVgnKducHws
ZtvTKtFDZGKKBJrRupLd64TW5Ew3+JbdO51of0pm9itGCLVBuFM4Qhgy/d45d33Qh2dRzd9/TowH
hoWpP9Xn4zN1NKhf+TnUeKZ5x1udMmayFxa72FFD1xeHlu4lzHj5qmnT/Y+UhcG5SM53vUHCgCdq
OiQ2fXK15ThhWe5ueYKzP9Om0eLaM4KSHYs3vRXIePCSF43VnocBsLgy39sR19D9+O9wOXPiJqjT
7zDU69o6eB/aPUVPKvxGZl3cvmz1SiE5n7MJhJMvDXfaWFc8yVSmLMuFjO3bFmkhDU/vOEijvf1A
J6bwt/jjrvSLLGpkhIRBNfI0ASBr0Z/ikw54tJP+n72kX2psJ+GOWrW84jnlASTFeaXUzg1DH0D9
lYuMSctqgUzFSpSUnckFhZOfK5A78z1sFsXFb7SXzi19SDYgUnrop6CAKweyED3JH/ZixJaJUTxc
M4wb2RlStICKP4FV7Ecx4HtkAPtSrjDfWG+Br6Jz1E4ZND6FBzuaU7FFFXB3tEsIeugk5tvbRYg0
HHRQ6cia6eH4JC/O7B5WipEU4ALd1EreYra92DlunfR3z/A3oz0N08eLeHUbpiJeXe4RMYGkutai
4QgFsxyU7GeI6wSFsSO6P3FX6mzkgXeeus0Dy9UGM1S+ryZrVCg7UGE+8aKO7xDAQwjEn/NdMgIY
00fgLwwR8NZCIbnG2LPTC+3CVBS1L//gYH7Qp6Hk+8WIFfDhdhdfu+u2yZszbCGl6ToTSlza5I8T
3xKSId7ALBALT0uQG4VpjulmpPyUln8xebE4FPmsRfx4eto2W0Jdc91xVPiQAN7V/2LaEtCrwZdl
TiQ+VnS+xHC9Pr3tnMyX1PLCkmB0lV6H0lYMfSZY4uwiZJEc4Ej1e1V0pqBuiiyFZlOze7kaZVXf
GR0DHS6pM8jxliqg5Va0ofni3y0uybLaU8pAD+4p+o5A5JL7pdsQxo75GeaLGlj/rrF79cGetawr
B4Khowwr7xcGcNsCXahnqX//G8daDmMlhJp6zbxRq5b+6F9jobKjoyfw4nmWEjUV/nn9DQbWtsj3
a5cQGSrIjgL2YJyL9XAZyG1xd9G8lMfUm9+xA7OQRXO/vXljBQVn+tLSSDQw/C07N01EN+1mjHCs
BKlP4w20uqfIy9yxCzcmR24sVj1/146wkG5ngqzsyPIpmtdvO0s9+qxqCgThr352jI34CmZUyizL
pvsvXqqAvg8wg1H3r2w5mnAmC+P3llDI/GEjPl4EM4qDxU20FtlagrinbsCfMGjxZ5ikoXiQnDf/
3bgiJKMCCggf72uegap9zcC1uH58eN0mKNTGWXXEDn70+vqSYmBT/9zC0MofvIpcq23OVslsUDEB
LjGWDQTEfGg/fKFK28zEOr4Ti4UvSJrXc6SjDBxQ2d/Wd4Ee6X7hnGNueBm5i0yp1/kih733w44t
XBrTm8ReUll0meLnIZIBvHMmU+ydLwoG6BwcIy1OEJoQ2mJACeG2sDw8bXjK9g3o5zxtLP4td/wA
evQnrVreN19EmLW8xw0QhUfWRPvlZ4sgGRIICCgihNiTAHzJF+m8XISYX2JZmKR8T174/pLqc5o3
Sqbs/HYPbKEo2HyP+sVqP4cT83I/2dZL3AP5s2zAo0z9p08GmyzDUhIBff93WqKTZ792NSohV7Sa
ZHcSXoZYLlLJIM7Kg864v6+z2BuR1dLBW//u3JaYPPlGIboSImOQJcVih1q9i1YLJ5eIs6l45102
3rywA3OZ5tgGUSRnsEkEpmHhyNmPgiEHq32DbSiWeujmICGAXDHvAg87wnmx/ta26JFXyZUY4lhz
hfSIuZCy/qGpa4przmONyJOmeo4CzqiZTOIiwUN1MyyEKNaiG77I6OtKhaFq3RAu6mlHVVpe6lO0
KfwpjPwbFp6Ks0nO54odMZ76ii1d1Xs184cKM1xLGgCzAGbA7cz5C/QGbJ9uDm9Q5WhgRnQjuYsZ
ogX7aQ4Gizrl6ZOFmnhm001D9QCNnpFdZ7Mampozei6yUxfWjVmfjHYomsuuF3I/Hw8f+KOvJaJm
4cw6NRXcXUmC37VThryomW9KrpYEzM1DKQYVN/dTfcIa/PLk55DNri4i6n8ctiPvVJ+C3xwbdNyA
OLQjgEuWAoc6xCTkmyiTKusogj5x67rvGvm79miyd0Mfm3qHhoO8jNTJW+DpHiL0e3wSSgLEumHO
W7MCWhA16QGsk0jsqTkNaPMPEIV3wJDJUz98pjlS60sK/Td3ZRqfNIjufLt33TH2Lx9R4oAvvr38
r5KFta1qRO+8sewCKKdmOQCLtLm8gzgP7a/vR+oV/fvUL2sYzjhOqFkFHU+Vzf/GVib34EhcXpAa
+uGum2EsUGeZNlmOvG8isaqL1QQzfnrzF60tQlRhwoVYZyZcGcEXWgewdPzoTQJkDCmoz3y7e3kv
ht3BmiXbuKIdQOs7uilCbvd0PZkyRapon6z3kra+hwhmw5mFDF9TfHYg0T9nmnd8T1Q8P2WE4kMI
nonL4y/IsaFYMrclw8jKXmyVijA7SePAX+NqLuZmP6+5cOivebjKJEmILvgXsfhYBU7Z1OoH4eoy
IZZ9k5wGbMcD8j9ERVZOeI/C2tuAD8D6tDWONxzfhCzbubYCg41Fy0CXDB+/jzECqo5H2CSRMu+l
YPPdt4rjOq9SUae4xQ/lBKOm56xkha8ikg8fxF5qw0XZoX2DFH51QbgLA0cXph0c5B6YvWTHdbMw
56V4panQyLUWl+V6/pf19arMdom2KRCKibIZXMTdSCWJAEq0TVzUVp6sak2Mko1QYU4aFng1VWnn
DfHJkfp8apvwEoJ2DFN0dba3GBvdpY6oxZxd6kWfOa9Kqorr+Gat47fnE6sdJawqghvkyKrx+2pf
ghhPoxt7bFrQ15HR5tXBxOpmInw7S0eOMA2yI1ZgZ50jXHXxY/uTKBIjUNc2MBW+TNj+uqdZEC0h
DH626YUCFw3eWsDbpme4ilnR3G0aM980oNOaRL+DJOvTozM997pp9x8H1PkK2ga9ae12ewMskKYa
ZikmpnveWygpHTV2qxg+BPwgyyuSEX5PAK2Ao0TzOI3AErWmXHU3IuzwvOmkpAKiE1t1oY6wXX0f
GwgKBpt0EI4zOO3tcnDEOwUpF+0aP5T8eZu5wytbsIaV3nj0A9RSyKjxUJJf9erSGXkiFks3s4HP
P/Wo+4vGXXulINl6y5s0gmci4FN4nnFlznbEdEzB9k9GjYfdwCpXqER4Qy+Yytd7SNv16duIdisx
AV/cB5lbZrz57vUezsIz9p8Ma2NFn0BHVYC002nvyEjjUEvZv6/Zg2YB3vKF32BFAMTKsg+Nx+Pz
aFnSEzGLoRTc81TOJ+Kj/duMQexqZVyWX+3rFuF9h0ttllSghlEI3guavLm3XY9gpCAeajMiyRUh
xsf4WT0Vhx8va1/KzNWdq8dNcw3vqCXCj5km2REFkdcoGf57ccv2nXdd0PKa+bIhZpknEQHYZXxY
HAeG+F439QFkDrGfsRL3ndDbp2wOA+ipiyscaBgKwlPPIbtC8rQXQ/GPYnt0K8YsGFhvCpZ8tSIA
6Hz9OD/RdS+tgpVSNzkibPqOC2qGlJaC0fYconvx7fV2vHkQT08LAdZ/l6r31NChVO5w6ffyPm9k
/OveeylaVIwUtX/TfeoK1RP2p3/voUgiWKnjLtoZL9kiGpaKmTnUzYrB9SEGBbkQ/7QO+j5DVXhI
Zf/Bv6Ia8FemNeqVPtFfZgEvYFAo5f7fAw7hCeLe9aFoyQoemOfccdvExUm/OVSitNv/WpLADoxC
IfaDru2JSH2RGio7RQPGs4rQTmxE4hIawskmWL5NfBhwY4YqEsteLZiumXb62fxs6T6wMpxLlfIa
zmzSleiPdiXhUzg7bD8nXThlKtUTJlcFU1eDRUM6uPRMzyH4CAMlDGhZXhw4n3z8cK7+U3pcpudp
dkTv1FaxR+fTjHX2yPfzYgG8dDjYMAxiscmYkcuWn5cvZyswofyHhGp7ZWHyieKOBr7T0M+lDs2U
p78DGF16qqoJfPOd7S5T9V7504a8+0vtZm0lZNwZuZ87YhvbTfGMPr9WZfvozsrxU7nYseLFDqC5
4ZsivEWxEOPDhspaQ1aJNhvNTyzekX5AAdsbkxneZCoDc1hnY9DdOAmXzGa9HcC5QWAWPXd9h74y
rlYAT8mzRU0k0fCyw68xQYbShh9dmXQ1Lfvcmu8Xq+lqC+IPT6aHoHMHYkQN1il9i62fhXhMmkH5
MasEKE9CbtzKdjefwSyamdmBgnIdiUrwzbMFgIetUfa9jbk9eK08ayGF1ze+BrDRtCTwcdpjQXM+
WY4GXZOBCz4G3XNz/itYERmCCM8iEqxrGOlZZKAl3oeySgpC7KIZl50jUIPa6IxdKyaiTmq1fj+1
BCsY1l55DRoVxuY0zg8rG27uag5LteEO7RxA/Q/nFx79Bh079QKUt/feAwmFIaPeezAvplueo/9n
MsQSR+EDYpmqEUs0pe2pWoPm0NYvtF0bY6NByvi4ymeMQE2bJ6ht+oUtpigsAL98p7c4vU8azddv
Ce9z7QLRBlNa5SOoA+77ZvTg5XuZQc4qzSsbQmKy4WLGudMNsFLwVxhG7fs7WheeK92fxVJ1Vlo5
NJXqAhMQA0AYpCcsXYrec2F/wFrFB9lgarF4k/fUjMK26LaVSd+8WssiazhNBKU8Q83xgORE8K8I
7/QWybU5Mg6Hd8VHVedehC3ImRhc8sLsvpv8dZBXfmwlDZgKnzIV9JO5gO5854uUagj6x942WnXX
qhjk97O135+OYmaO9cy2p4mvzL3gacEyDvh8crydYHtsqIJvnNZXS02bvHn+49sEJ6B1xPWB94Vu
qQDY9iQoYOJsOViKu1o7NxOmjcPFwsxo3V50vx3Lxzl/wghJWiyBaDl0mjbihB6uGN8z/LK8qYfy
cJohLqSGn/q1eJmbNwL/+K+GHgzlJRKdAFDnjHIDOWhlYyhfYzDOT4zu+F+AqZZ+pypg4YqG087m
/gblBV2TTjNp9GxqLIfuOJJvW6JJG0NqIGdYQzgtEA9u34VfITy+Hkq24i7sW9i9GNOwXkItDOph
XTPxrTx7lf9o382mYhSsd+InV5ndX9UnTpfxpn0OQgZLiAHIiiKkypLkAykj0btNE/cSurjR3Stp
stpX7vqBprpflSGTqls1DsYjy1h4pVfRSiq2SmItg2UEyh/w+/Egu1YoRiYy0HdwleOjmWPcK+3C
bwI9dpRXV7qamT/l+dJMoyJrIlEezFHloun9VCMas2F85+wr90PZx58li9mP28xT2YIVsIy8L2rW
Yrp1Tv2K/VioGpZAxpOE0tJEAmhKth54+7SQcixQezMnbgfx0c/aK5LgWiUfv0L7Igg8pBkH6N7w
JTa5mYJOq5CP3O6EWEtVFbakYTBf1SLqc1USeK01c6OMbFwzwaRdNznvOQtflLykWj0/FPJtr5qw
ivxq6gibezBExkL0fhV2k4SsWUAphohd02KvYNS1OhNbu8RrM3/hHp+2Rr7pGeIAZmUMF7W/7cXF
mRJZafCXtCLWTaoBLMly26wZRLDWV8B+zD1v3fWG7No3DgApl6a1NTOcS2O7KVFi1BdD71v2NRlQ
EW0HVt3fKuYHdHul6QLYXQkT4MMoQvciFP7Gcv+nTF5SS5MCWZZ1+RE2ToL3JuPlEd5BvYX2e3jm
NfbaSY38MkOi5CL92ks6xNEZ91XzypPO4kWArfvrJcKJdIpTs4uDhDcGtmTOJYhOIYVV0R2erMJ0
tcwNl+/WnyN3OZ1Mos5B7SIIQi4qzT+8WdiL9gEzoSB9OqDWe2KSHyilBR5Zv80JXa9jWL3jbuwv
AZ7s0w1bxbobTrlb5rhjQnyJtEujObgUrkim7/QnazA1ZZ1osnJ5dcLcIRm63kEJV2U/GeP21fDC
gGUYLbgn69Ot6bChQuRbnyH7eIyBAHot29Q3kVMZ77wwnUomDKDypXgnYeq/KcQaJjgMcod8A0uV
K3SpfLCvezj90IKS9BnJYn4yajdlMOxQUeh7Xuf1oOjpNh4mDGxuVk84CRabsvwhoePHGlWsz9nf
Z6vEmVhaH3XwNYNPmUsoK81iik1YxdSTmItVTbGzVRCmJrwJgNT8/hXP6s9qoQ/KDXRvwB/786Jd
FNfNsZtZQLobjnn7GxP5f36pZ9se2/tJNcg8ycAvlPDEZFA2UGL9dZwKMw+nguE0oEMKhkWWPAn1
0oifqJhw/jyNKy/FWgZZNarGDxfNkjGSsHeYltILvaAZ/9WMQCVYlhnkvXGHdKQIUrGdi5JEUKXY
2vmMA1BE7OqzjmuAKT91NmQHmz85gmHXNGIH9xZZL45/jPgRVs+gEaCNbyv+PNPCwoBfB79FePHn
4gUfzmtvBmcoMcAJRygRWRHMZrAnrsDdg2zg5AxO2LyiqvJ+IfEh9jOoKxYPw72x0lee6s0ggM1p
opdkOWgzLGsGWYUDeSa8Vf/zdsp5XeDt/+fu6TAWLS9mkkQpgn+mN2tksrDRfhC1TB6a38/smXJl
E7ie8UC3Xmm5WK7Wkd9NasjnQDhuVgXEVUvFEUGdtUEJwWHsRqgWfLaplj5ULxzpjS5crDfl5moV
4Wf+lRZlE4Zq7A3RmC5Wgaef1DE9++1tYg9ahyMwbYiSJ6fI+oexyeZAyumYt5ymMtPf9kwTZMPp
XWiKeoxX3/Ybdn8kAX/WmXsNi+va8ZdGwsofG/ShRHQ4DkjWX+/zmTV8WCPz6Vktg4IivQ0lGJ/l
bxI9z7UTdt/iUQoiiyncxwrnwsCtmi5OYS3oyI0B8F91fL5zg7Pfz4xREwhtv6g+OPT7mH7k28dC
M6ym0vKaPqE01v5/u3jBbsSkVQpt+eQvYTF5gah19lYDq5/ukQssYxexDIi/tHxXhcvMUzPpj1HM
/ZtmudRmj3OkQhffuHaOXhSHWqPMgyrwLdjMaAJASdi+P16K0rd5ZFcYvvy48yvgYA1Km75gfRJH
haa69tzpE8QUkZq5gdbCRDfN8ejTGM3/1XE6/DVDHIF7Yi4ZQr6KxeWB0zTO3SRQA5qjAA7Tmjip
+rcO84TEcx2kz+tRhj+ORKEWT4IdmuGYNrsaonhEchdr0HmqLcOfahSK11Y2gF49HVZFfqMlqhZm
H9hlGINHkkazrSGPj1zQ8bUGVglhRoq2/cBNOZw+QSLaE0hD6PJT8qPq958uJu8Dvke5ERu4cuR8
dh/0kK09LVAPeHDZ95dTDpLLWIxw9FnUDaoJ8aMcGZ+SqKMKggbWEdNfNeLbu//fCoiR17RnSmAO
eGvPp2FKa308tjYd4wIZ3NxHhXRbOH3rFkoEuDFUDdO2CyvQMT0phAVus81+n34YCjFjo2NZvd69
8tvbu/y6GV5Qrd+qezP2gBQMLgwvOEOGq6clR4eZzo/xpdlxDsb38ASVbSHJnKaKOWxdj1pHPbHi
L8PhjuWQbI4hRhNmPS5u1HAUvMHOvOUwYXTJ0QhqRv2Xejdy2k/tXBbdI97+P8TKHNo4AsSdLvKC
u3E8uth5/Ko5kypKmuhwr+bDqc+js5mWk4A2rJRZSyc00EQdO4Ct0Cy93xPHsSf55gA08awRTnh8
4RfesP2tG8LFM1KNy4oAttwiu6QRuBlCnPYcPpxjnXNvHOpoYz7B+VUOTAi2uBTq/vIs8oXrTKaK
cX9MYOx3DSGiZK/CCyHoMevndapwYU+UAnHFmLOq8ARSfr+b8WDeF8dMyzBBAHA4Qy8DVZJ1lIV9
lSWqH9m8+zXriDBah6rsLsyFypTiMDxucALbZpupH55mszLI48KouzaeXHcgDVkp8YhMan3MD4tC
niLT0NImuKyLOyw6CENEi8lO9OFXp9kLgeE0SxqCq0/rKDlvJ0LYhHh6p0IF0rArm2Zm0+gNfyhv
I81NTKW79SrGE0bUszKNn6ODNcLAZVHWgkp7yCKQE/K41BxnAtdVnSrqImlH5nI7ONHzAWtrfHZs
tsYM0FVteNHkoYXnjoZ0HKyEt8iL4KN7fmNbpyiux4qrAOil3mPeStFGnnO3uj+PHsRovRn5OZQI
BHxtvcWje6DGA0UX9spAcAhnzLxXTj9QiBWq4Nefg9SP8k0YcpPUdMxROZFj3JloNPmAVmjgYrSO
C+iFOBTsfvd60iXCQxsd4nyQlgn2rZQCwzoh67AIL8OjK8yiShV1fSSFvqgT6Jv+VJuIDCWxkZAd
sVJaPXhzmDcZ2WOJmescUtobLlGbd4xA7a4cikpnrEiktzYvUpdYHtSUUOVA0n8YKUSn7CIJgK+y
cki8+OXSeWZYc5WDJ00ykRfJbYEFdHAD2WS3epQSkurS6LaZ1sfdoH4iXIfuWvXwdk4p8rsGv8QU
+HUvo4Q9/jlq19eZpCM9dbx9ZZtYh+J/IC+6ZIv6xPw+7bI73dXyT+Tb3HQYn2yuYIjI/nqxIwGY
9X1MnOWOWHmQ8o5SgP9wWvMfTk4Zs1KpB6mnPVSAhXnlLNdH/ss9r/6EtC1ViC+UEHE+oI+zfLmA
HMJpIqDsu1J4TNxYxwjaikRW4fUOjUB99CFCm2go6q0wfoXNqln4m2ks0kdtVBnyzdAUi1qoDv/V
lEZBNYPFLYGFfrEO1Dtq6D/55ndcxZTYp5k19gVABiPGWQhprLMnTCsSJmFSkYyfGSfUEnrYasKI
FxKGPTi2bndRUYQJ5EPsaWy6RpMZWhbebWLsAsTDCIx/wOxcBViQX2NOFkus85SaLnLGY8Wj7izE
SwwGGUbesvODW/BcB1WA4J3thvfO/SMgheYV5Mj+ESSZUONomQ4nXj7uL5MCFCA5l4jRm1+3fvVt
kHH6hM/S1zQoJrk7owgsT5XewRheVyFGSYY794UovUjMo7D3Wf2p+L/FDBJJLpLjYxq4rttviubo
ihHXk5LiHa1zO4jHUj9P7PAefrjfHusBkYvaOTwVGT1TX+WOPvyhr3usNIfIQBvasQp+BrYiE3X5
uHXvVrTZzUNErz/5rpOG97TAfHiKUQkwJq2WEniRLM73vu6R7OgOi/tW6nIoxXTKI0toRttpZ4IT
XKW9NjtRiXMjB9MIVjNds9Jwv1fbF/Fp7QAFeBlER4LiaoeLdvii1Sa0xVMSecbwQ0TOGv8YJRoy
tLCRjE4ATv0mNHnCJBOmv5vI0VTAkY2ufgBik4u8OwqVq2W/ZbgDCMq1ZFFSdNa5LVPhgKcr50XU
7GtZYVastgfEiEQ9MOFrujhOmOfVX9evIJTZOaoDxHKtEoNwhySmtUFzyRMnQwRfHyxD1w/Llbd3
qQYPeEwFerW+sCq2dngNwSddcrj42iIge7N6kXEPGEb4r/c5yn27X7AqcGkCGY5WApI8WYm7siDs
OhJjzySnU+3ETelvlHmGHIxhNk5WYSMTXm9feXX/yTTR28C3e0xR8xzC1iivfklgzhhaeFUBVKkV
cRaCWe+++4BwJt+0XANT2fLqAth951HNzuJLXek7FXwboDsWuff9hEN+7CWkdIW2vMAv6bBnpWCQ
7Xcyhz5hzF8dwwps93dsjHRN26IjPh0pUsmt7A3icENT/Z/5Y/a2eBnhIxVUpXI4RvK/YOmg508P
LAb1c7WdMA5R6SymF8WzPtp0YW9vguXmJ196U2KAuQbGNSVm6mtMdVp0x0cXQitPZhh8/N1DTmLH
LCrgAjIPN4ijMHGssS+TnVP94V6oMhJGBueKEZFGYRcKy5KNlFwKsUCQEFdpDULY65JbpxHTICd2
nPqxO6os6BheRB46faYKF/4glJ8G7HG/s2S+zm9o1ndlmuchdJqzzMFeiuUmTKkXH2WQHT/NCcDv
6UKCLCkIJ36XVMBD67++OhblgHkFI5oXKh1D6xPpAcXLRU5jGW+Ym4kVw6yj6exbomofGKafUfUz
Jjh7jXwJ0yatGK9Th5Eezh3heYptIl+Da2wvh7CY4EvcpsGxuDty93SQbX+hSRoB/6Ama6XBSrQT
aGt5/1LOnvcaXMQopdjOD0iUXh0AZV2bxXsKpej8/F9Ekbe3fSVKM6Hvxg/G8dwGjgS79jRzWqBC
mO7I6x/aCWrxNehNX7WF7MEpiPCb6w4BIJxtv29xFXpqgKvOnMT88MLyapqZBnpKMAoEx2cUr49H
nRroA6dObN8bt+PCRKdH1+Kid6i+WA0FwOZajcUc1FQ4RcsCW6Ely/H7n2ZdLb/35jd2sWz9ZnxM
W3uSTbxEaFdVxV+/gRS2ttk0j8lgD8je18DNRgK9eqSJ8D8I9AC+i4IhnbxX1RgpRiay9LrBp6Xb
4pySs3bv9jOAQXUYXDVKTxN9fLZe+PXCHkHxpYdMHzxGF1I/6otdoc7Mebqi+enESxVeATBpwvYd
cBUpoR2XmNCdPwoPLN28bVsSk9vWN4jJC56yjgrfnqEQTWpS320Ni3GS1g4zx8Mg0NlH+TaXShBH
KuU8gGz34RyFFsi8a5hcBmqk3mJpPqQyKVx9uZ8SXsw/LzeffbxtojcVHvz35TzB3HNsnfugub8U
ACS7QehMX6lGJdXRXp9Zl9xQLP1rP7OTpb5fxl67JFK6VZpch+FmFvlx/lDkqkNACftSTKLPkni4
qZGXvZOo+Z0KFbxsTvBH/hBJqceuXx3CpwD+ET3vd+SHoT/ikzNHuaqoofWNwDmjZhig3fDCA3tU
p4dinYDQlW7xs+fjFLuqBnx7J6jmuiGVy0K2vNuyad7cxzHCH1ziF/N6a7YJnrwBO/U1Buh0f32Q
Qk6LNrTF2JZSNJsj5S6qJQcCT1kAAk2lq8O51YTthr9UNV3TMbddrB1tqTWJMIrp7wGZS6vGr999
bsirBLDakCgZOJUoOgdBDyvW/NbTQCSxeomEP3xHU6ysuKObGGWn/o/lcZ8wKiaicGa1fj8xk41n
vYRM3lLEjO4tx5Mvgk4PZIAog2/n4RSySkCz+hFlCJj2YLF4pfurUWvQy9lcxnfoUfzQHYCEpeBp
IdPifTu7lyTgC4maJNjoUJIbFxj9zCrEmyWZ/1iFTWwVNKVsvvtj4O+fX0eJZsz2KHpXwT7PHAWl
n8R3z5vWTiWO/64TdNWkSbtq9AafmCHUeJCTzc5G5EvnqtTKT8JI9NeQulanm9/F2wIGsgQYtPFR
tmjUnaxfcdWl0y+SXOQVK+fOJxETpPWfYnChZ7L2Ci6AUeuqpJSg3fZKkKSQ339/8Us4C7fhO5ST
auNN2BpCXlSHw4XWhk5E10iinh/Lqp9hI1inI9PokrCUOUgcExdwiBgjCAgjVlKcrQdG5KtHm/iY
tM38SGmanosCSPB2A0SI5u+heTSageKWyXyqtklaGwN+EOUZAyxRsD7gwswYBQ8nPSq5rq4sl1k0
H7NtgTF2glUpkQfCHhoeTIWc+DryqqBczdjE3RSNJuJegISdQW5qKFgP7nRprALUQRv7Bi/biY7Z
W+UZhQqv7goflgyhW8aBk15HnxFXweyFj5wIvHdyGDuwqqak5grlpbFk5h9wSa+jybQ4YJBC2/H7
tfjWRz4B0a8ZnH2SWMD+JERo4XTARsb8apRetC6kM/4iqAPdIKePQMk1lZYQrdeqUtblgZOM4ZVh
+mDeL66chekJd036yqgjmdqNXgV2pCfIPwizRFAsaYUwHB1ELrxx0LJ6vW5sBSJMGnfP7QgZ/ePT
+QLI1T0bdtgw11atnQaM+oziLyCgCn8SkmHqwmTv1FbxDAFc81iZvr93EueyCSf/BhLuVTuf0lhs
zDJVAMYQV5KANZY71zm4PM7w61pA0pEf1KBixPI0Ep5ycibVkIu2rd1jZiX2Ub+u01YsuUWuI5/h
6lKO4L4gh2HN2U1eaDEiFDq7WB3aPqM4XCQVdw+vGIURniBB7qm2iarvZuORVdZK/nKxbQ/3gyTK
c3h21hZfV49O15h9rNVJ2mGwA4Dcni2A8O+Y/nHSJI/ex66t82TJhUratLlDEjDgSbPwk4TyuEML
mjiTZ7gtJuyh1E4bD49Zs3keELG9Bfqyx1x7jgaaM8aI7+QCs2cz/6o3R74g7NqVw7VKRsUqFqIk
Dvz6FXDZTBgNZTw4NckkOSdO04jvXMpZHCG1xjrwstodHx4J434NSbwvAJoOAjHevkuJ+fuUw6fR
AXhOCpedf1tzyoyF+fK0IZm9UDmvZ4RvSo5wx3aGkp9Fkd7s2HUvM0YK1vTYrfvFVB2dWryB+z+S
fbClFplRuz96klUXY3XPwy5utV9NtmikK6I7YXhDtZF9qtvQSdGk5dknc6V7nP0z7V1UKi0qqBUG
LeiehgdXcNBebaikoH1z4wzgeLtCUZgYzvivjWuRrGD6UtCpjG/W4Qb5bLy+jbImuM7HWPHVsykl
0nmNi9D2Rm5bpcQnAGL36D31m5sh2sa6Q02SP22TStXQkfGwGIf9iUygHcHfdpreebwAA+USm+RJ
lZ/gWZy1so8tAFs3zNCNinhADQMLS9sePUcogAXuxQXNoy6CflGLwIy/msru8o5CY0KrTgCY/KVH
/kfNIuEfDSMxDEx9BOb4sz/34fErcw6Xanl9Z2uLcs+KvF5bTwpWVlw0LrPKvWsUhrmIwUa7Ejc3
Te1yyfuBiI8GJoQL69DDucqelbB+qs0B1FLjPKGFrhwB5GH3IAWVdmCMcp44GuCE4bJnBuIIDePD
tx/+Ui8qLmhRAZY+mAu7nRqxThzl4c8I945kiyyTWgb2DzXRiaz+P1fj7dKzP3V4AATs5w9YTzaF
nklMvbXsyzr7HTC/GpC9AIv7Vmk69E808U8Ial504vBD1PazP4rbW40KDRtalQf7Ha6J2due1/5u
rAFaXae74fiwEyoNRrCH0nvwK6GhYP1p6Cur6MaaowF8XqILL62NJNPUXkPD2JX7cx6c2Voq2ZwD
1/YiVO6O3/4rfXEPx0E3XNSs4oVJ66IX01Vm4UD5jeDVqbce3/aqV1tjzjGRliGtJ0/EjscKC+C4
JT4MOi6IvfatTKqtiI77KPTNnxoGO/0Tv9vsxZzaJQdwyQ+nVUBANbjdYppYbtHeUB4dSsma/DSE
IHpJr8R2RuiOa6NuyvpW+dclQtwLhpdy+L+BdpCYFgFHdN1V2jjiF27Y4FqRsHYfyJX0kChhzdFu
yfTRUOEIbtQoxOpe9P3rHKUb4hqwxcH0pW3jrE4gSGuN29dGIIPMQpokXDXhnBlm3/8E+xrRaIYm
TQCIOOyvAwPFpSM9uSsrSugNosEnOkaW4SLO+l5VDMYZU8tvSAL6qvE1qHgtXcoWqQXKdt4nC5H9
2NfVcvx2BCT7R+3imKrbQzihPw7l/19TTudRGGteyB4xguS3tf8ozdFNIFv0J86TYFedkvYQGoL4
LEPkW5w4D/Yft9x3oT/gsBwR/l3C+PVEMA9AX1hXCs1xvSYCFNYkmGSCBMmQeIuUL/hD2WDm4fyT
UmYmnilTHHC5JfRpz6NXQOaVuyz3X8NCYyHlu7a4Q+NLhvFKll7XnrMlP57K+rbOyfqzf7Vwcqs6
R/KFz7nWDlobSyBftfdvhRCWK25m0m4DvmUJykTLLXM9sBxwaNRbowz3AmLissjgKDSEd69cKp2e
02RpI0vRyPgqoOQPRbXwdMzFvNDBj2Yr8xnGJYr0SJg0OlGIyGCmSJPJSr3EpWZQHGA6yBDuaiwz
DSelIbA7UyHmYpzaZe66TRvaXrc15bmw1Vt1SemAPyUen+iTgf1X16jiZ6tMrnSH1ZK0/kKncqQH
FqFBDo+zD4WHsLReHPoySBPssnap1APEjSZRGSVkQ/X2BYALC/OIMnDO6UFXJV8TU97Tto+LNQnK
gKQaSjzMktv3lWM9Doi/dTzVUMtw9rnIfL8gkGXt41DlCAvHF7wfJa7HSfRiAAN5O/zG2teRCSrW
5RBlRxH6BUHwM6EQ3ZZETxzTD6a/74Tqy9uzdGk3nHaAZtkNzxOXIzQOOWYAWDEG4dyHTZKW5eMZ
VqItHsHHbr+GoBrueqj16mQ0uV+G/FQx8C6UUgIrI1kGHv6MLRNp+zhz+cwXZpYabMmpIWWQQpRw
qgEkisdmEOngKWQ6QTKbjQyl0rf4Hc8fHXnbZ9HLWrb2NBZ1t/hAGVaXnGACjzJ2AlJRJoa/OOA+
6LHv9sp2LfuNDoFs+ZZ3by3pDO8ldVXzK9CFe8OUkjpMEccEtv9JfwUc5dON89gonOYrBgrHpk/l
FR8gSKcVJkXbwzePPsCX0MfaQvdkrGTKsHtcWLAKLj5r//3MDcUz1YqoIg7XuHg+ZJ0NfgszjvZy
utWLtkMJyegOhp+s/NE56F/5/USX3PVnIkR/aHiy9qg7c++MvYK52EL7HERwokhEeOQgnlvZteiK
V6K0Ox2aPBCEx0RasmuPBG8EwtY1zPGo6BXca/vAZxiI+1gpIqlRuBdLUUHqoah6+w1gY/DY2fnH
Cw4Sxgfy26jGiyAO/A4yoCZGA3ORTAAbe5t5rtEXU6EvshIerHqYuVxh4GraVJ2xXbc/zMq3R3Ca
RtKzvnvCjvTp0Kx1xJAKkmoGBgcFTDGFGvB+qJWOfRYrJU2SoSNIgMEQc3XLfoxshOuEUJszJGqV
+jpJ8NZqTjKZ15Moa2PwsSAY2ex4vta5445PY4gr+2JktYni6oG3WQ7mPyF18jt3O2wCE7SvpUUN
FgakfdWNZu3i1A0d21CN7GibBnH7k770FRXqmXp6GJmYB+LSmcXsWlfASUQFEwmNnA9FAsLuJYNC
w3aOJTxon1I9r4zI1LwV9vh/eghxd8zoZ4AvI8SHjnC52JkMNpSRgwuibeyDCj9zdD367oPT2bVG
yOmBwMsUK8E5poXx5kZMnjNprKqbY8eJ0gygzPEPp5S0hs8n72f+vA1d5Nj4pE/7p3R6Qrk4JuC0
ZmHKlG9EiM/JUMCVFukmlVQZlhMde3dkUyavOGMvAw9vgHJlIWEYub4azPB7jGQbL512ig8fzqaa
WVnBrEa5MKEZqGSarFctY/S+QMmBvuYU6bfSWJ/d36AxEr3WdDNJB9dAcwtnAtJRCI3qnPT54C35
Vm7FQplxHipEkPMnBoBtF7/Tlloi31zkMHuWkFIFVHVRqVMEYLB2ecBkj3sM7QmvsuuFtXh3AnQ+
Uk/TPCiF4qij01J9MNzylVP+mn3l1ibWEjcjw74eSvA9rfqs6mfp42Fb0/qyo33ypzT4XCQqGGBg
l2RbENgvpzVnyKEZmBg9Kgi+frKD2xNpos3df0ZjAqmjpAdBiEvQdQ5vE7qDrdRrwgee1mLw34i7
iShs2MfRKldgP2WNd3cBJylslTf5zjzamIouNXZiQ00RZ4ayvW9kvTprJ5VDzOEH7U9hsDKIX7+f
CtbowCnJ+vYbFDCIMc6WzfEkq4m9fNHEWvw0Q54pMHmbhmu9TSk1Rt1NAWMDGsZ1YBr1m4DWMzsW
7pUJlApP71qisQxEM44AoYCx9Yf+I/rZkwDoQ8s96b0VkYYLXC9TD9STW9ZHQeI6bj6ipoVH3Aom
e8xMRIl2VucLNLNps2T1tarUUYv8mLpS7jNrEO9Zmpx4RUzzIwkZj4IQ+YsyBeYKFxL2UFqKsyGM
cxTjUyVzt15PfIjJBBOwlX2QxgFNxDXAVVWv6J/yOC1Z41eOpinTGjTieOg9Qc8YzqGWDqYQa6Q9
zKB0tYgenZuYVHAXyEV2mR1/p5hXKXnTQND4Fc77+ybq/rmJWKTZvO0xTiu/kTSo85eUItpAuOeB
yBkMBEgiYBOCFP5Et53KgocsWu4bV52VrWHnG/VSDZTsCXNtdoRk2rc9qr8zIOxOHDAaimdAU2Xc
+NXRlQULcleFNIArdAM2FC0nnPZf8Tqgpvs3/OlhYhAvaWYkvrHAQzujWOtbPT4PCFgGIGm3mJK/
0MeRjXz5cVrgbCwvYQeniOjN1DFt64mBGPtN5ladySmxZGmUCC29Y9ekpIo0S0xsN77CauivPL+D
i1Tjxnvt0ybMpbj058yBzHx8pvNSBV/v64u8SyCfpcsjYs4l5mhiUxYQdHRUBCZKFrxSN6ylc6Bc
UXAbENO+LFBvtR92v/N1sxThsgZWsJPo5YPsopkysp0OznHHcKxUnyxj3K+tJIGvpTZjoUxw/qhu
EOFHNf03DZjOcYffR7iPoI/Bcxh/Gmsc3ShtGkgJ3JFpPkwmAoax3NOmwCTp9hRes3fgZgc3LKE4
F3mXi8ixsgeLhP0HqmF0yps/YKkb0GssWvWnVwB6W5UjkQQqOiCSfOj311XnrKCT6jUn24K9DwP9
IWHn68QWjlxIDWbC3HzkLVvR9Z709rs3ruQzje3ktR8OxvKRaIKj/FvbVQwQYrcq/VaDya2KdGB4
JI1rLh+KVAGAVPU40bafJ6f9E+2yeVSJyIpEE1oN36UN3X1zRQyoRagWzj4OUl9I91rROh4FRRnS
0i1ailpkqofchrQCpBwKrtyzws9EJnnEUR/fEs/LFpX4ykO/Ppyz0CptX2lkllGD7mRi9sieB7aQ
D5kP4ZD0lSILtJ58TtkrKHrxZOcRAvWWwPeDR8I8xT2r7Qjq544vNSRxpm9UO6wlZI83yX3dogUZ
FF+cN7jRKDyD64uOLEgnTacmqr6GsKOZ4XhQgxYOSWGeM5Amm1rmc++xXlW5fude4RMsiiXfmv4c
Pns2/8ns9pLn2BXTTacEUE1g0XU3qYyrhMxLdrCFNBoywAzzyz1CJx/O+uKoBDFIjFjLuBBfFUVb
YrOkS5XG7X6h7dBfGTtGwEBvgnrjSkMCbXuVsTETwu3szENSCsYG0GFl8ruRMQLC6qvcCUX9iG/s
wRW4eZMZwAtGxWa/Bkm1CiIW1evA5i72jouRbwZUYskCCBZgkNesNeXfxdExF7WZNFtM45HXIlqd
SqzEpEPLMMBJTP6vWXddBhEzeq+w/GwvSE/AkK5ZnXy0UL+SYEHSHNdMWYFQNEFWUHvv4iCZrUc3
Dll1+Ny40GlOPsXql9gm/l9keJRjR2x+5o2vru3/zEJoqm/4qWjtylW8oxn2xINFbtuYi+gYjbq8
ZAzXwkx03Cn1w7dtX3FGmhOnXza/jazJcBrjDS5+qbs+QpwMIiSPTIeH+K0ErykJhra5sWREBxWd
seKXjXF2jUNYjcEGb0F+ThZHU1ShjFSvWwMnXEZChpRCpIkQ5KbRTNuE17OynpJ+xhsoo6SvsmMZ
oclA9XpLF7HFGu+w+7dOZrsGcRST/+dv69b3Zt3UYbI6ArlmFtvzgRTL5U/fGwO45lmtRGMYGCH7
dqs5W5lEgf4+quKD2PutBYv4ctd77KCHnX3W0cXm/1AJMYod9eQWdOhe+JH9cQsa76bPrH4iuTJF
QrG80LHn2r5TVr4VlWsM/I1kNNXhoAVBqeZ+54P1vqFbGJLGdADBmx1DGni93ZihKEaOEeavtDBE
yRF1eIATNEgIidMYcBYGHj47UINslJWkW4y/3nf66vGrqoDz1Zhc5g8A9EGHGZpaSBPenAaLH7BW
R7rlfxbQQWRUggOz0HoaWREKPEhn/1mGQ7GVMvMDCpfSEuyRGUkqZGJ93++uSuScq+ql7NNALF54
6vHJZduPtjOWC3Ym7LovS6CZUYRUD8aCfybSEk8nQDCP7LzdmhA0JWnmLfop4mLbT+ofdDFd4lwB
Cc7W/ltOhX00w4L1yQfWSt9355TvbG0MVcyJjG3rtJdiTXXbA3rqtAq/BIize8kou14TMg2aibMX
hUeX3bCV8zbOqXFRue48WqgbzHBGPmO085iYHDAbdR+K+pJtMMUOmWFm0Or91ErXkxmESPxmHM7/
aLVpgyjXMY8TRhUHhkr0W1jBa2Qr5adR5XnhCfw5R9siUiZIMeK53jajL49yp42O6aHOJFMX8tBS
dKgOvv5UNnEAuiie/OE2fKjFlDUhrg3Kghwwtx3KZxNP74RtDTJ7OUrBbZs8YB5qZk7h/mxQeu0W
/AnUoDkQO5ZGWiLDEuNPCnQMvFDWl93cJf8cmYQhZaIrsj8TSCH/r55maVh9iGKcimMkwgafObfM
VLLti2CCL25L+m/pj8k70bS/YChFhjglg/bZRyyt9tHFtJa7hRWp8bNZqVgWUEnMuDJCxTlgFvLW
C2UWqdChcE0y1aPUPS+1OJkiUi/pzAUEalAfaw4ecynHBrB/3RXuICEk3Y/03R3PW9ZOpKMmlpDP
Mq9ku3fohXb3/90r0gbCPEKkTH0+L+c0nKUkfuQ+fRj0zjCMTwH2BCFyVE1uDOIuplyxRGWu2iGd
9S5i1Mm2imGN6VKzqxuoGAg0IPeNCq1FC50EYHK2afXiPz/S/laAkcznd6NJEvRkp196dtmallaL
ypkQ2LdJ9KWf45wNAQAaaoOBei3PUzrZH4U2hgegEme5aGUFZY+ZR/Cch+xpZ4hkg36wyApyw+E7
BEPu0pmyuXPylgNj0XS9c0CbH7Mkol5mvGPkvsZCXrXJrrD6tKWWoUuZ37cypPesW/V+Xl7H/dpO
kUQRFhFOU2ZpsS32CvqJ2IiYxk+Ai0zldrNZIj6K59U8jJPCQ5MWIp/cIDA21fbHyzqLfuX7EDBf
UL4dKY0eVLlABJ2FT//rc2P02wlwfTHOGkLv2NS8/xUz1jlk/bv/4ezs/g8xeATIhF7kVDHzvBWL
p1xWQ7LQqAWnqUGxwKzMzFKkEvLbKm1rY9vRUpfe0dDnAJ9nGxePrs8ngdUBeEa2S1f2RYbwvVun
j2J080/k5MtD1Ei8ujlp9z4HDh0DDhYtPvdxnLcw/50wxA898k3hvxkpm6AiJVnS4RRNuJ8nMzLV
ezOCRauiy8uoQ/znKSnGTNRya5q5DsCWDCL1EzDWz1OtwTvgxPMhm1nEiq3KDt8AwkVL/c5vsutA
CfTUCL8UnafPWhkeTvrR7YatYSYKoDkIFYn2ECBPRMQJJHdTaneSnHa2ok+soTAMqBss6llEQihu
cUH37XAaetir3eOkfeMhrWs+jRZHw3ixu+P+5cPlmZmRNotIYeINQhr3v4Zl9YvtCsdH8kEHrLMY
2nWOT3g5myVVPEejCLK9pc4RamMtUWSNwfGg24R95pzPk0WPBzFTqUHowAb9gmlBSyWikCoMdS7X
1PTZf78mdsdWbMJDTxHiBAcoRM7/0rSFZ3HEYc/gkSAjcAKmr83z/KtLJCKMWF1j/fXYBrZCaiH4
JDtlZXIeqbXn6J/XntMKdc3Eu9hReMSdNUiWyX1HX5j+Gi6n8HxnoHlILAWu2D9ofW6I/EOQw0kK
5PzXeS8em2PdxlcPULJ51iS+miykWkyose58qglzTikU0lDTvYlv/+Z6H5i9pPTpdEeNMoTXTW6R
FZWpv0AVDfbFZ04fhf9jePPQc/bhWNYHTMPOIPrf/ILfnC+7LEdj1f2ocfHpSja/YHb/9BYNw4q9
UzyJq7/FkIVGaWk8zz+VJJZy2iWNaHSSwIs9zAPLJfPciE9IjvP9jH8xeJNoUlosxRbrMzizHEUp
JraHWj+aAM6kei37MRuQCmlQMt6NBJiR4wZvVXELHc+A5dim8v0BdkxLuJZu4AsQ4EyyT1j1l1b2
IimFDkunCY4PZ6aRKOYCkIgmqphqbyffgSVMfto0Dn6txJ4SBzRJPLg3hNzJ3ADEORrzXNt2yfIO
lm5HAvJ2uuiZyggeGtHrV/fDN5ECuR4KmgFnzZ9RbNDXspHM1plP/vFqcJMPUiUIvapQEDsReT8N
KjxMz7LhHkN2UkHKSI0mKnPpQcmz+r57Kgwuz5WVeJ0OOOQ6bxH7IrsX0RalVBnBot1W8pxL3nma
YMpmk1BRRiwKS0KWS5X8cYxV9KESmUw02HCfFh51FXDFRqlPqlf+Zv4eMt7tzKAi7x1y1G7Bgsie
u5/LvNLa7Xf5pqnSSa1ZRTMNUBMgZT5dohgmrwB5/wNEWsAZgw68hjRl0HDFl/rydHWzrXIF+Tli
ZR8sxfzvyOpskbahlOMPhg5c+zzBqhM+TdeofBDjHsw4apKnY+bi1TFS3b/tkbHsDo6GaxluDvw8
Tbs92is8qEdsOtbiCdfBosDIemjEEpss76sW9FFOVpIDK2zoYo56fDBpsUBbIn97x9b+TC2RbypA
I6OsgYMely/Tx1dqtc9SYU+wvnGl+EaR6P0SVa3wAN9STADoa43CBA1Mrs7768mReC1tRVk0fr4p
/9OHIV0jTsHnBwc9n1eUVXkHsx3wZXgOG5pwD1iyPXGZCttgosSPUgmJ86bjhQ8h8TKdo0hpSt5C
LqhVwCtrC1nhYXnO4NBNAvEQP2PDZLwHwtdr6Cm/htcQxXT4S6shGOxr4mtiZIgDgzx2dzabs4Hr
A2hNvjNWzf83MalCmX+OTxCP80vkioG5+iDdbicHqlwFqpFhyiRAlTXCJlDSraKHaWkgzJMQClZD
mdgM6myUllu/NfwTg9vBgleXlTF0ygaW0XtAUlxP88aUH5mgELpwpJ1OxXemnB20SAJAdhC93jrm
cT3W0UE2uBTkVE9IfenzQMqqMTk7HVWTPjBXSH8JBKahZ0bkAH/8d9ivxevHWP3gbsj90A+WMWs2
GTDPRN+XHWJvcAWKz/L2KDXJIQVaBbml3my8fG+LJgl2l96V2jAmC5JqPr6CTJH+S12VQnSCed+S
THYsjGMkiYgBnCRpUUE66JLchxx/qglaK+f4OHD70Ru3Q6OsOoN8Tz2/ZYp52lxbN4zoRGY98dMe
SK2/FJn0PRaMO4FNkwD0/5EtF0tXKKqLLjsaRbQ3z6kjJdm0q65x65ViA/gig+HyeOnhjz6PKf8N
TelL2g28JjVNUGIKPE166heD/AjRjJMUed3qI0g/zDwBrwU3BM2clK2AebpYfw2p/zEFVi5BVC5Y
/VA2Y8kd9LKEcNoR6Xx+/6GCZkcBedBxXnlcUGQXhP3JFZL3GQd3a7fhYW1x0/v+T1KT+hrBqQkF
E6SCh0QiIOtSYlsR134tURfJi+a8V3wVBKxW4P22jfrZiHUntvMBixbvUObcvKnH+z9+IkL1DP9Q
gjHK3T0Q3JWIGo1bydpx0wvGPPgH57kzq7lfhf10VDhkoE5vdQvluvpfXqWJ5v6RcoHZw0Rz2+AL
tt7pTwjjGVospTg0YxGzNGlpo202hSr9pXVMAiTxS2aI2Cwa1WcFczBPIteuANnCQKqXqttH7IAC
GwSNFIh09Tz3j9J0WOHwkZt8+OSwSYOa0ncB32sdvjTnKPCxS0y6p26a7U6XppbHDgBqJiISkVDz
8X5ERbqmB6zfceA71q1V8xU4SBcsRnUhdz8w5jsU8LJswyrm6gyge/ooGSTU09OvDldF+Km15lZx
CMmtOS11nw8S1uOUjXlo3aGhTWCG9lppqlCkztGZqfNd4kvp1PVWPsprAUdxIgn/n3Ntaee+lT6T
SU0gmX9N3cSD721O5yI2DUua16U+o+HtPdpAYtZtteFBPcEDCnlzzjXU4Ie+QhXbaET8bUc7ELab
DQTVG2bKIeMOycM1Ru11RCffPzsIgls5RTfsRXKhxM+jRkR5xUceu7EO49OkJHXrBfNWWPRED4Fx
4HnBsIvX6rvEzn0WGRk7ukCtOJ6iu3rKGdeB0KCvtZzNeMqyfAGOYamfYmc0K4g39o5d3XwQRUhC
M8oCVhQyZOK+iosE3i/g/YLnUFhyZoXvOCGNvcx/itaRucqI34PjmIBFguXWLRyYOIG8wHkZyQL0
XjuJCeDfyFrVR+80XMBtKJvkcP0K0Lt651HYDK8zCCxM16IXKkUCDbJZ54Q7MiYoDtyjjeHtocB1
yHUwZh8cK6NYpFdeiUrtONDzVzezqypmpIe0MW7V/sAxaoL90P3pmIoh6uypld7R7tMOgxi/VJfU
ix1XGqvZc9OjB+HuJi/h0P7YsouQ2seNck/fTXhmRrxLh1O7eTs1wzhe7Fk8L3oZmXvtRD4aIUb8
bZ/wImKbo+IhPV0NxSlrmJU9lPqhNdu7Aq+7f9ZtBLWAJdxicqgPCFSzaqoSPXWpOVq1+kMjrswc
gwlFe1zugfE7RUsngyDWlq1kzRL4QgCVpuTqC1XZAU5V6pAmj509Aqk4KlGuXfkY26TOuN5XKlBb
NuPntYaFHSUFhcrlK1y8+WKpiuAGwtfuZNM4N/l7bxGT8TNwf7N8qiFN+W6jNh7ng0vlfkjSZQEl
i1LgPT73O66+fz87AWGvJNW2r+d2I+9Hq6I0PNnvpfczk+BuvMLlL5rlEZ5npjdnmUTXIGJFusAo
xbaL6C0er7O8DAPDHkCx0Vv6hJr4MrdNyuOaMvquRK7M3FNPxx9YBhqh+uunPJId1BmRbxluk3/m
DsfeHmdw2V07DCERRwz21OTp8ayCJg9ZFInNB8gSnPToBAmIhYSZIlKFzAhmadSg/tiUDDQ6Vim/
CgUu22cuBjWjaqeN3dZIG3NJm2J3kuOKW+WLRbXZck9ku246ut0hKFXbrMpoCM5ydFZ0u0dDbCUc
BULLaxDcpgcj8TfC+LN/HqRbR/xCQmU7TeQS2aOikSRqSwlvNSy06vJjCAFjQDFW3MFYt6xuXWgp
QV+mC04O2ZU2gdGCeuCf+5E/g+dCDtPV/gZe8dm05+wk5zu7faPCz4JKBUHWgHJc9AzV0A/CCRw6
vrEtbGPWVonrQpculYZy1zsDg6Y4NUS6ifmNY2QLunTSnLiEEr3keOuOOAatwBjG7Hq+w/7RhF5S
Agm3bRdqzb+hmeE2q9h947IhBQkSncYOlTX5bxF3fhZoYqL7BFW5bT8JIp5MWCe0GmczJIQWHeDC
Gu2Bpaybbot2Snr7GqLjA1EFoHiUnNrmEzshZzx1S+QsQ6ZCjIdgqjbk6XabiqGRLOYmJa6LF+ba
3EfA+ASpzyJI85II1Hc+CWsRSJ3ZWVeyZAk3wlBVwxpxz7dnVLmCN35pRkVzMEPDMOp54h2kP6je
S9l7P24xJm6hcElEzjd/WcGfuNBOv3o3aMXbN+DCsp7Qu+KN4VDybd6WO3U78m0wBdHbv8pCDnMX
jbiKqZ5SEQnBCLeKaL28HKEMcekrq6B8CVOdu9ickqZvSRag9gaxD4aWI7DobjxwHJ3/EboWyE49
obCWIUnLrAmDb5hckoH6BlwyS5K1nb9TUYlRMg39BBVxF7teUrTuLhtQXByW9AHbPRG+cRoujLh9
YONCftFT7TVJu/p+wEDFoFIBvUGXGIUZoa9TdG6pjtiOTIGFQEJu1+9YXvFpDisr41cBlai27Y4q
dgsRi1qfXnvqGPO9Z1x5Wnh4IhxeSLHJ76BwdypuG6R35kVhOGppWz1uMEJN1cYGs6Y0yv2bK/9d
aAGKjsUHb0mVfM6OmTQIFJ6PPyt0foWGwhk2iCDT7c8W2Isxbw8dM5/ZE8+mdbcjwOne/U4jvUno
eKFCN/cNlFjLw4xFr/cGqF6DkBglo9vRse3+aQ7bz+iQQe3e03gqSkcaa7rR3jhtHGK9u+LWPH4B
WKdtedAeFqB0AtbHtZF1xs8Uf/lRF0cCe8SRhzsLbApeIiwB+FMx5GaJSw897cwdP/RGYObg8mzF
KkUggBMJsWVK1SC3gtXosstejlKVzLpE9at3JlYigGetQUD6C57GEem3L1j4grw5HoHedplwxaRn
ldxgna2314X+uQSEcvzoN4y469q3UMUvGj+KTGgErxdM+01/r139zLmmIU733Z3eVCZ1OiKH5s3d
KAiwKtKYDf0Sr9jHGCk5XPgRZoHgeqadhvP8JHd4hTtEmTnMRBh9LLZLk4m9ci0mPtfoUmBF9Weo
4AVei5iiQ6r0kxqbquukA2tWt+sAjZG1pkInaVXfp6UlUJNSI9mPipoliUCHNOnhcUifC0+4R8b1
uSXy9MgzQYK1CVf9HdTF75pBn+nCfvwEkmWMpnQy+QZzM7GrXBf8wZR2fSXEAFPnQw9/NK9T5ALQ
Zcn1p7gqE5sH3nN82V6S6AmKw+3R4FyFU8rUlqGzyjO4DT30aAypjKzkLn/loCFtCy78JqwMps94
RzcfCVseyW+O0BoqQ4gWH+mfAoL/ypJ1V29IqqjAiTNlW6RX1R/yaOOP5wd9GQApJVMBX8UlylSI
uzYkNSLZ72ln30jCgVgG/cIM5xFd8VODQ/1xS+qJ3f4F8E/QbBO38GIQpsOMaA1eNEhg1COehWTX
xcoJozstBfdLQWrYerIZOP2qBfnQv8Rjz4UuxVXyNhn0bIb5+JxO904P8DqsJMIf6DqfqW3qdgMM
4NYjrPFvUkv2I4fA0SyAKZVGBybGkhTkMiGbTD43d9K2yl1p74EnG5fYs0mLTAY6KZlBq/E5KpPj
Tg4Sb0yZQVK+tHGV3G/qbs7apWCpNqs3VP/3+bTun5qwU3+dqJ+FAoQywwK4SszbGhXJ2OFG0GYp
FKQry49oJ6hWK+hdIvHmXxEQuxpbUFF3CVQKwQrtO+YMLfmQOS+xV0XsUvc8RAGP68GHsZ2PmAGZ
qDcqVozZ4bqjMhoYWiG8dmBMcgqgXp7lQ6QSA4I0xkbenc+KBf2g8tQ3YhaGD4CGzvftU2hDDJmN
bxMGRc7lrKJ9ZvLCzJGz1nnrP5U9VyGoVu6QfwfUiyd+XTx8egrrb/BIHIWrheljejEdgYvctlNB
QCs2/VmiVWS1Fd3lxI+oVlieLnTzx1if5wQmDoGt+3F8AaMLWGaC4hEMC7ZoPpGt0s1Sa/gExYFb
vw4WA/akon6RtBKY53r/+WrVy430AGaBdv0NCR6+Eag7NSKQVoL+jQNqo5khKaqpWFsyK0GtGtwi
W4CFWFdDsVBBaYeDLsWMv68W35nNoY2kDhVJiUiC2YL5gL7v7ZTLPHJGGtLVKMjzoVwIwzFDTlWb
8WBRiLFrwTmG72uif2LIhAs76hyZMXV+aMgrscKOJiWrWIQFHiVe6FzHPMyZJ7rGiLanHly4wMYa
tjxds7HXzZs7WBxmhZhppvdFsZv4LBCKg70IL69hGSAmJTbN3erLlD2lIDdF0eGhszdhtvDboA8D
tPCtaMjZoj6N/+g70fuOpzs2Tw5ECI5aR00yuIQ8OEHtRyO3fn0bEHY5k9L60DOdnEh29jHXhkj/
2AlTxwJpD6yZ4HrCzCnyj+irwlTigAiIfx+fCcx91z/l1kVuBfjVA+1YzfJIURCl6U7uIaPDb9CB
X9BhOBSXRBKcQ0xC6Yzv13x4I8btIBdLeA0DfOLgf15qulYKtIEdliu4D8BB/gxLgsJVwrFONzTJ
vH57i5F3R+f/M78uu/wPNj0xcpT4zG42TY4JRyIHSWA7ZYqwuXJ7H+xOKhA1Za5KBxcvKyVbbW/Q
I8ZEnRy5pU8RG4ZWeuHwSS6WyUpbufS9P/4+OavIyTWZW9evkJN7U0CRENldDqxERq4nbg92oI8U
ZNYL7LftXQ40seFmg6Msa6Dw6c8r4mZq+TSaozLp3Dkow7k53EDWOxNlKjB7+jiH8aF7gj6x9YoN
Ve/j2K1UZBEZfe21gzJvzAuvQGO4nY/hJvqqqGRwAFpZg+sz0NYz4bXdNovf/tJALNqVDJ8IDFS0
Ayg+FxZc5Rg6M5bdFwkLkOgiks7VMJWZkjGuOv8cqFVQZvoN/uBNAF4JYrCejZu/pP+TTvBELMrC
1B1T+k2PcazGVBfKfr4d9RdW7kpda8XJCZ5yClJ3EmH04VLGIeWrXI/lDK27J4g8vmdSQL1I2u8G
bSxeVL5RW/JqaZV86Zf3IzWCQVpWcgxxv9RAAm7k7vBqzon8F6B5vcuFlWtp3eW8KkzRNSXgIAR0
Lo7YrKg4OcwUyEDWoZ4lKyD1BDN5LjYkCDABs6/BK0qRMwTEh2MNsuv1ftdQXsM8IH8PanvjrLbA
VQ5sFGXIaGmi9gpwlVeXiK6ApUReec2j0O8OvWrbYlffSrUiIbYN8LO5zKe12GiM6y2ygeHRiVLa
VG7W8l4nhEiR7e75oAUrT/tHoCPEvcWaW5p/lidz3z5336X6yPtqtdxmbePUT5dwQIxojTKbHozQ
xHprbrHutuflB+xDMv7KCq4D9Ihs4a/zX1QZDIziuHmhg3zUOnyEJldgd/C678QG/GlxqQnIU/uw
YzrvtAbJWOUDPXbsnEU3Ih1jsR2XXnnRlqZEvbvshCjeqwAFEWiX0/oPo8qrOseeOQAFaLRgnIGV
6hBjTV8kBUmfaz1D6Otk11VLmfPr+acODd4oXSbVdSMgywcOpytmQiDS5Xn/R5B1c3cfO0JeYqNL
w9ld4Ac2X5XaHbVaGnGBheeO1J+74lrN0IM6WgYoL5aZeA4dmsyMblSCbtIJp+MNRRPFLfyP5OkU
2Qi+HO3YKAu/kZ3qs3wQKWrWdrLl32rW+oYtKol1DFWzs6gOXeypw8o+IjLnMpLU/tzeQRN0jLrx
fCazJYzH+utiSVwadnuVKz4MQeivg7PezNR4E0XdNTm2PbfUDk2r19bbilR6RigRYJm1JMo4yxW9
hKCrl7SzvHZpQWpogsWYafOJ11sCoEhIEaRypIKwx5akzSoFFP1+qkHC7OLQz5GgMTgGwGk8NxoF
4ovXZURjQ9Tq9iDJXXCmYoGDQzITHEJP6Y0eYQYQ8QlpEewYnZP+8kpRYILNydFqNUb36ssg4/6g
KcxQQ5/poHnPhKVTrt3ua1aGbwtBvDLf5GNAVN6ne3nOs62Nm62gyUbS65LqwedxcLrmgZ7A046U
5lsPgcuT02Guy5j4CfCXgSqZNIHhQ7NvdAIx9NUjNGx9lGIqDiJgZYJiKDr27dG8bww3ta0MFbxu
anidTpFzIK+cKDPwmhiYm4ZbMov4tgQRIxsBb9Sp6kJGgujPPPeoQbWhKTuqttlYVL4PDug0dPf/
KDzvcrfukClv+l0hLpRQB6LVWZyIEQsnKwrpLiD8wMS/GoTTiOYvHZT/fg8nE+pzhxMMXurAhZrV
tOUuwowbCR7bWMTLbId1JXY0uz0ObrlewnMT/qSX4mt+wCbPfKn6AV5XtegawnJBDWelp1OoLPSm
x+UmsCKus1yfIlOdJ88MWzYFDViQjo0IxeGU4eXW2zkGcwGTXjGUPLfsrqybt6VWwKt0IXc+Gv96
VBs3g+hu7dfMbrzrj/QdlscF4iNQv90//8VeSXamJLcDI1gIj1jhu8LP6k5rmYSpP/BV/y5jCXaM
x1dyXK2yOpYcFVT9K9J2yxNuKoA8NxlNNo5CGpCrdGiUZFILJi5Mxfiav4JO/On6BWBsIpBpFv82
S+pZLn60sjvXTOx2IXy3Yh5rKMLZZNXfWOqzEWi1owWK8kmw3OLEQbDuGm4/seLiWHK1hkTvsfbQ
PC7BKKryPxBev3l89PBJpa/T1F355pWhZiGZtMi3hLVDcH1Q7nWV9i3LsZTOe0aSF6QKM0teKS6G
Ty6VWi+orpIywCWEp3pBqxMhA2hrjdOPute5Q6KP4VxrFQ9MuCqC9/wMGH+LRhJ6SjL5w6gEUAjy
c1s40zt4+3wtRT9rDQuvUXovzs73YoMb7/ZMH/bH3tO2eQylNIxidvNe00KuIxx2CCcxlvOJMF2M
orTgfMhs/i72v5nsew+dNnCGZlLe6hUXuOuU6hLfJGmM2hX2vb9YJTv4Fb/CiNttA6R/d5M2OtVy
Cc52eVewXdRAXAyBLxfn4h4cozW/OUqJ8wiVSU1rzbE7Cp8675U7TWP123Ijg/oBM7awKXGzlZ+U
zNZdwSdAsWmdIbRkv/6uW8HIvg8lntrv5gPx3mJLk2cya6YJoqY7EQq5RSVMWJClc7f1Ri37+2bp
GXe//6PPoGStV1uV381MRDpoV7kAMuiFY6o1EdwP+vhxZeWgZsQXrheWGK9nZNlz8J2wfj3c4Sa3
9NAMvYLbrR2S7gWgkFjR3zlznshvm1zAgQLjxmFFYTTw+HrB0vln3nXQsUyZTlkzUfHOhyqfj8Vf
IRR5wNW1n2qzzb/WOQem8NfygJQN/0O+/0Nm40rRrvvy/zXeHPpmVoei8EGMZ627z9pqRaNp4kLr
VDlDX2SDelpJ7Qxqg45JqsJAtqzkp1iB+TQIsk8leepilHLMFSmqd5ciFLqFOlqTj0eqyY5gmEhk
7eqRDb601fFBc3xKP9jTdsLbg92oZuqCDVC/rFcsPzpyFinW2qUQg9jQ76iuxRJiWnTSpnRjBkqS
ublaaoHjMLCWO7+D5e/r7H3uMU4V46ojVmWAHc70m5JTDzP2XwZ5olMkgsEMg9zZMxci+8RzylbE
3su+6L4zb+2EfNMrD1HbcGZJYrB5oaEC16Fv59XbkKAEzI5QLoffEzeJLym9GUwspmNB8oVdMnRa
LbN4GA28Ls4JIa+607fZKaYtuA3bbnGtmbdt+0Cdv1vSffQMkCxhQjj0lXsqf2fdgfjY24t9kCo2
ILUYXUjt9qQZK7oGjJ5bwn8LwjkZBaU4Mg8zvIUug9B8Mf4DT+Zbml6XHBG5z+UMlnYWnhlGPdty
vDfF4zWommpBcXoSDhneGBiFyRJ+gsIIFsPHWv+WbpQcDG2oVOGvgCWvJhqDdA0IQJQwZQgEhj/N
R/0bzLRc7Sjzwuv4Q2VOU6awaM0IJoMQKcd32soyKnlOYTJ3Ndm86Hri6/Y8k4dE9W8juHoAJZjf
VqQN7yOmaTAnjdcIILNUuU/yaoP7RIhvRTodyNsc6XEyP/TbCzvI29egCfdqU+QWewPeCmfUeRKQ
7nXxU6SXd08h0ZzFm/4xPu1s+gGJFm2szJpH1lOW5TNurYO88TjOBxoxImKHQMGcVolwV3wPfyn/
pIL47GzPx7H9EgfxyNe6FiPhnadJaCVbnPrxjBBEB99CFA4g7RAtLktwlahyGpxDwiOPfe5bw4Ay
UtoEDRoFV+5jXoQZHkLq9daScJLuUQUdTvBwAbYgK+gFV8k1kS3s8V5pnAdqj5UsxBQVCsnmJZEb
uDKF/2MXsLQxi3OweOccS2OwirrDmw3wfmDxnUvrT7PnZG7HrU70qG0SbU7v11a70zAbb2lgD/rh
ofm/y7WpOqM40tSBGi0AAsSYdJM5aPZMvZU9LDnCdvv62m5ry6Fwskh+fTW+Kh5kK0kORBG1lKVS
iNxBsShMDMrmXQeXYoJ4HrZLa2UwDcbVBitaRXsoM1kj7T99iZW7jhuy2jP/ijlOm+1KyrqjvTLM
A2G55p0z5ZaUy6cHOH22uvZdtueQRyW+aLnbVkJBXfscovlKdl24jZQucTJde0bsWM2QpAcCrWTt
SvTXBByRkj79BltBLJQD0HcBlfS64qOXbVf7fNUxaMg989Tcq8rKP+/EV4A3ph507qea4ydh1822
bbmnpVlgT2fapNd06xbvvTCssJ7neCT3ScGwQVMUTU4i5unmP81jJbzJV37rwRgtftGvfOamgfdn
YdWljubTK+sQvD6YGh3rTo7b1QJBnzN6dhRl76uYvkCk7HMGGk/Sq4Ph/srCvO4H6WUDO+3g6qeT
maWLkC0K4iae5UL68ZUc5zMPGyKur7uezIefdinVywLhrH2vY2Te5quJZxkXBAxJIDUvtjftivEJ
xC5vOhrVBZ3RldDkry11ceOHKSQE1FJ4vc4mjZ5TAm9hw5XT90kSFFkDTClYDCx5Tjd2sKLGzI7K
8dvOUn87uhEqbCBIk1sYPewb77TP6t3SweU9CtBjlnq6mNczk/75+/N5Hpxf5AW+lVpOD4/JiJvx
z5Ie0xgLE4NVSVXzvUbAuiwcy0hVghivPJQ7hAiqR+Eh12DfC2e2jM9Mmpp+KWuOe+6cMuPARfNO
TG3pQ6jfYeRFyh2ymW/Qi2jYEoCnxEVEu8qW03UZeQi7dr1mDOTfRUvdwnxhpEmY1TMLvJdzlSZ0
RepwDcL4rGen/pJyCk9a1nugRaRd27r0LVRJuignQhlz80hwhKPiK7k7LK/ruhBWgz3HTu9yyXcO
cXUyuPuk/bZqhR90uuyBD2g3y2meBC5ymPcng1fkut6xFIgn3ayBfbcv8oCkp8+bLXIqaM3HpGZ+
Nsy9tQGOyPgJ6K9XvHy9fQblEj6oQhm0Iujr24BR7s30H8mFZ6KLPqTFdABate+Nqpzh5wL7X1ju
5NFdQKZKzF6r3KJwWQEMtODy+XbWhJxLUL6FCe28AsS9frx1lbAgelp7diHZ0zrFFYv433WUkkYO
74Ro63bL3F+Ks5kDSwXybrr0rv65hbexIZ9SDUhlTUWno8zVpqRYBNcmBh7wBz7k7agieNbmfehs
bj9gf2jvQOr68H4vCiYGc4ODDZl+Y7e9b48pziNZcXRB27nwS31U9zwmZC7gFYCW+M77mgsSgO98
GL/BFTC0+/eoseXegK1SltNVUjoiBpO+xnwtwTFlsw8ZInrV2emmViDkGMmQ8yXpz9WpdqomiMw8
Is+wZDH9hKpQowRdUf8r+BsG5XS8XrpamH8GTBdlBF0fE+NA7DlnjlAE7Jj6alb7Db/ILd+Dh60G
Ldffd2tCo5L/3OIW1SiMLzyzQsi/24GMAgtbaeLFjlJ2rMjCGzz6kuYem9BM0OR+hvVsQMDG4lI9
POR1c0p0kWU4crubPQ/mfRxzuS+/wETcUXMi9bhq+de32sDpvcMCZxxZ1IEPPUVhm5ARK7Br7Z+v
tA0+q+MixyH6Id4r9JZ/C4n5DhJI4od0o26aNNrODYOTG6Ly7gbJHTwIFCTzuZWGYhYUW2XK8Nuv
EARN20ZTag2obRWc9qbLXh5NkRpYBZ10nnvPK0ZpRac7NWaZDnY0Lu3tR0bpZpE4ljUo9NOvLN3X
3tYTOtlYLwl7Sr9DvFGA1DKV/coua/0QKd7Q1JaNRz8U/lG5g+I6/VhwHCh+Un1YbDuy7Z0B6dmA
8w8qwmKaopA3l4xuV4xuBrWk+vppkLMID7+7eLdNq7wKtrIzr3+E4bmEpZlFV0ZEvkKyf48SHcoc
wnTgQj92E5hZzmWUne+uqM2i8Y0mW0eGlO1s3gzLYGZ6e7ZeTeURlgJzW1CK/md8ap+0NKPy+mf8
NmqStNI11uOII8uf27Xg6yQCIOa9guGmJu2pl7YmOYrf5pElPyK4B7pm4aUWAbDemIcGCLQZFzn2
K5tAAWi2bFCm2oM2moADtEQatMDd8a5SOVpGcnBe9XEwNLmCDsPX/DLZUuqhU5ngjAKFYbCAtm16
FoZLR1OFHqrYTDMqjCSVd2jz05NJH86K4NihUPveY6cP8dpnRhi3US3aju36jrUjWNKwrrTl2tfF
tUVU+zwZV9mTTET2VlP6BIp5zObo7LIR3MyaLvKOg7jN/jE9eU7mEAENpht5nkxDw4vrT3RcPq/J
Z5mKNU1jPVOkt9SMxZmLLQpQhRWQ7/RrzzQSZqH9Ssg+nym91g/OnCIKJkKmY2zLJswwQuXijZst
mw/yagSB56w7ZsNibTqsiEi+An9/AjWTNvz+7vIqaobp5fduOC1jFnS1ko1UaPn1D6SZp3k6qoC9
RGQ9SjdrRpS5I1JmrCzSsbP/fyHRGF1sqvx7KzP3pejeunpkDynuNsVAnCmCmy38BMg0K2od12aR
Z2KyZVwHGtV4zExwuolRpNu7p8LXk8PvfXN4W19rOH+SoDEPCU5UgzKAFAHsGks+81Gd2ZI6Vrh3
+vLS2lcs3KlvjdJWheJJ6r0gKDifNCN0A2D03gxbsGHIxjc1BfOMcGGKKVhBMszIATq5Jbwb6k8L
DckiN1inNh6gLR06trReZRzHuGIYwt0k+drnMpyJySYpYx4rlyW+HtOIqRaj4+yHp+ArQBunMYzk
bIDnJ+emCDBB+JdvdBrbjRH+3KD4XX2dhRSNKS+S1MEPM4KRXYHpCFWDLHRspSwDtozIIS78/Qm4
OEr5CFpk26j4NpeaYPkXJqeikktAp/320tv445sF+iU/SaJvmJFYWDtVppEq8TSVRyu2yydytUvs
Pw1KLPBzv5bfX83knv7CSGkYUGE+dPKgTalDlHKCdy84rEURyj5cBOuSVg5kb6kMih3jNOi2mkDR
UdydJrr4QO3A4lT91y+lF9m3ZZHYwbvHTPetghFiB3S3MeZ+UzZcfwgiN3mIzBGNcoUm8LsFByKd
MMu8Ks5WtoT+3tkiUd7ryf6YoCH3HA6MancCMLrd0+ByabfdPxhlccpux/W8vsA9KYbFGT+6F0j2
PREVTy5iwwk/prFuk4MNkuyXTDlI3Tr+QCP4nwddhFz6M38axuU2pS2dQI7uCSQ3udysRx9n5mqK
lNksTeBjjqABvnHX5i9Gl/fS9Vz/uUN/fZthfF3mIiJZsQ7aUCkfqF16j4ev5Z2chJy7/N3vus05
NRjMpU6w4zytMLGW0gQR6KN3okNmS4e8lG4zRdNnktohwohwbUBZwJA3KPzaGOy1GKFxZxhLMZgk
F7xYADPLyDRYfiF1WJKXoHausFLjX8yrHs0OXmS0nne1OcEoLjolHAfkFyOZCcSG+FXA+cxPUETV
1koU/LaQn1/CYQQXj3Yp3h2OMxDPf4fPNVNFfo3ayrWRplcAgbMaMzCv+t4rgv4x97mLuH1gMQ+8
IBPJdN9W0dyTTNI5zxtxoyFYWqs8hzN4UkOL+9/i4rxaGcWA1nVtsCkNEe73GiV/NXesKr3e7DSN
1+huNhM4WgTR/VGrh6tvfySk4FiP1a0l/HfZAQn23X30lohEaY2PxAx9ycqOZ2ymw99byofS8lSa
LqxPItmIUY3wx4GyC58rFNWx+SJs/bzfFLXlySrT/NwsYMZ2TOm+SqqbiD5dXO6/zYs/qwrIZOCx
ZXZItdQFQoO4PxCXLPR9jJKUF72SZfhNNqs6+mAn1JKdEdSW37D9LwSxTEslvMjVcdayv8NzLVpx
Iilz+oQgHW1raLPtJ09yNYBL9URfs3P29RrMy7b4hDvf1uHmZU7ReMNjF0ekY9qSdS47Qm7DeJ74
K948MsnAREJ3PhPBaGB/NTSy6YH8no+Jemingb3EniX9RjT/PXVeNCLbvoVRRmjQqnrOFD4O22WV
e+ypaDS5+rWTmGn04dKAcrsjJrbeLa8ryhFKeQiqN+ISSR9FtJNwGBHUwg6p6VuSfnx+FT5El+Ji
8yWRVe46HTYCZkVrgkif4yPe2WtOW4LB1tyNroSzBV4s0hUwtDcP3QsGT14vgBDrR5w09tpq3Zaj
Ynho3yLvvbIgg4XM46sceo3hXGQWyFXL0XUndxkQINJa4vJ3Rh32z+GeU5Ulg27WZXhvQMslDcII
5bvlgDEnijnFsIKqYnKk8Ii2j+KWZIj3B9c89JPDvojpVgGTafvCgOR944IP6AretdknvcVw9jsd
zCjBOHyir7BlXA9xngHWn0uQgMSEXLO7nufFlCPSgB2wIPwmDZwUqdK4SgfjGKrCDrfoM8wWoKNC
faMizbcD5JmsDQFG+sVgkWsqEBgRIwxT7hbXJp1gUWjzY9yx++Ib++AFZQzn6x64C58G6pukL/BW
F/EuvsLvkJtXllH9z9J9k1dSj8n+SoP79BmD1yBhLF4DEnZbbWgRSkrlHyGgA5btzSUQ+zzGUa98
MiXzPHDSzbaaFCNbH90nc6k9qtqGRFUDtHzoWGVpBEgsnTAW8hpAkzF6WUkvZNyFaErEuqIan8UO
dkW0pcaeUkathhWvaPWZS/cUJqpTG+QE+kBFb1cP8CewzItsWMxCUMmMmFat1oHa/v2WoCxep1t0
FcJU4V9DiPunCWBfg2zm1m6NzqWnA/c3EjCsMKFAmTnUGLo5vFd6/zXlD6+PTJzdGJZBR9ckQyhE
dsFrCT/LgODFTC+RhIQPWGsmXWiK/evRAq1+aWvrxiHsS5275yV8y/z6ochYBJlyJid/R9ggUfvU
HEKWuSxir0Vmvm02HcvkEBzGgWQHoZtvx8ydis3F5kPewzbgpsu4uXEryK+tb09LaW8C9kaUh58J
Wa7AUiAx1gJ0kOsU8k9KACijRvaYyeOEmHmreLt5YMzj1A+Vjz+V+y7tdFcRlmYFp42qDh6MqXhX
BRADcaYql0DUII5WsvF1NjcVZpyxrmy560txOpSYZ9Yphoi1CTKLC/6idARbk3goG/zRuFxGRJs4
UaS+rOgatrTbIUyxbmp/qQXxjbjloWS0je4VVg24Hdl8xIJR8gz+ztkmeS69cbm9YMMsaZdpWM0K
HHm7K7IOsncM3vqAVTwuGayjxGapP1SjV4zm8eAp1/3KYcnw4BDytqTOOlxGR9qXSXpg6gEC2eXq
/RiMFL+7px+cNBxPyLJIj672nhS6psLYvd7yEyA4cHX+Xo3BttVB3CQRtfj4IKjxzaYTkiv5/2vp
HgFijkxTarq9Rm6Gl4Lf4vAvtsrtWfHq/ehF7FhjbiUigbJ/31NYht5mMfKLq1iJqgbsLIfTEVr+
NlUjiKb5PxTw7rG1ONvRHkq1sYG8+wPnPxQx7H4XPOquQl0g1gyy4JeUQd/kbofW0ZHk70+y6QYM
rPQNVjIEKj0xHsDjds+gjkMKolpe7owDm6ugS9TmgAgGLKkZZZ18pXO4E/02Iwn01adIfLgUMzCz
Ci3wA9qS2F5qXyWNShG1G+Yo+WVM5Wapsg3WLudOc6iiyorUALZJemRLsSIB386TgsK9A5owVcQq
1POjymQ0YvMrD8canjKGJ/EmgwNlPBHJUaCuI7QUy9lfm4pjGJQrIVq9NOEZ7rRH0WjtzPq385Dd
l/Q8H32eSyC2NYhhn84Cj8+x0Bt0fsnRrUU+wvnSYDE1XG843EvKpZrc5MYzOKKc5IwP4EIrMgVB
pDylq+t8SAPjoTYNTf+CAiiO2brf7jJaJo6YRzXhdUVOvrSlShXoZlcBMQUuetHUY3Uz8QENKq0U
62MTaAygSnZnRdt+6spQMYDT7a0GvDFcLDWGPY3ABw8hyTdhYD3r5+xid0IfUODDOxKA9yQbTF9R
d1Mn7pvTEQKEhBz5ZeB695uOGk4wEnMZJtq75DgKUKeYkDG9Yy1gv/o6/yS5OSutAH5J0tWXpNgF
6v1kalOhYcv4vrR2GIGRA+LoW8nhpqNBAuPLrK3oj6Tn8EbOAVCeIReg9JRutbH/LwXn3oFphabp
D8GDnjsV9wjZT1QJvXnx1lsJJQAoALyOfgPZckBNJOq4+GPwzizEH9BfQsY4VmXA+hbc2Pmr58Fo
l6Q+mvSpXEBECxFRwYb4TtciypnoyP2Co7hHmOHDqgmglMevpClruxwLq7lTrlVpMEX9VRJfnoKY
oRaAJrEpr6+qX5lB/h1IVw5Yzcaf7Ujz3LO+AHVH2JiJXq5slLN5UhFxWpY223vC0f0SXICJjReS
zq6HWkjQVyL2eStqccU2pYa4jH3GR52EEVNqWRK8bOkozzDY6M3K5EnEeapfofFZ+ROXu0swkNf7
8vSFB8MesCQoJZi7lRyg0ScdbAMjRJVM20IHyCRb5/HyaJ+sJ0MQCOAoDgArr+L3XHEwmSW1QTIr
YIbQa5da2qS0FpB0bocw0cFNPM9ei9eLVJqNHw61YC7uGANkDe+krzsI7uVbRnPXuNIyyMOU55bf
XRvr7zQAP05U+b9jm41fzaljGeLEdRH9jG7LWGpw4r5iOvV2kQQOdZnoGAsODPVZ5k8HlR1HBoZN
7CVeQLGLgWYBYtnFQwcuJ1PDUaDNhWttNxFOJlqBVGsNfDSc/fZTI30iZXatsPAAzqz4qHVwnnrn
E4s/i1UOzgH7heYskHOxyVXt6bnmFUdjXtidEc49dc+LhAm5/OhzNvSjd2ji7qX+VSW5wXTg5HBd
790Zv+OcT02RNP8++XM4nG44MwseyOhJE1+NgeCs1Cb5M6d4mGaq/0lDdun5kobtnnKgASt+7VVo
qijJcvaJiogluU6XkSy1hyTkJySwtrpcFF+SaXRoRMNbiqiQ+1zBPHxQ94WmmjtVuU8x15M0Yfw5
6qsTohxsCZftDJi7fsLM8OQ0CRej1jtuGMpRCgaXMH4crgz1sshDvLi+i+tKGXUUGbysytgaPMfp
VoJf0Vv2ylLb+pB8x8qUJtcyMwPxXqKMfdiCSVGusouwwuEKMqt07eR/6j8BlBPwmAhFxiZi3ZKk
qZxh8H1AGEb4ApDCjWB3WJrPtGaCX16WuO2SS+MvMd375xu8i/4yExs+wnHCOBiM0yJ/0SLAFr06
AkAamuDQsSRwSOGyXes/cgO3mwohgSIQwqnGAagcRXfYcVLewsQ2xiwtUgStK+3mM17/l5UJyMNd
kHBesc/OzMoNl3N6kWWIHOwDIobFpFxdgB+lrkIIV4J5FaP+MMlWO1u999URY6MLpHaYO4gsXFEu
q1zoikC4/GQgjKELjG0FTDIA0wXmgJQv1+WpH7VYh+J3ii1/PaTH6XJi7cTSloFBi5lPqf9x+cf2
9WPAgtHOpHVfOZu1+AYLVFa/GzNkm3BxyNf6oM3rXHcSkN40Am0YQTUgOfEBaSxOAfjbqMYK5MaE
C10J4PljOKKOEfpkkK50oInwGPeeOv9si0XDLVBr1NiADX0WNAPP5aYMKCWeIZQDPTv3tHig2IF6
mx2/xkeaKUSN/QbGXlmHTvrAiWs6HpdYgHmhLKStpBVqUgoE+YPUI0BW2qkSGyzofvMwPeOShW0H
Fp54jgVtl0p/FRK7OOOpw1rzJ4QC/6GhUbnZ517Xc0qT+0tSdsydgNieGCEfL821w+gSJeLdx70a
kUfQh3RFQo7F67l/Yn94JrkeflwRlB3pSEdx1M6FpEyOkJb8Cek3LwzVl4z1m/HOoC2L3RkWC/ma
WItVYNDMhm9qImZzll9gz+W8bO7KjMbwWAzF4FZ2+jUHJ8qE3jTiYL3QzHprH5c1jg+wJh2emjwM
XMp8KEImRblxNg6GJweAjq+FDl7cJ8jKtsiXwgsiRDmbHohYH1UxT3UYcZcl0idlhDizP47mOqNW
UsCDpiORc0GTSAC8hB07+H6q5UVZaqZmHFpdnddl8NX+OesHS/J9pqI3Wiu/kEUFS/AbLWzSqhc2
/aH3jfEyx34tRi1+zn4BwlvztnNXZTGiorZloxpPeKY6oxGE6/3Z52eZ6J6JDCM6jmqe2gsZBE80
Bt8kbTH1fU04pLjwoP+D7SEdRSNi3xdb0voCDkwj66S0XWQvXJZBmQX6U1KTYR8tIvTt5K+CCVze
K9Uge4m/EXtpBF62nP4OQD+6P+qxTIt06Q6ALZ7atpzufHQNPBe4Hmuyr9gjksewunNVz1CsL6S4
+AI2YXObjqVKn4TLSJ2Gog7VtvD/BjK+zb7JczbOnFJRq13xyvAKQ3I00LvW+rVuC5KSzWvEcN6Q
LdK++QtrICOTW9/tlJSsoDSATHHS6xiZGF2fP7bNAI1rSScylm6hH0FKVMRwTkwOlI4XFCL2hoAR
iDnVx3iSVrs5CWqwrLDs7aPoXuntSR75Gs2jIX+UvW8b2Azd74u4wu62UGMyWPZfBaRhB1HGZn88
u2lS0tXb5Yt00HYgKNfld8pxiBgrCMPho/JKIDsbaz5Bvb6gJOWq1Zfebfxz1kOrgDEDBNeiJzcG
yl7GfDAMBPYsoE1ylmQwjZe1gDfFgf9FFmbdys/8dGAk8VtOOPspal32MTaxewEdkYU3+gkRRzzf
Oky/tZxKKL5nIw3aUZb0wM2ETDQ4EDQbNWZjCzoS2uqjzIIRAXl48Pk13ZnS+8vbFoohiym+i45n
bpgir++MLONDcgItpWhXm3vAIaf+zU4bQNKgk2svVGzpT1EdZWn3R9dOv40ess8bmgoYsUx0JuNj
k+/1hBM3r4AsoWPdsb5WxZhl9DwLnvOIWdSt742yxauPfjbCjjLIJYke8/ybfVZ/U3BJ6xHTxG1Q
E1rdJkWLdLd5yoFGCNipSrq1RVAxIt6+p+K/Lz7j2gw7DPmubnMp6TyPHhy412yKH+07YIPd6Eim
HZVhBa87UoHwHRNU/34aRnUmzmcDMmuY6Eplo0tVs71A5eZhsANGeQnIsyYrHig+DNqb7DaHYZFo
j62xdN0Ont4HlfMqYh5/nFRTPif/L2Dl7pXG6Oake5sn+ngh2QuV2/lG4BdP4sRePZzAxyDwI+CL
U3LAweVm8dstFcZMYV/UI0FEbDDcpET3p7i2tnf+khXarkgOqMJhbHwurdc+580o8n9XnznWOqGw
If0Vy0RZ3ri4OUVO+ZYoBWbE3X9rVNMaVKo/siqyOe1Rkole2dit+o6ixv/aanRVZbBM3algiH7v
PBeIvXrKAF5r3aCvdFy3nSyBEYD9NlOH5dvyF96Rfwm+yhTuMBFGtyiOqNlfUwE+9Wj5Zf2rtX8B
9DcMTg9Xha1DtSnK81xsZ5S96vBduJZcs7YK7O9tDM815ZVw2KlHFUemUrSQRW72/eVNHAcNKUlk
UBISUl1UygmTmaQiESNbIK4wwvtj41ANYRTS3vPO18DtfIHI2k55z0Xa73Nfs6YYvslDBsw+xrgV
vSpz/X8nVp0PLH/CliDQmMX0M1p0aIkIU2pz+W9ztn8BYvaK3f0xaaFJWMgkyhlzTBZBU3xAmNiR
ehWKEhq2JAosKBNNs39oY3tIE+3E0PhP0/FyKwN1MXSmP7xWgW5dPd4HSOIKoUqQl0IPkgfKP0aa
o6aeebhRuEVuvUGn/wDfTmLBAffTVyIXdvhb7Fvts+SxUF7OtSq1vX6Bi08vOv1/K0YfoeLgMwaT
nQEXh8QBRCtUG18RMmlobMn2rI276ftqFcsXxdS2/Tuhxhla12ynPoHKQgtZyfpwMjn0Xt53d/Lq
K99NgtvssmMBWB7N6bp+kltxUURrM0uOjF5Eag1dQJPpP6KZwfj6+FZf0V9Ezltl4INTzWA/Wf/r
i9xYp+qtsLX5xQW3BS+Zz31eaJ19wBtSn+5C7rd3rm2R5thc/5iYhn3aKMjXj9agELlL9+he+0o1
ODrAyPH8NV4xehnFuyFSR1OW9rWKHFMZ6rUY/pxF1Pgvnb2UIbWU15OaqPMf7kQkzhi63UMmXBjo
5bdUOmczvCEordrqsRbl5uPhjLWmHbvOSbkPyg66LiZjYxXLFBRjTJD6xUs6XSnrl5Cjd7S46n35
ZUrFk3tV99hCKvOl0bq+edl6qSN/sW2jOyH29ZN18/Kzbtun4lxIjxpBzWePyxu4PMqlRm18q260
wVD6Yqiw9UvciapEPrhoiEy5OPnjbK8Z0VVG7dikL6c4Ihrnxf7pla7Z+LL+qfKuVtR5PhBkR+BU
Z263yMY7KHP07ZN865g4AsePYp5/NQSF/MaeWHVwuf4e8qJh7XTM+37uIX4wHic8LlYzdzHlNHQP
Ufx/6f6ByxrN28TdVzAI+vle+sBuONOp1fEcrAJA/kpbnbj/HlUtR8yVt3mlOEMQ+eZkCROjVAik
DJRlVs/1Sra5vE0sRaMIeR7fBp2JzPPL+vUMi+gpFeADIUG4WDNMxUggGTFLOUNFkvhVQOJc9hrc
BwrkZHZGbHJyYSrCGn4jt4zXCS2qLEmnb6G7xOiwo5Uq6uacBLTKPYTWmyoIYlgPtBX8Fxws54wQ
7EGf8Wh3vZIWRzDEWw0pfdLsLaIYvzfmReoZkCsu1Lt/dUUmRch7Naq8EprOJGR33LKHdW51s9b5
JLhML6eMh7wDrvAMPRGh494Cy5PYVT2zctedsPCoclaC0sh1HbIP5Vyedpy9923ifthUsVPRif5x
k2tqgAseq991H2twS+4lZhO/NJF6TiQxhmKWwY1e11EAWxGg4LFgpZbw/w68rcS5kLuDCYHPap1l
Mtg7fX89vyzaPp46dszwjZ+iAQe+C/KfEaRnKoFcOpHZ4JWHL0mbv7UTfYth7G2x6lIb7I6kvNGv
sc7DU3exQwPLgqJgzb9qjLfdbLtPlmE5TJfjV7fYahSkpp49JQxJigNWZdDUj8Vq1L70sWB7EroN
sTzuwV8d2qwkKB3MUYxhYusVSaue0ol4QkPML7bM3m4oht2dLrwPldy8VSVW22vVtSUXNcN3zwKJ
QpXI2k3tpie2XoZ+LfZvc68tXtDPbxkliKTRGqIkybNOt4YBAFwL2+66D4V3biiD3Gbh4b1ZBCZF
GYGDn8/xeTV+YUcZ63gJD/yYqQIQMUqWkzjsG+3kqjWKd/NrON5rjnmrbnM+PQGMSQJD0cnKDskE
xW6YvyqMj7F3XrFcPUOlM/xdjtdhl+2+SqUKuJ78YjL/tM+Dca3Qr3W1hvYJEGHExmSS6dZCpmJ9
xPvfCXlktrscB8pAEOWASGc/TX50TqyQza2jBzP0VRvzqLOj1sppYyWLKuQuXDAJnfs8XxgdWG51
wiDEC+/i49n22KCRsInOHLz2+T3HFT6fNG/Uuspb2d2Q21p2SNB0GGiT4Kg45KjdjP77MyVCx6uu
abmnz5KbAgMJ2Vets6zZwPbNI/XJv0dQKVw0BrxwuvuzUX1unC/HcVqHaccSLh65Xq0Ogk7IRq0j
g27/wpPbvQw+GXQ1jqRjZNagbB7LTynxJ9HoXHFnisvkvo1SgjLeEFnkRQNbsrACZyi6kBFOgLID
xwaUPC1ckY7XAF9844rm/1QYExBKNhqt1f2qGGPkVTLUy30IJU0XBl2NZa9rjQyfLxWPqD+RNs/G
ossMSgS/rpX3Y7lKTcIFpn3N4RcoaQIjTB+zgp96rsE0boh9zXXH3xYRP4wJAEqOoOu40ysMUefC
dyLZnwfN+kpL260yNnruyRNUvMatf3xA64CyaEp9/S60Ji/yCEdZaiyMdwLFXEjoVBUR11jkvz/+
y33fru2n4ckg8TPzhSLe3iOMtzmqSpLDjvhQOOv50jI2RrCgwWqQbAxtkwgUL5XGnyzktPzl5ZAF
RggQWUOUtf4NSV7Hy8wsoV2nrlNZ/9ckgCJuzsO4TYn1wi+TEoc4wfAvJHYJEod8MyHfilkexeju
NTetrL0sTg7Ykz4fIRikLBSR6D4CP1KVPbw8nUwW6Lt5GlFmzXS03YVmXGRjbYe2eDJI4IWvhyiy
DsL+MYP2WeF/RqUpwxB0Y9MQr07PGBrBFo3Md9xLsBTu3ry5OaVfeDzTSsBWgyZsOzLcRht3Ja8V
7tzBT4EhuT97qElezqBy2/HuLISpdNGpPIawVpvuf9KQXom0Np239wXYRChITeLlsTxrbSTMVGJO
Asjqt7it04AFcYycbYLHUYQV5I3l9N4YFfysIuUFZuW1oQEDfeyOfjoStNgV2ghSkelOd23YLJxg
vDw0YoWDPyDitiLmky5zDM+hnpXk25lbq47HSHLbUDURV9JFuCoMs/7VQJM3VhiKBDH05RlByxpP
C/jmA/m+9A4VkNaYeZVLC2mN4I19ezdtmFLR/EiHEHza92OCeorFAgSLzpUKr5EcVAcdBTmSfI61
P1CCor1vH2nrQ7fQdhBoUdx3mO9p1RhfIxGxA1pnKY9J+GBNzLMSqUILvZJT5zEl/BEzTQlW6Aml
C3thuPrJA76bnFy0GsutGWW+s3jyz8OJJaAwgQ44Wv43HHdVa/UygteGao82H3NzUiGC20tzXx2z
Y+sJTHjb7wbvlU7vKLu3MhL7vBHnx4M1T7/baQRjs8EyKD6ljDralH0Y0MSTu1whEA6nL01CwV4b
Tl3G2u69Dvm370IGLWGZoHIPtCmrES7exJPL6GiwFlrPiabXUOHw0f1ytwEmggP1uOyH3IPuh6jS
Jk2nOVo6KPiGiSplGz06Ca9zBGYTyCD5F5fkjhEAAX/6MHLovtzv6irU6X0BMHOwtZNjpLLH7aeU
MCmkTOsEs+vBNfhKtrAFs6EnimBYcKdWO9m3HtidETiPCRzBkzxrdJSzfHjA195pguszMVSn/CA7
VTidMXkGjBA2enqpyFliJHHWsxwDNb5CZjXpa+K+Vdnw0TzMnOkSaUuZJPJ0Uv+5iwKxIp3T/V6g
X79UywcuYJcKKH/f0BZBm9CKPtW1Gr7xef5b8jiC9jnbXhavdsmmMTcf2/nZA0gS1W2OOsLowBsw
CQJySWsP+rsJWCmwHwObfHNlJkmECAF2IGX74R0Zuq4YR4LfG/QEbqlKyap3VLLMnY6OkUgYZsJh
gDG00gOWh0mGMmYXRygsJZAgZRMeK7SMrWVMS50ew+tKfFpSD03Nr+1JufA9mY7lFFOdcguNU3Ob
eTXiskU/I6Z47noY6Vy8P520DnquZFQ8yK5/7ryOk9cfE+DB374hJN6SvCf3meRYicVuLdFKLWWc
6Z2SRNOxCaFHOpMq8UVZRwGZGrptajyWgnWlxVeHJ7j6l6clsLTw9kn6+FJg2IOsMQYty2kDi8JA
JQC6RYEApqe/9mxivSPInA1WPPnV1wfg+LH78ZIsakUIBLum3hN2EN+US+VlXWE6C2Q7zeA75+2V
jcRmNNzz5eDVw5EFEc+3k6e8j/T/XSG81xWdwpyZ/q/pSZUwbJS+BrryISzsWfRTR9/frIw4SWUl
Ki4WDypyay/tiwxeSp9Je/ydDCJfL9geaO7Sysm6hT7uvkwoHvbmqfPgUxp2GLalzZkLG6mWBorY
5xZh7wAAfJJcbDuTOQuv0LzoxoWJxav0lyg++Y6UO2wU+550y/Ga5xiL1KpAbjyYdLyZBhSo3OcP
jT/FUKRLeIaPF0MkfDIY+oBNNMVpOeCZzX49rTNbyOA5lfxGbfnsyTS5gNVUFfkZmgPeV2KnhilM
xdPq2obE8Ubplgx0Qq6Em36cCfBbdSwHJoeJvTy5Op0J0HxNqBUGBGEfwivKXHBqHVnN3PNBH7n7
s6deBKXA26sxpjQpzwl2G/5aZKIX1caUKSnODiHUVVEJiO5XX9czAtIRQMcbOyHXGmZA2o0qdesb
CrYklcuaE2nRKNznU6MJglIEBsZC7wpHm/cja60Kf50MYD5AVlzkwESbfVIbrk+EWUh5fevi8VHU
H+P2rEZd7Z6UW+XqBdOIskVIe3CEmskqJEQupasc5W1i64pnvVivcgdESfyjmerjMCI+6qVGiT+3
rux4EylQ+RPBM2MX8cdpVKik402hUkCSEAEFcZeuXFB+0u9wOfp3mJYyB02rfCj0rMvwo/XmKNNv
I0cdisyTRoEWGYqeQ7z5LDxd7QPtlu4fkjJxcF/T9McLIQLM+QdPTg+/pGwrJmFj4j8OxYrpn6j2
jDPAjEKYphwdmph3SHZKQ1cYFMNLfy3Ma4eZSqDqYW13N2HMKNLqdnqKyKG/DeweH7C8SxqhJUKg
tXZakpRdbIT5OEWMSQQEfT+AdJmpq6bzSlN1mSIXdFseiGCTj79exRKNRwSOgnrYFo/L6gO6bN2O
Iw7HiNjy1/2Xd+AGzAezAIf+/llTMPz3l4q6dKq0Ladd5mw34qR/SccfNsOevp0MsFXdQ9svIfk3
cVWEpX0fP5zp48z9hsRUmtqzwgEq9uFllwjk0nn1eFsMWGUquGHpuwZmUqHtq/j36isU9/jKaJpl
zFDpm7nA3S8HYPUoODKhms1MKHQv+rtKtT1pN1Pt53x2dY7XjDLyCAv5ieaLf6wWfJNCFI/j3cZ6
PANFDNixfmaP5Nccc9RBb5uF/TI/RGNDpjJtzzfwiJ3riGSDYcracZ9DKA4NasSelNOBxQV66glB
E8WsA3ka/FcnX1eJAmSUZytjy+d8N3N7V5dYqn3oW3cWz9BX2Up4puFJ0ZiqX1In7ZZfYK0xdoiV
ZRisDzOju9K+abUdZslSmAu98M53yH9k0yYR8mW5Vg5czkGWu3mX7bEYPS3mRFpUUsLO/1C/BDyT
UJD3pSd889Cdf2ef7h7yFKgFw9jbDZdX2SIeeHYbARfP6FnGzPb47rMU9rHFQ6UJ+T+q4351jcU1
zHeP5hq9WWbbPXglYwKtkVDrTeXiqu8uZkB1KgYlZpbGGpSKFcdTqnUC9+aegIA3Ejke4pGP9fr+
oxRnLEAgrFqqULb/GoBE5u9hZ3i6loieZLHeSkWT5N5Kk8SUKIfsqmZrlkQUliO7v9jTPueU6BEq
E6qLfUz8r+NX5tQWl9X+aQOYUHmuqvdQdzldhkAQA1xFAfaAFsFkOuUgV8t1xtv4Gc2b8p+Y3LmG
B79t1fz6PJWs527NbqxDXQh0TvEmOfZLT+gCTrEUPwZ57scA7LDma3xXUU7z644Shz1x9UfcEWq5
ffCL03vRw8nXAneO5bgxyCaGnB3dspVMVGb9IDx6xZtuqnj8g0/ZsKmlO8jYNEc7RUWe4SdPKkfn
Pu/dZ3+6J5H4Zyf/EO8sDH+mkfWGPYF2ShEpaHvxGP454mq9uNtIFHdAFymS4tiHT0LmlayCG5Ah
Pyjg5twBQ1PexIdMXfQQBqauw4sN5O43htlfygqsqh1P8Af8UeyM9g9wU5NFgUzZxc0eH4Z3CYj+
Gy89dkJo2IFNJjnI1TmUFq+jcIrX3KqqhHZpxp9kSZmyYK8aAT4coGnxbY6GQO9wgGUHvNVuZrW9
sUb1CRhuOlQX4+1OEg1RGaCS5miWclcw/vvoJJmRQCkVonZK/iNrPVoz8GwM0jJjLJWS24WzKlP+
pC78gsE7tvbPnBJD2Vta/xUP7XCNlYHbnmAdOYU5z23A6Bu0/CCwXTl017cHcIhw8tH//FkeozCe
AE0AWDcTKVgdGQxCWFBnVjrsO5AvhwLdbfDIHYW/5sUYOUu16DOKXf1z7XgiOD9RsnMjINs6RHo/
jUi1LOWY/yhSFYwe/XtEsDVmkhVsKWfAHQKG77F7C0ywBgkvIF5p17DdhEUaEKQpxrtUzTJQouT2
T8ugpKX4PJP4TL9A9nYOtj2+LrhrmQUEODwMd2KwrWsdTS2MMTlt2KvyIX/p/+xKOPFKW8ThIvUh
HBzkkXSOkeagHQjr5vceaTyf7Y89HV3csBs3Y96T+j+cQNmZWru3QddmFb+GvgNNDJDue+iOJBPR
i1GQmT2lErjpt4mWmFqD7x4b9/yJg5THTu8o27HecZ2gTYYFyfzYrJD+Tl/P6Xx3KO8HFylpi4tY
2gOcO4eR59no3jpdY337pARGOdIosZxwCPtJsEE/TPrTGcQVaj8rtZlfnqRYjD6USQf2ztIWd+W6
PsGZNExavqXEivpvxs0BdfQI8CDB2uOkeK5DPx95mGmf/w1RfE06L9yheFZqGhwYtIvUKZ1Y2AlB
6bD55ldPOnvxe8v5HynbWwrIoL2RdojHJ4xjolq6MtmGeb0GT8Nnh4x1RUk2eiTRl0nhsCZWoEHt
yXZRFDk+dcqy8Gd7fpvMNSo47lMwKQXiFA7nMwsAK3sGr16dJaDZdp0Qw+C3NJf18aSAMVqIrE3t
smEAtKj78QnlZEWmX4IokC3/QJRm2ltTHqA2cqM0EMKUEubJAnn7wnJFAeVItpnFvf/zLW0KAr4e
UJJ7FPU03n5hEnozcj0g3ofmcVZwFVCzmWx9K7LtAhvpbwAVmpxIpOCi63zgO0NMZKxSG4O+mm8f
kt07slWiBLd+eTc0CYVna1vFGYpb+3RoE9w54X0GT6CQwDxDq0X6wAkWjSstrTXukLmw7r6HH/Se
umoW2cDsQjR68dD5wCiZ/Cu0UizprqdFHtvGs2Lu4LVW1kbtE+MmpYzn9/4ZLSiK3GtgI+TI5iOY
22SKmAX90pG1qy22S0XOxEQrc/E2dSLaig+4GwtTq1RVeyvm6l94PLHRyCPVb7ESPc46FU0B7X7e
WzOrBFHTl7iEu+zlVE00C1NvuZ5cNfCOTkAH4VuWHbQFvb0ZnicikY9TSC+v6eq088huRuXG6z1v
UN1NsOVAcHxNbOpN0EXERji/dlJW0WK2ZuznG908HH6Iag6GiXKk0k+HMfhACgtkl2uP77b8gAUW
WrT8wASZtcKMxkjOTQu050o/mAmF7WhEA21vel5LET0TaFsYzB+nMRrfbmkunNJwHePPqDo+BhIa
ViC6//vpDDXTX2Vu4OjsP4pAarSIMlF6fUMNBQDtvddptb/QNT+RvLbL/V8NhcKHiaPNLF50l1yT
ilZFdlF5xIUDJw+cFGRLI8CNpz47E8p05aTB/uJbG9c0zpLKRr9Ew2a7Ks4qWSWH1DHfgviEyWKp
r5ZgrDNPAUr956/akSQIHPXUY4To9FMytZM8c7J0/Omn+Kw4GXsp0uMqHXxuOY2Z2VGA6YJkLWw0
D5zKZ3t06lwhyjmz4UcPEYWx2BsXrBMGO435/5E31COGG2xDShSLu/RjCkR0PxaAHsogAjDwU8za
SQAOiPI1C7FltbFBac7XZKl4CqDcPhf7UIfUkLb1MLXeiMfne1iGdBJWKzPPaZJvXRtDKlS80Ka6
j3GAMMYaq3BOeOR5IG/ByQ6xqPbUGeKhkmxBoLhJfdxjjgGsRUNN28tQoGRIPy5TFznnT3AkpX4i
idHU1aTEyqpb0887uHGKN8ChKiv7qKPb49oLg9Ar0hAf7FjzFX3OLtvJIPxj90pNMLgY589FX5Dz
7LSgD422LRbh4C/veMaHsGrSvGg7uHz/BAlyaBb1tRimMddw3BRFrAtJy9Fu95He1/qjIdv3vWgW
25A3Uy4IId9qASFGIZ+DbyUUQSyo2/6ByRMY5hqy6NtGgmxGm6JDTjSFlh9DpusRnyfjkyS1vl09
ibHMZHrvVJ2JA/vpTf5Gj34f1GJFRYN+r/k0hNQ6ztssYMJiHqzxgiXKMJejlba0u2Vz1ACpwFiL
ZMezW2vj7SfGeV7wdYGVwGJlngsZ+FinJ74sXNxeWZFYgAKJE1uWUEYYIY+AI1nHR1ie62ibz9v0
pLGOgN0sPeaghWnQZ0aBq8szg9TnXplO0fzqy21E5plNS+78C67OnO11bEYnFMrZnCvcsdh20hD+
nuePwQAxnlZQkfcclKUXatxTLdCnBIJ3rIJA61x7TNANgtcKX2Wk+rzmbMCuUwqNLBLFsca9Y/wk
97N3cYveHdakCb9pZdbPBTXD/I4VP9EeBc6ls+ayBc3g5j31lm1cwzGxSZWZu01zG+KKyqjVr1Yv
9fHNsllyYVJg9JR33iqOEYOCfuFqhfBmh4R2Qmn4ij7p782kHLHxHSkKnMnHqBmYcOTKDF3QUjRl
u6Rz4TWswgTzBFP3785TYEjiwQDZO8gwBMMGmWIhGr8BzKR7vE4OgVK4fL1yZHErHqml5opw56Ud
yCB57LKqXYpr3bxWi9lcYvawTFp7KwirAOVe4GeH3g7T2HYkTN41Rr+0yxLRurHMRpJY44Oo3LTu
anoIR37Zf8x5l+pjb2Wg3aBQ9fHNhVeSaZt3n9NpB6a0cn+2msQ5EVNfBPXKoZTt3XrazAL/0LaI
FnKOtrhctAuewAg1vquLfIawAH/gp0G3oqCZmaq5NEM/X54Pm7OtcG0IWTqt/QHLGQuiZyceiwDT
Ngtn0Z5yzevKvKt6WEXuw2daJlY+vRLsKfUgqZrsM+pJHopns03f962G6QPfTTPsgalNrFTS2GWQ
gW1703mEJ2Uc8BqE4bhKKew5mTJWmPEWonU2Cbxd/GeDEI0loqHxw/9L9y/1javRhkD4kA24uPfe
Mlu1JL2EOir01XrVTh5qKfY+FbmECsuXMl01rLjFoG6OlACZcPKWnCnnKYo4fEhX3IRI8W9QXkhm
dqLcVsvf34fsEISmY4TAM0YCk/zLQsbRuNV5hDcQlKYRYVNaZMu1PIvlaYMvpjJ5VusXTbt/vfBg
BESnTrRTGOnMRjqrVY+GFOXvqGDtzbV8yjBLeczFO/yD8KxG0zSMRJ+mlqodpRuhH+NVy0XsIxy+
LHU05h8WIhQ9lHkHwRKdT+/b1fcZl2txyu6j1x4HUC8V6i00FDOH3gljqQJZjM6PPpwCAqjioICg
Ocn1vKrq4w9hxe8AlpmEWWNKio2wyFe+VxgROMT9WfXvuS/LKtqgx+IWvqLs9EADaMAvuX91OPgq
Ey6Ov4f90KnqZ0YTSYiiaO2QMDSQuZVPRsovJTJRdNTTnJXJWTqC0qXLWA0cab+kKmg3dXPEbb/I
UjCbyAPTMMgWjbn/70bUUwLJuhDQqOqhWs2GWLwxpUlX1GIm5yvaI4xWLUBl0UvcHO/16VIDBzrJ
aW4NpdXJgqJS70Vb+uQOBPPqouLippv4abMrdrHCDIGSH1PaAiiHSjoAIu8i85BJwt6ULY48Htmd
J8VW1TAx5WV77UtcBra+eMnl2YzjCdfSqNYHrMa8N7pIBD7TItludtXIzJ24rQjUgHurDfj4a2VZ
3kh/fFQuAgauHlHDkIMLTSAThsr9UCx6KBcjQRjGSXZ9ZG/tydVlVhZz9p8Is16Jx5nT7KjfMAhB
hcImCJL22YqGR3VLUyrRq6MNhgzhgDZczLNY7tDz+hchyMlxjM/98qPsaHmCN5a26ccGuRXNgzVA
qnuUNn8n4EKdO0k7LU6V7JvUJ2eiAkZTZ4UengavOhgXU3KBLaeGZ0gELDFrQIs/pL0K3oNjGF7V
qfiU2wHKHHNl6pLdn/S8BhML80s2Y5Q4ceRfylZxblAEDtXoeQQxs2DJkD6AA5xxrbOS7JaNN3rf
95tOR1/yb8xp7h2CAtqBhYtfirwqKG5aKsDJyn1L204fUZp6dUPlkWm3/nXnMIMolzE2gHMcQHfj
VBGrPLB+aCnDoVX7CHD//SrRZhzgy9+1ls34TC/CENTOv8We+v/2siM4nj9chzCvvs0Re5X4Cn9r
/4vVIz9UWH4vXANqUGq0rXINXiRNxL3PxVH6WfF+Jks/SAhMz4mzGr76qcfjTf02pDeZqWGoV5fY
n8EIADiJZQ14vM6Iks2pYKIlhmv2P2yHKVM3vGxsxLFKfCZN4gpYwLjGN3B2Tnh+KR1h8CipU8Im
8uqitloaPZgtACIODsSfD3wjqCBP6Q4a970KVeKqY4/TEi6CH+/16+LfoiuSCwntdlR7Io5f3A9K
ItvkvzFL4cGnd5FB0h3kopetTw8riWHBG7pY7CinNA1o4wCDqPhhM4EbiDi62ByCP4YhttIlX66j
Q6XSPj3NSSekOafhthERhnd0wHlFeegmJq4AkuZyVzjMpfhZjhpztD2BhC4ZnK1QwndTdmcN2+GW
cluCKqG9mWBjb0FzXRJVnBq4DQxmdRW98+Fwp9naf3c5UKcyQyUKZWleQT9/SW+JU26p/R+4vifR
HXP8omj/BNdnqHtbz8JirdFjrBJQgrYrzOln4P4jAktjRS67vMXo0ObY6bIcC2FhKxVrEwxu16Th
60ZoqGmuCBKxcjhUkHDRTql5s1SJ8wgBKIZnDcMJ/GeSyr/uAABLTKk71QbsBs5gFeMH/gDTJWcw
utnF5g5K9G8sIHOc2BH9nyQb98NWvLBdBkmYE2His50PaLjkHwUZGm2DrD8ukv73mcVF3jbSsSsk
wbCVmNuOJQynaZK4EgNRdMptEPiNJHbyxKFCvWE9GXl8Lh0RbKI7dCtUTKIIodfHyLNFMjl99jBt
MBE4Hvo9eHmahLnnffJauaT0U8ZLKZcs99spOmL9Lzbz6D5Kr5JmuqrViaYqr9W3IrsZB/TF+Vbr
DxtW1p76x6/MmiOj9LQe86aWTBZteAXmbJsrb8cyFc2lIezksEYK5IOLYco+D7aLvlCjcx2N1Qp+
W4Npf+C0GIdq95fdlO8otbIoyzsZcnWXhodXyDJBMlY+4GZPbIBiOYv/D9SqBdm+TtaXuGu7WgPt
eDy7lpmqXhqGlLJdRg/XgQRi8yLGRrwS7welreFF2Mkl1ZUJLUR5100DeH9oALu6RXrkadlf8Kyt
AfGvu/ihBz+uwz2UF7gXKJz5n0VmZaa7guGqr5/C1PthAjsa7C0fV4dCjPKrVlE4/qulJJOL0JdL
dw+peXciPu1nr3njs9vT3Y1Ipleqj8ET+OzsH+KvDZlFYYZP1f4Q3hNJJAF6y7fyRg+gKeea0J3K
4P6jLQqUsdcr0AIQEbJY5mDB25qFRQG1OZkKrP/sI8N6Xzq1OVBI7UxdfpAZ07Bj8K+qVw/aA+Pm
o3V76JNHvDi24fnj1Q2uPXD7zO7KAfk55m6XDfodhwWHhF7gskZfJvKDU/Id3I4dhccawhhuOBbi
0oBAQvfYvRawVCgrBya7N0n0pvoGPYSiB5bi+/l5m5TfQpSzki4VvDEkYrLG4Is5D+yAmKQNtqzD
bfKWHGNIOMylZIubEPpa6UvM2NmSi3Umvg9vezRgA2edD9B9adDn++0f58TNkutqCuLyrIGF/pE4
9RC/XUYXHt+4RxbOhXzvgNXrfKJkvVFG+2m6TkbfBdszzXDhmVfUa/SqBcYb60SvoTp97PJxQKi5
UKC1GXpc5wJFZuP6slyjcgFnPOdd5dzw6275uNFMYOxASEqe+FEKuo0ciW1hQMjHg/+vd4Ay/Os7
zRdIS+AwD9ESnjQ4bQIWi8z+lS08lML3GubSE/CC99V9gZEyxePr3EiS23CcFRI5irhPye9rmfoo
huDuDFZ1Jdav2RLS2eHhMX2kOOw6zC2HSB+iiIcXRAsyPjzQznaElaQFtGGhC38/zV+j4OenDVZX
bqsS7iQh2nNv7d43RwJz1eo2cZ1Yt0My+paA3Ov9wJ4WGV0yvHv8Hcqpp2qW4hq727qAmaBaVVNC
RgOw2NrvuYAZaLPHKK2RkIOITQPoXTucpSxOBJCft2dXsyPnUQ6VPNwRJ5JSJrrVKQX28lyto/6N
wKrMSYwAKVwxi6HpRnnAwiWkvRhSqfYJwxvPpBgGix2YGq8RW0+L8oWnopnW3xGNlK12vVdWWZs0
VKaR36DK+oCY0d1WaoueyjGuPuquAigeOgzs5X2LyI76FMsSTtwjwjum2JmxTC0IV0PgpHhOOhcm
FkC3gJSXQlrAJZvrFbsks8Ti4jLEG3sKeeWEtW+DLD5JhaxPShZLtBKvTWy9exc8eEkcDxx4du3n
lwqrZ/5wokHkd4jaEKKvqcvFQnIegDLLvy6o+DPI+1ZDTsdW82ipxBtsePWaPdMuGjh8i4onYAYa
saWBznsveyrrUAjbQKUK1BdIcVm8StHOcMvPt4qMkRLOh1BObS2zSA6B8v3Z/yRKTfP2lxxEx7go
NsMnHSACsT7VlNUQBFZNKyFNqFKOhhKquMYEhIv+GKfW4utNP0dZhN8PB4bZKxX5OCLrYGm45xSY
NQkDTC/fjtIQNv7AtN/X7d2s5RceZnoOVOVyFAjnub4h8BsxULJYcTfsp62KnKjm0cCeshOyEvE6
WETCbDrItfiaRP+aWMNngAM/N/X60a5XwXn/zoYyRv7MaB0Re2MeRxVSFqOuaxShrSx5d3uzX4FU
u8aIsfRFToHZI8bN8Sax1H7Cg5ch62Ml7amqzzHo1T3Mgy5AcFtfrVwIfMbHKeFWOXj73EiSFoyl
PM2jsaT/tP405l9H9j7tbdJAWFrZ+jTdvFZY/B2LPS5r0BQfNbsHOfqJV5Q5ICkM7wx0deNnuYiq
OU6uyrcswRT7pUvUG3UeadPsZZjYKpMXLqEH6+Kcuxnac75mhZhz/Ial86n4kAVn9CmL2L7CcNtX
so+tB0a7NlCL4KUUb4A+w/7IdJEeIbnMAX4AN/BTFLV0917VfPHqA57Q/FeYA2GxQNUAefdyeg15
XUaTcnVSd4gomem1uny886futEqCKB7Uu/hmylCSrCqGXJ3KA3FLq58o5AVrebmwQaZrKutC0wUi
JfvfUKP5NeW/WYVmVZdVL3GMJFFG7jGrtZYfqAbgK8Tmsuc/E+hJAZvd/0+yOoX52Y2lL4ZYVNoq
z5vBhrHFEaMGVcxuxfJymXQbaWdh32LQ+g5BNoEP/Flnhflrz+0RceX4W0mAPiBuB8vHIsXt3sle
0EsAK2tvhmbDrGMvl0G8P1PAiefxc5RVhyIjxNbjGbXZUfD8QTDiKXf5FwL2xIeoQSVYNDF6KEJm
g4hYUYuLPSeQ+j4hF8TS+03MjhFczJF0kcgbdYb1iVCbg3ili1/4QkpoZv1zOySxQ9nAIGfHvUXQ
84cEgsHm9LO6vvJNHqHYmvXF4eaavDoc+oXXWuk6OY0t6H11MlnpXctWdfBm3p1d+4Wf7wxmu9kC
ODV0sqU+qbZeAc1W5hZRoQLAyX6HhZeO5OL1O+wklIOQx+5JqfnsPYFsagAgHoCBRmHZU9NGGVc7
w5elyxG6IWoBZAMJg0zgnb2qq2tsZDcubQSsqYLvCm1bZ5aDho4UJZZuQVMFD9RxWoFkzxuzxb34
V75g99848w2lKivEzqymcdhZorChruMS8ZvEdB/kM60qaXseJZIopCKctKn2YIH7PxcBjVtwkf1a
Qdinp8BJqJ7ihFX2ONqSPjpeNF3onZiRRFH3IE11C3wZ2XDRDrXJEhVOAWoy7J7iGADiPe+bQ4P0
3GW9PjbPfLFm4BE0kco13tOhTiUkqedU69hAFnNGsZUgProisVqrNMPwWqyv3piT9V1DwAFejH/H
+tpu2JvkLk9VHeQZFnVTJGvs7jX7Gov75FKo3x94nD/IGpX+FLv6WEobso1YYpc+6jA+GA3yozuh
6XF9v9YprrJv5RxhIht5jv8vq0XyE0sXyu7mzcZR0PWAmk4MIVqKAK3l9Q3W91fGrnCRaynfHIgo
axuFr0r78ffeibuDKhxgxynbIa67rQvolgWZx1c4Ixk85uT288EwGaEXmjjikMr/i7kpfPZOCKqM
5zddmNBYpoNS03nPvpAvHt/c3tngc5w8P7iyPNkKOCVlddi8opZMFlZIywZC3xcw0A+Jl/KpI40C
cpq8GezsVwFjEw8b3l4lxutUi+GEBNdu5sMa/PkxMymIin+KtGQR21pqaE15aP/KEBWhUwBrnsIX
vnuMFsr78BPLpuZVXENy1inzcqgsxWJOFom8nuSRwRDcQlgDeAwjWwAYFjWX8pG4RIBizh4gNj/R
ZTOqZHQwsFgCmH4dxOUeNjlCgDdKBteXKPptMCIpKpzJlPX70FAwsUMYo20jth7CJwg7tW2s8TZD
icbIM3g4jvwFYqsj/gJs/xK82SJC+duzKZEO3jfWmaOrAEyeeuT8ZENNOl+73/FEHhbHaVYu4jm1
MoFOZqdXUPI7FdVF/4rsrRhzi1bZQd4JAi1D/JavIRzp7FwoqhFW3qdTnAsM11PR+UomVtK5u2gI
oJZRta+/TlyD5AjI7bLUwBlLCrjcaALtmL92Nfyw1cIpe1RxjamNG2sE+myhlIs3MC5BEmrWgE8l
BIo06VbLp7f9GfaREAxPJOGNBg2mKjqr1YPOzhuJymXlPh1V3yPKjDO41iBr8Mz1BWB0rAECCU3d
mHjmBwMmxexopWyugSeSflKqW+fNw+n08VpuwnWPq/YwnyaqSW1ipo9Ar1wsHCN0fXK9DxPSdIer
tOp27UXHSVpGbjiyGwAR1CSpFilJQXmWiTQszeNNg07BZjv+iaGgpw/fh2SAtWTN3/+OXlAMt2JY
fgJNhc/WhJcxY1bXOPGyJqnyGDPPxclOoCMzrgvHRFWfKOL7FGwRlB9c/Y7efqEbLfLBUFZz9/3B
RQBqMBJYYhFumkySi+EYFsjRKavevkZ0pNDMwwBDmUI3AOCBZvMD7J+TJfPbVAMwvQSV55cPPxJZ
xId5NUtuNqm9XtcrW/7S7roxXMCLmCG7MFWlS+BS8U+lXNnQkNY7pNy3Jj69hpVreqRUoIH/YGix
jKvtV6jGfOcqyECSZAgcd/asWYom6T0+2d4FCoBerYglsSP1rfFtmJKG9kYl0UW1rWolrukb/vpQ
Q5UE9MAOhD+yTSwXDwj9Kzn7tp2LAE+ycGS3CBlZgEMiGNctgMHtTWuxtPVSxKK058+WsCQi33kb
K9BV28mIkzj/oo+6Ckl34GktIOvOeSityXYOzVCmoJVppWo5Yki7DNHiJQbHYjKW/iatvN2vBuGb
7wVInd4b2e27JgQFj4g5DCd2Yiet+RTR3jzRIvYowS9SR5fVCPVdk0UaSCc8SdaEjY0x7KPBK2zC
6UwakID2/tefr5HTM0bnHeXexziGKaaaP9LhrAHjqrYRluq++SrZU2R7bN4RaiMd3NN4ecklBSPb
l8IiDwQ5FcM+p2JruVeGbX/E3HWot1Ebgv4sVDmsy7sIi71JnEKqBZBxPQCJP9YPyIoCbHy5Nh/M
VY5yB0KpXzG9VmZAOkhx3hXQPwVwyeiCiXZETR5ljPHTdp1zdDVpXjKepnJQUMaMJzIVeXIcamXG
JX7p9nRRq1XFus6VI6Rbqkw3JJ70KCmKvnIQxjQ9uzBvzWiaWbe4dM43bz9mQ2JLTxJ0NVFr6RzS
PaglU7Mcy7rECpcnG9JNGJNirlU9nvo/SI7nVS7BLsGM03qKCfRkU+RL2vjNDurqwHnDHofXMQj9
8HYOhVqZ8D9pIfkvj3EFbIlNFwlNcOeHW4Ii7MNT5W7sSmU+pVoHbex6A4oHWWQ7XCCT/Eywa0P5
p4EUi4A+UDkir9Ly9PFAe1MWjxVEg6ZNmtVTMcWPyjjIlWyfdocyQlaJWt0eRofQL77Qsz/JPZYd
ac+TfL6w+tuJNd/rperCMVm7/FhGVU6XSPbqM7fKCtLL84sjk/+wTdBMu/7xaWUH7Tqsn62aVpf5
U8d2RRw6n2M+MMYlCsK5uHmAQfO9wrNF+z72hG9PlMyLz6kxB220cFZrxV7yI5dgLvAbtX2fDLc0
TBNGNbanwBeaefx1BEEoZG5zY30RkaRmqG6zUwand407fgGuE7axOvnuz6uHsHbBG+8vcW7V9oGX
Sl0EcssMbs+ohQdxzlRTDhJoN/o6SGhLS1y8wAIork9JXX1/LtpWD5un7m7vU+eMHuq3Dn7PghiB
AYUHa29xOXsPeayknK6StYHmY8/Q0InK2yQeFi/GCZWYDMG97ooIgBK+UmexxxXOJob2qfRGvMLL
0Gg28GjG6QUiyX4gzENcyi71os3Z1oa0ugHJIl4aASX4skllmmxXUjmT8OCaWF14NfnHRqUiJ7jl
BRB1iM/Hu3hzL1Xm480uj9ensQJDcyxCva9ETqr3VbxDpKLBRVF+mOWP1nULWs6T5tFkS6KzFjGv
Vp3bOi6YZTL7JVBt/lJUQWJeYXJWYhqMTQ3dXJMpi6e2MZpiKrufHVDZYgKZcRC6KIPbtv5l9iQw
gxDTpfw3lbBqXQhtQXDzShedNd4wxd0bXM8qSqUM74V5RfjlzhFgxkVcS0JvMbQdwpvswCZMIHxF
aBwfgDmexFUmgKxiGDVEC7c/8EJGwzrWUFe4j0wKLE7pm8p1iw3A1nw6duJxHNVih1c4PaK5vZrY
iBnnpJUbXDVtXs8Z8mrnkIXgbjr8rQ3exj9Q+m++hAOZXMvVRoV3EMyuN3V8+kcmuIkAYwraByhA
AIEivfr0DbNkQx7/dYtcE4uABNs2eUMGoz/lOs7OslWkOzIsrs5kfFCYDoGpYvZvywzg1wyZgCwz
phwiU1A5gFC4d+B+eYyr2EVxRKVSTgZwEdBcs79rDyL7eAAl5d8ZB9WL5zDVo5GsFjF1J+i00amg
+Bsb/iymHoL0JURWw4BCgtZOsSmCS5DKN4KRSUfHK7SFJ7BGhLNtQpKbdRabvGuKr4WnmsN3cvuO
cSc1bvrrWc0LawUINxi2/q1VGr5MmQmusOKX+SxsK+95xYyMu8HOQz+flelSFR0uJX3D0eblG47e
qF/3T8sYRJxRv0iL6UYWoKaxK3lNj6zgBrwpDk5A1LgDeWqFrRtnPCoTj8RqD+e/xADGenbi3H6n
EeYopsTX9WgQlYch8l6CLThBaG3aVrwYV1r8mLVk3o7FJYQ3u5i4J3wK2taPruozFsn/dHwHV1BK
ReNxkjUs6rdvC3Nz20+OBXrR4ebgCzdk/x16hmPSVN8szBgLhyATu36dJ0NowKNZKYeWXJBrowTT
PIJF/VIyKs43cxOYrl3PLloq6o7L7h7je60ehCt0UuEALgP7SZ2zTqUsojMKXt3tDxZWx31r8I8E
5ld91lfhVE1HKNf4ZaPE3F/dv3JbfYlaAPg+G5TKA2i9rkNpLzchfGgklU2cwwOhmGr++r4ZdThU
NOh9yPAvx/VyD/2r5RR/McSWKai6E9S8ol9BKgF1dHg6QxWcrG6GKRWqrt6TE5kAevqFa0e2Z+gQ
HD80UgK6YAojRJqqLwuwU4gChZQqhxqmqQIkg6jees1TUw10BoLTvvA5WArlyhI1WIOitWqjl7Ea
5+qQwsvJxKTqccoXgRgXSx/VAP+FdF0rbxgQEisRrR9Q3c73q6L5LJGp9GcveZdqJzW0NaPGLPcs
vb/LoV7WlM/DHQy0NpKnrBEOBgatzbv403G+sOixf3IigUZckqIb863M1+gF/K4NzVQEhx6M13kS
al6Rt1zdVAAHwGKLJIPDmi8XvSDY/7AUXtP8nC6Wckm6ScvrJENd3Ns/HuuFWbQ8GP3XQdCwhy+v
FfTF4z/CuyJhKqR95kZefI6uOkl0PAxpY2+ZGO8p+FyHd3/0oCZzChO+qvqSCjArwjeHHRtB7MY6
j3M5dRulSjjJ0HU9y6d9WD99rn8LmotEdHmqrLokGMinQGC3nN4kpLV0hc/YyTeWa46kWI2BZqRo
02AyiDv/9QSZuYxYWZXngCwjjnAg/LoZGr18YyJIg0zaHoz4x+cYrHe+kSy3ruHSE9rH0yXj0Wql
uUfwTJxAsWl/l5T1DuqdVuIGMDCHYlMP5xvKXiM+aN7amj5P5uKzuIFkTJ5pnPaRm3agesQGRzn2
F0Bn7NqiAdFxlLn7DAtzIL2OYHbi+wRXELriSEPl31JRGF8L3UWPMZxb5fm2wB3I5G40oxm1KhSa
F6DfHUFjbuXKeOMvODYmCw24jhW9qAAVRi30e31G5IXpsLrErH/jNe/tV5693LLjcTJr93hNveRd
vATFkeI8ByJhxbAaQwXaim5i/QhS9L/CLT9O9QPEiPCCBQoTKtEToB0n5/G9KZCLUCmGzv4sr1cC
4gNBFu9rfOg0oxNjMqK/tnFya04a4k5zFIQkcTjKikc6u/4uQJvVbIR73o5IwNwHdWkj0QjwB5pv
e84+lcxZ6ps7PnatoOk8gLmPcLCL9Hqhw2EPGIHmKkYBqopSyyGZizAUVHhM8x66HibVcvz2WiaM
CY2QY37JdYmK5tZ+Of0KL1v/9PC81UKV0iuiNaO3KlrdWqk8inzMxAnjGVtfgAnA+nTK9e1qKtnh
w28/fhox7KVPpLrJ8i/t3tayvFNIQtlCT5kCASE6kU6lawy0xzIOgKxVWDoEgkFInuqWzeYXwQG/
n7daW9NlIS/S5XRFU/zRfbdB+ByO/USkCfHm+NPMoCs8kvi00nm6fFWAfsTntpdKC5I8ndPy3oCE
BeggP00IT6RX81u3CPIOSZN5jzXcCoYiZTz6svmykRECT016OcGtdILz5ByOn/BkcN+h4WY9n/uZ
F7MVArecpkb3rI7JC6kecLqI8SZ9Sej/2lH5qTZUFCFfbbwqslTICosQcE74dnELQ8Du+aXdLA1Q
eGRY8HhAe43Ymkpr3Hq/yuq5jFK+2Z9MxeiVpCANsM0GsAlG/d9Wu3ty4z9flTK9EIJRLV9ysHKS
Mlgdk1bbaPZkTNAi5/Wy+5893DqjdraG2xjCnjVRuHT6OK5iSl/8gRz9mZydBFJLYAZxDNPK6gah
ao+LRKDqjHzWL66Iv1/fdZzg29cFnOVnE5rX8exM1f5kQ7HZJqFhubXj1ieR7VYlVvM6kFKW6pKO
Cyqy/PqiwBDqRpjT9vgTMVI020SjJU8Y5O2dkp0ee0ARWnY2foQ03Rmuf/Cd/imPnsGgSnFoVu9J
8Q20KMuLWcWmsbJG2/jWWKQH3Dijz04W8y0uv3ft3MiudQrC4uT/ipqAv4/X73/H7/uKe7xHe6sZ
tVi+VBB4AVxm/VhIRsfxV80h+JyNJ1e1KbQcOK88cqF9aFLBKffqRAes9mdqGTGRS+6lBJ1Ko6eD
kREhyQWMwWfWIA0wqt4yOJcK4HXkzqyMtfeDrCsVPsnsd+1x5fjBQS1uFnMptpA4/vdnEMGot84m
7fqyV0UDMQ3BbzUWnCCdR1sklyI2Vd/h6atYKD1j2k2ZVukyNW2i22aLpOVHbMyC3yWHJpYzeBET
n4+zrxxuIJ24QvfMBU85QS2Q7w7RvT7p++0hgoYYSQtRAdrrSckQUmkHEwZUsoCu9QvopCYzRbOc
oMIjN2LyMo9fElUg9vRYD6R2OymBIzAVXj5sxygsWW35bwxZIrHull64BQGM+OAYtBEW4I7b/R4u
rXkhGFQf0m0ToixU3NTtXwT+VX/iP3xJQo0NNN+ldId7Pp8e8EQ5JvUHLQFGhbQ7pf8WsW5rYrAx
HyvpYjE1i+qEehVDx051b0UnslYlsrDrNUBZMKTP3sU6S88goPkvLhjvOqPI9t/J+wRk5Jf/M5ct
+NLX4K8U/xUHKBlybXLpqguovX35sELZN2lqqKYf6dmPiflnVgr9VadL6HQvlvASt+aBB3Ts7rzA
sPCFeonCqUJyyiJasqg6m5Po4Y1PAVm2iPzy+h+rL6LbuxBicEKCcSHGRK+uwJAtjRUszW5S2ilS
uUCt8pjti1XPr10gF88VefCYUIvOprIj7XonsBCOsfkY5Vl9mksqVs5HxPKRBOzFtG4J0jz0pO0F
2EFpWMiXis3uOjf1XJLfHv6kLeqTfeUvSrN5qBzp8VDtob+iLOwlolaUYyTTnTWZscusn0Y7CgPE
2KiTgLBkEiLcUQq8Lw8l6P8xPdEw208R0jakdU5DPXDWRe+4bwsGdgjbrN4Kct37d267KjV6DbY4
ERZ9xMFR8A/PxbKr0Pf5ynSCxb41gy3wMRaa9cKNQ9HiduNNJqCBdyDf628TtKD2sxqdViktjiBj
l3eyuZGLrprZbrfuCODVBHIExvy3+5CTLRqWM0O/DT2NmqmH7F9j8xELwjayKOphtEbaPV2wdmay
hk660BRKvLlsG3/2HBId/j2LydmUXdXb4O11YQ40/6LZrcadt4FXzKsa7ahz8MCow1/2dFherTCw
xea/HG+zyEXOlR+X/YUJ7jx9mV5UAX7zC4NNB1Q1QrW3lQ8bNXxsA7kHWmFW/RqMu1cGgUX5wCVa
OkznU0ZP+sEFZLwcKv93YMeTKbgWO8Fe27koUDEg8YCNxJj4BhdFs0S38eBBWdIunRuxSYCpdxk3
Sax2eZHwap6goMmsXehMRkxJXrQdmyu95BaVfM8gnCQTdyCNSgtK/wKrSNKB6gtoDrtU/bZ+HYDE
Sf3EWK9KR4yGcKMlpSelhciLmBa8IUbvSnkSDZX6npuxX2K19t6WSHnkwYDYOWbIPLW1wnxMHiVi
/R16qI1KrCF7g3JV7uWubUp2S+O++Dp8ahT8zwkXWSWsFhYAGPV4ZweGJq5YO5QUqEhcsurGWUpE
w0/kZtZN4qlI1s7/jaXKfbEvmehqzyDra+tn7doJfFFJzkEzfg0rDbpHfPOOjXxLBnSriWPeAvcP
CiyZBy98PD54mzR1TsQFFGqWHxHx9UvsQ6gvndc+qVX1saSiGvOIooMCvv1qGqe8BSFusXU3GcWt
GI74pYoAobjwzx5j0V2SIBem/wDdJZ2NEMaOKc8BdccsqlSOnHjtyh8lNCbUGcxqPNlkl28eGGqK
2O106eAu9o1E0TMVgXz68QFCSyvb9n6z/h3qkI2sotdDeXcczZKpcuCqOL9Ns0AHg+fww/UBneBd
+C4WJ1ey5Ebbv1hV72Dihd5dEQZpGH1NUusWGxnoWWHa/yCTRlCmqE7krPapYHgjt50DjPJ/vzaJ
DnnU2jReLzR1CTEzCykiBBkfwrFUPv3OISjo0Gvo9CC3ApPSAsf4q09UG82qbUWw/s4SIZxJOQlC
pVxZ1vwDvZpaiu4IYBu4Ke/ePWo7MYyC8ouhpWBDwtlHGlT+DAdTAalhVcU3GZ1NHpH63y4xXSkk
Rb1x/wQkWcSkxO2U1l5ERC6/kFl0bBIYOynCtUkCvtHmCp1HY77Vtjgi14PCjgvUt37fYrLfF+E7
hiJGo2CKzV7I/BKPEnQm0ULJFiz7RXoUwO1hlE3tGnDgbe1OsiS9GXTS7Y+XSkHsQLRB6kLA4K1d
diMpLX3TOU+cfNdAj3iHI4O0UjalwQBo/jN2ipat4eLFYxjf0Wfgo+VoSHf2yNXLeA+pCUagclR4
AX/ugyBKLrmd0yzEOsHLoh/8aG86AMmL5qxswlcYH1a9j5K0dcv/cSCj31DIkcbX66djhbPP1zGa
kEDoPWaX7TFeROJZmywGOPUBfAu6mPypiaj/l8Jra16GiUA1Jz9LZadKPZbZeUTtO67JHlLhELhW
aZ7VKVDAePG0GK07OMjB5neYP7j+dYt+5PwkJEMC9twfSvCYwGUG3sC1MTzkJGGTVKMBZAYgdgw4
eyZa2+vasLV7rElSYhklB926H+dGer5EfPRpX5g/vJJh3ukiF2kEzphl7iEAHptDoRw4hIFaezEm
iRifdZYbryqWVVnWIE9j/vJMch9oDFZFhZtuYB0Up7KyIzC+K7CqCMo8ZEuiny8C9rUiYr6fmkgI
ok6fKOHHgswR6sBz47MAj9xgqml98t+lTgjzEKY8+oEW5NSZW2LK3S2VTq+LvmtTT+MC7O8dZ0kS
aoE5sGSCUUL3DhbfWB7+Ohpv2CAwNtaIXk9qQ4xtCp0P1Nqh1hCu/52DUK7goVFcQBZ/UAr9aQY0
C4Q/M5jM5J+mIROMnScnspRDnDGXYpb9kJhG0Y8AmGhTlbWy5DNWBMnXcBfA0xr6YTyJjiVBcswv
Mk/YkImLRYqmaUxyD67eXMjFJASo+Puf9vQZC4gaPje7XX5iBC+E/tSG6KiYKUy2oVxi9uJL8xkc
8xuPGad6Ab82Aj0gbQ/5TInQ3F2BbF2FBuhp8KMqXwdfDAXl8PcwrcpDvg32Dq+2eOhzoZBtjmfC
N25va6BdY2VSSHNnI+a5BJUUIIx1P1PPcxklK6EyBUaloPtCw/N97L6oAf3Fwvt9UzA0hOe4XD5J
t4GX3IpKoKyGm57gSfJ6z1B3MZfSrW3ycvRdhB8W/L+5S6waSQJAzUPw3hORTjsaUxgDtqcfdTox
622M6UI5CjGMYetZrnB+JIO9sA0V8uYuwNbAGGOdhzTHsLKgcSBYnGfuzIzPKque9hW0HbC12CmV
OAJLVjSn8tlOB7DRoCq/9Fd7WwphCGyd1UiN3DyNCp2vVAGYsuuJGQfCjy5ogxPIpxuTlQWzOMOx
LxdP+kMViPynD+5xbpo+KdSnZ2EunRVAnR4YcHKZ3Sf3nPuc5q8XqNnn60FN/pVFQuhOh19ekADt
ukmO34RK7qtenmAabTCg9HMHL0SIU0RH7BarlftEkkkc1UXOFxUf3bl5T7T0alUaK63YkVQdQs44
rL/bEBTbAGvnUdrrJgoCNFLldZao2Ama338h64hpoAs4byYalowVtQjHbP8gFyPHkLWgTs4h4x+2
N7/cSX4jlztrYzR4Z41wV8GoU53igIHFJTwm/q/0tuq3IdwkYqYBt/o9jZZzCGd4/yLVTnzKKkxH
PhPmSRoEx5Rl+yZmDPOyfaYe/BPAvjGP795MryxLkb7euquTh0F3mco28sNCJ60J1uPXfcQtPxqW
5wnr93Ii99JEXi/28zj0o5fZgp0JaBxqVbOzpO5eviGBaqJ0Zw9k9lkNo5hLuCo9QWlpquxhPiX6
LNWRx2Mj3WMymHrY6sEjvMJCXcML/XD5W0u10oJr8b6mE1SETZkuRS1q0LwoxbomANCTXcayadap
JMOmllNeppHF/nogfK9j7V7SaaJLYWbqHBTfgGF3TRXXZg60pUP9Zs0I1xUGv1A8axyZAcyUFaLY
NOEAUCfZfFaaEhqTVu/uzuwceSgZuN0l6TrC5MUu8wJ82+1K3kk3EzUjWLUN4SXvCdJaz89B65XG
LmRyLBLNsdJg1ywmhB5gBvWIQeHeGR97ndKy2ntBMdYiONStm09KxUywUZDvyByEJyL5X+yFa7jy
fjbKTdcfkPddbR9iJxxnNrSZ7cvs6py6NyAba6SjdfOZZkCBnE2+h531arULKoeBKqB40cPxVT+q
xpYGxLANIRRk1h6Hbn+bXgRYelbvCcB90nc6KpKzFaFJrPT9d5LUf0QVlonRO8xygrxnpx0tPejZ
hWlL7hOLpIuaUZ9IO/Te5euXIXqgttNjYAjGPJ4bJ2bnbaxGr/tQQyxz2ZWSHyLnK813g4gBP6SY
N83qg9lLulP6PCyzRlNnZ0D+ixJ/iihWRPG2FqI4Cax6900b6frMEbyKBpllZqIip94p0LOzhZdo
6FOcqqabIVLjSrjiOMiqiQe9eTtNgXlYD9xNMkRJq7lwmpZ1HT3EhOSV23+j/ggMYueSuZvG9kEy
+JtE2optkeVdl/18n2CcbdzznZ5eQb8+klyZnbcFQNc8irGx6ryRbw5jIR61idDr1j3Pn0WGL91R
wckONNj3aL19k4I+4fKskUboczrwvsGO+MzvIYSzjPWbu/DsEVcbQdgFeXsf57rwAgDUMb0F8yCq
0gI7LaGVuWo1QxyHlnqbb7XDKJSkl8Fwf/oxF4HLL06oeMOpSoCF635XoLgzkQDoGC0vjSYGVJYf
lZ7GBLwQe8zltvi3ymjMp/VGE+kvNRiBjDJcR8aHxYxnKV4FkoFi2KBA+kZxCp9pCUt7/DGeqQe/
Tk7GWYMyr/u2riEzFjSKE4gnVddf1hbNI34AzQofWYw+nR2+903VSsAPekKA6zo6Ydc5nJIHgj8V
LksgaVtCeFgKgjj18y8qSFW/VFZYNy2kAVZMbZyLssFSsUqDIRdQ+9F1g6PF0zj3/2CHSB685if2
VWcITL8kJtRwzMzudDpco+g+WSjaDn8rfjNnPM/zzwaqVqh1q1NFvygBXlmElHpabwY+H8bbYDXT
k2SQhrBWfcUI+NhLA1nimLFNtdnPkw3iz1m9D9SYjlIMdl2vPqVs/6mnxeRXA/TvpAmElnWQ14FJ
lDo+EZ2JaqlFPH4P2jwg3UtEmlYeAerRJnQaGviM3dghXMkSmonN3Y0zPXB0MJdRL18cO56D26Ri
8tcKQPGJfVIV0TakoNnWPzwOpiDTapE8xkZSyPClApJ6KoWIkyEhweAGdlP414czzAcm63nyrL5h
Jwk4kretUwG73MW+a8NzBTZ3jk4Xc6JFkqCa5hez+ZY01waNrIMkv+KI5QY9Q0zMu3lxwuD5jTRV
HRXgJffA6Xe4dZKPsHFokr5+26osF2JGnrBKSdralkKptC86zAPmfuulzahRJumxoFG8IZ479Y9O
xov03fK1XzbTpN6oN/lISkRjZzmnFCdac+hsazXIh010eShHm1HlrHPiEw5roJm1AcRJekBU8djw
rZpLlBQYtjw+wvSWSl4Veu63ealgeftAzn8lwszU22+89EyhsMomkegeoapKErb3ZMV/hlxKfiMB
3+IE+VOnbGskxreEwlDGBwabXfo15BPDvoBp9tU4u7oewOn7ertMeYd2fVeP01KoPvN1iZTs9J1l
dg+gDwV/0w/1aRgbeWbQAa9p/nF+mgBLRx8T66AXWoGwD0iD1QG2KsgOtKGlEBy7U5u6ci1+8+u0
80A0I4guvb08wA4Bcn5fEfY/gauOknq0Eluz/5FvMKWPBHQfgkcFbWbItvsxzMzsHSZVLs/5phWP
iVviXqgVBacZxILHBTCwHPArPAS9/xsJNLTeoOeQPUx037TAioTszL3DmK6cb9VEBbd5j60+heH4
H3jH3ryQ/KBeLwW5xZyBXWTQ5Uyw7kNBkAVUOW+OnTXQCpL2NlA3VRQRheDEcBRccSUxJBP5tuC3
TNuprepexVrwheHdxhbdfLLNKDv3zqCr0NQyNAJ2Xp96lBoBuRzyQsHO0BaugwljhPV3XIKRea6t
JQsJuKZqHagLl6IAXZhoS+Y2ysPYq9QAWxZBfb1KFSRsjD3jKYWlDDqeOYAKaKUNo8hJSy2gb+RF
Yss7zV4+SFMoaX8w8uVZQi9tc0M+QjxCV2xIAn0wVY/cVIt5htWtQKqMPGNxpyOJ5NLDMiKwaGFQ
tLim22vRwEAEAVl5hLkPJ7oRO5q0UVGf+B5nyqF4vtXF6gwkRxIlJdzri76pNJy49UPaLGin80w9
JXfPI5t5VjGaMrjGMRH5IzKXksIgg+Vzi0Xf8K1V/RtfR5kuGrX+mJNve1nx4FykW4l3tpuG93Rk
UodatEbImmikJr3Tqa3XIjMQBc3S8AyOWTpQxuTQoFrK0QIZY2WK/6frSCz9sW2GMKgUlYaYg/yU
7nFMkoXVHtn0ujf9nDMLQvL/XcT8I50/g1jd763CCUpN6wtDI3theAwWwJ/tXS1vx8unp7jRNR2v
X/kk9BHrLUV3bmJVvHZV+x51dqUKXLsDbWlvWeae02fnrtqlSKFCon86RQiWBV+uEfvhnAjZJjTD
hTdiMV62X9I581IGeV3Eq5uh2Fk/Lqbyvhqmj7ydl3Wq2QRWdEg1fB+GktIaOdM3sjseQGV2b+dS
PSc3dUDPgmzByEZg+zkdd25n0IO/Rypfv8W0BYeBlFwg1LFiqUgZwdqxOK67XUa2liFI/Lvx7V3M
8rxm13zgglJQi8vy7QNDbiGzYlYVQvpDtLuZILPupLUxXgMUxscwTuXLUwdcThtmiVYaGRPzYZUD
6pvMLmR9FMpcWb/Gf31DT5CMoLdmEfZOnVrZNapZ0OvSoCPOTRmPC26BXsSOjhl1U4D7pz9+3Bso
zKmEh23Kpi/fZqbjX2rcgMYrzWB+GNWJ5+ALBH+BAW/QQnFQGP0oP9TnJEhO7J0FXO86KAujm1Lf
jqVru3AG86kEbD4fAsU74YgwvU/iAncogem0AfvF6lbGRg/r3l2z6fXJ0KNA922ap6axnMn6aSfe
Jb9zZbGHjQ36lg1JGLH3mxy3mP/N7SpEh4iIfeWeKWh7irt3/hi2acGuKBkif1WRMXcb+V4GhT86
p/huuksxb90wAlMdhfqWIewFcvdS9mNzXwbZgo4aYcDjOx+i9UqdL3JpAsKrn42vm7L0cav/gpJz
+WTgCakIr0UCxuO3kP/6hJPtMhFQNyM9tnw7lRVXqrXLpGOADhta5VlwpBGhtX86vsXUWow6kjki
xPRI48IvYvtPm/BeTNIgedbidNAr67DM03U2ZzmNdSLT0ZBFtASYliRucj+Wmv257PxJR9iQQXMZ
qN67oRx/FVo1TkmNsuXlPFalBeJNfWI1uC1TyEJpQ0H/NJfhUKBZKmAzhGvKsROX+FWpn7RdSmVR
ShwBYQiWAPX4JFTdyh9VJMcNEvjdXL43tMffWbjR1+y1T6/QnTG3AU5e0PdOMpMKMbvi4ZzQOqHP
2CFXujaAVHszjuOFDoXqTENFuuah/t8hF7N77bmp4aL+Ot9+Em7rURtDeBJ0bbnTA60PjgZmPCHT
qjlSPteOP62TSR86Xa1f00gQJ7sBGuYkDgwC5egkWFynV7NBcSsjaeuB1aZOr7O4GJAaeWq6uwls
AtbKx/S4a6csGPGdxUI7I5SQy3JnYgBFILXDXP5Y9TRVF3s4hGOrm8q9tw0ZTo/lLhyvKUqqS40Q
yBwL+4+ok1e0egS8dkn8iwBpDBS0509TC1Vb20pYjYnoFi9jLn99NM+a6OcEvjN5ZAG/CLivfD/A
gXvBDTToWENEqH/cCjO/cAK9OwHS6wDnJLEL+oiAW19KZUU+YQfjuU/WIKw/XZ9gn+25vHOBSwaF
ltUkl4StdfvOqhpJ7Yd3d9eRntnjAegHQA/O8hxHmFbc6IPtq5am+B8OZvcawTbCCY54gV4S84em
5HTyi+M8upr4re2hbmyOhUWiombuFWYudDYg1sTXkIFKO3yxxvdMc8S+STm9nvymo4ae4XdEPxk6
suFDn5m585SDBZYSNBlg7vOCMID3c3pCkVzI+Q97OUn9nlHnYFeAs6qsaEKs8+GvwYKcdlZ2LZNO
vLSVIYqT+BaCp6M9Veu5eLj15JK9OuMnnBGbAR+lY/R+9YNmpQY7BGieGlwE9qXdmYx+qNPiRU1U
jD97XruVcx/VQyi5kE5FQNX1UpY8nA/C4BGJzC2VVzxPXYVWji0SigtK2ZHAr25RUSdfAzK22lr0
kvbN1rCjdWvhSECX406mxQRLv2MwYyumRnriyX2qWN9n1W0oXGtoF0RLq+jS+CuJeA9z7gYSf2F+
he6tmU+EO4hzj1ecF6zXYwy9ntdxyhuSLXVBhPUtBXSb9z+ZTTcy1zGZVmJToBXJ39rrPcxddtW6
4mA6oGlZsaM5AC/qZ1P+QE/Yv1VnX3DheqWj4IyVuGYJXicCqV1y71nNjfzkpH+DyNfs81kdsTjs
iCgXqykQKcQ9GnSS7HYs9BDU9WPhTM6UqwC9GwdDPZTw5h5hYgA0s3auYvepO2PuICQv634wPad3
ngJ1URNng0nETluFKOzFE/w7fFDXQQRE+4J28rkeX1Y93lrSRG3fHrcso0Mlw7C1NoFSAfdc+KqB
SKRIsCgS5LNaLVw/GAxPyF+nciM6MbIO4osPvHS66nLqcr/sgQtJvdmZzhXqQBrZ5gpCK+BIOU6+
nn0AKVNbP1aD+PpXH6XnmILchQZvoTv0AXN3wGD4UcCfJCEm9Aajkl0PGWTR6VXh6bIoWKXaMC3h
8inxIAaRIJNdtNTc+nZyvtph50PI1AY7JfOmmlY6Ttxv8LMQN48/rFKUKL5CiOZ4d4esbb/KK8DL
B0k1G3tzx1dI1eYg2TNwkodnVleCP7Q5pDPVtwD6cXXp/QBEZV993BEEyy5iaYwlfM1kU7dJiZIH
z67DBwPCNUUC5pXmXFk2W8TV03mMtk5oKVfMoy6drgEy1ZHYrPi+lkKVdDvqgnLuLBE8K5XU5h3q
pVUmCY32xpCuTQP9Ue/eQTJ+hNQeG2GDvKCFGIfaPAmcvTtsG7ezXpH1HK0npe5JmwMr0Ko5blYM
3peLimg+OyYU/2BcweulLqy8FzekxX7pFbtjuzqpNJj7ngvRKtUfV764xCNpVROLylPdEQ4uxkUX
zoGKmKFeUZ03ff/0gfCo7V7LmP7Brx036IjhR78VwekyYPOnO/e+B2n6o70i3AH1uCValdYrfTom
DXudQ56kUP+iw9LVHOPwgexlWqN/Sl4EDCFF7BZBESBgtU4tt7r3z+hqgR1Y5yBMq654wmODGeHb
kpLE88QOhHKaVHnR2VAkgH9+EliH1t/JYArYGMyA9D1gvxrNs191/sXGrTblG7tN6C2LF9as6BwQ
twxZHWVHIz+mbhvCLjF6xEcK3glEWzI48LQ+zPHtqqS+Lh29kKfuCRkM0EPAJy/77JgGDl/zBaiy
qAZ8U4y16tnNiCFQEK0IH8upj0eFtGKCHWtSSksVeeve3Pau+xsDfGmIgr3Owgcwj8i0aSJoDp0c
qh8jO6Q2vk5t+mFuHLNv4d21BWyfL4zEny11JdxcDfqcSzXMSSQ/7q+Bz7bBRMcOGyzLkH1hrB3s
qFeizfNb8j86FCvtsiX83miUIQmwypdQqfoKatF/3bKIem4VsVTX/sRTQhRp8zdEr7UmpkFtbpUG
TTEigg58Q8gkBif0QLXWml6eVHsQLmdOHAWxWn4oDXJHJ4pS4k1GMznDr/LwR+z9oMC+Yr67I4Jw
H1eReYMMPPckNk8O2Lq0nCiax60xzl/ERIlLqv+E9V8ao25YOnS/gUXfrZQwZzS15fDJ55QwafsS
tn+idKupaBJ/nz9kZKqPQdGVsFjToNKtcmFC3/i/T0clwNCksr/6iSD70RYP8BaaLWy1OU70SDh3
/4nD9czkyyzhUhWhKkOuROTwGom/e365YoBjUzQTN1/VE3zbHNeU30wfNtuDvbC3Ml1EvafmAYmy
uBO78Y8Vv4ktPaApg2eRg2BZY0vDITJbRHTHzNDCLWFlyn7bmEQSliWHXaCDV/9FItQ2SxvZKwDs
yvCCxlPWNFYyoVAbaOyAgXYZkEeR8EWXElLLcqL6q5OXumgyULV6ifUf5Guns0Ln23QbGbj3uwEL
jJzFibdFlkp7wKcP9HGi9HjqMzNu8fjDaogVB9x44DfcN8J5Gmkyz9Sax0nHBUUNNdOsRppPthvJ
f55l/wk01j+CJSo77t1fpBYpczXjhJjbFVUfWOaTRgasO7MSry3Qd4jM6ZQxp7AH0VDQgnszPfe9
92Nnygh5TZRhBSb9FdF0emkrRAUzOEexllToHhr/xqdPYesRPGZXFf/pnO+gfgNjmvSK/z5F74+n
V/SFh1ZE0lbQqRER5EfrjUruKrN0wInqOR4CA08lw1d88bDEl5YXtuyLG5ci7u6dgr0wi1bvoroN
WBA+af2OpeN/o3bedAa8bwqPq2JZzUIgpSwdwbRxVsgBMaEeQo4z6sjNLPkVZey0dQE/+nl2hFGj
vCpjJA0cHqGf8LI61oHP0LdcfmBhRTTmtSvz2o3LD1muu/QVy2Je2RSxwO0b6OFlZ9UvypKKoeb8
c9cNRNyEhKDfn4UC0qXoLMIGUM0/qRIfnxwTjfUdXGgYjVZddHqNv+m2nnjFdojJ8vNVVcjcd3Xe
l92nuDd3qt8TbKFy3NmY99bCQvIMhg4nwzeyEnEmqQsdnQWzvR0CPv+2grx9Dp3qr4lxBVH1Rxpx
M6/gRsO6qc4QCoIYK9ZKNB2fNZXyCRi/Yy9GK9W0whkowJe1XptbbOPm1gj5MwmCaaSr2ARR8gzc
FAb4djW7dApAW4K8fxpdU9ubwSSU7PZkb9X1osIMtkevmBdkFuB8UI9/HMUyT3vVQef7be1+6vat
G1sybyk6w4Vgr7IMYLIrYEwxaGtzS3eMsxAWPj+jR3sfC0HXLPFSmOO2vI6orofVcsGzMR4BRA89
RmYKcymv+V42NTI2clB9YX18QfV8dja7puN/WeqIvOBPrnlyY0MMPW98eNYfLYROtNn4YlJj4nei
cvvAcULr7eKkeXu4VsZeht+cXo/TU3+21LSmDM/BGvjL6+o7j43mCy6KRfjqWTXcXGpbUofHh3uZ
r7iibSCVVyr+oRbsWAGUBet/JW2sOjjCZuNspf/5TgtVWEhshOgyAps9L0zpSMpxWp4XSWvliRfg
ABPyEmetIWC2qk+H8sMCyKKpSpBOsCPKYGsLBGI8fRMzBk/kQfu4VmGsf9i2vUwP7A82e02oFPn4
GV3dXvew+uuf+t+4MVIQO174Hl0hmfxvPHf1yYeteChlIEJpcUJPF2LrU1rNF4YpEK/pIjz7bKvz
CRjnNSfDGgzmIb23j6qEwNFtPwGIdcGTESB40nlWkencfMe5XQjiGJgdPuRAx3quc7T1dg3D+9kA
dU17Vp0/wNJziH2byzLNh8U0/l/WSdrUdoxlhezmSJf1XPNSERzxHhVVNwAz3+Wo1im0VPJ/taMC
DbEa0duS1wuODg3k6UwJKrDZuh8zOUA1/ti5N3u1nqclih+9IAZpCP2i35idvCik+wDbdhmwOfBb
Epa/IFp+TMT1mIkA/sLkXYd+xNinHUgHC+F35PiRwlod4ahDsJB/NNWSG1mjcKb7ADPQlEukHWqW
bK/yM0jUEtEOLijdEq1cl4NDjuzQ3exvPVeUfRYZeLtGn4D8GPxJEpCGMBRIr/nywxOCpgKQqqMF
bVg0uXv8SwsBr2So/Txfsr1vf12uiKQMMNKNwtuVtBjO+jgbRntOl7u745ftJ8eHKEw4zHsrwdMm
dWTpWoi5m+xyKsDgHM1S6rB4LLiBSf1F1NCahQAagPNyE4xug/gtxUZWEVZAQhTdX4qq3K2yASjT
8Po9CS5EcCdbOLaH9qdLmZYGXQmJQcOMqaR/4IroZfMwY1wZdFkpWsgDGodTP/F549U8pYD37qAh
ZuFViLupj/dUv/m6MkJHSAbl1a4YkX7ZKgQtdqke6YgeTqMsbl/6C1Pht5iJGGOtnqV+sBLkvege
i8WCux+snMOX7wnRlPppbQ9RhJKJiTA2lsvXGSJ4hzBfXwGZOn7RxuR6yS0JLdEBr38zTMZ0SN9D
P6x57rf1O5XXJevum5PH4uK1YvdBEIs+s8k8DAGwRfJYuVA2snomhghzAqxWWzO6OmfvRh8KMfaF
3MSZ3Mf5vcVfrWOA379JAdTr6kxPiR2X1YuTJ3B/1owIyZc8/QN+mZ+fxLCfn3nvDJPCcGw1/kfZ
bfDaGrbX9hmjgw/9Gk2l+meIdg1jvxWolu6YMfm9HzkdfhU+T4SFNDc48Dd6ksC1vyETl3075Eoa
kATf0z9/p5O1uhmPA1VFTHSXeWRB5hLiE94ZdsaT+pSrPK2KqXL9x+fw8L0WzzO8hluEB5Tgm189
r7qt8Qu0W6eOMN8VS6LgiDQsOtoaRSTjibVzjxR1cWWVq99q54z3ZtSNEYI14/ZBr3l2tLOd+5Ij
aNBNzE4IVCCjoStfxf52bN+PdTxTkP8GVDYmxaF5rPcLYtHFnizlMrSZMvsYy46REksVf8XAmjRW
eizFu+PG04zY3UILMukn5nNBGehaKmCLFm4IFNYiUQkn2VQk3R8UKZD1xeF7LBDn5ioTaLkexCKp
vDmoNh9Va9RWkqp92vKzi8eU6zaujlO/RbDGB81Cy2R7dGI1BmA2wza+AmfYIgrmrD9bQkWtokLn
Sx9+GDGCjfvuJdYQ+jrTPHtFlV6Q40vExs9hFLYOp68eJCOjDZXOPwY9zK9N+ZhMjpVyarenMOEN
YocCY138Aa2GsU1zqdfjLxx7Mv11d4eJmrEirCoL6yLDmm5u1uxSbUZH3/G3SBWZMYn6I5Ouov/j
uVQKEYZTaHpyczZKlyJY0tPaURLivIETxpa/Y9iGLMEiiTyhgfiWOVOQlDtLizBrcsQP0d5fCKTI
ygqDsuhvcn7wy/s2satUNO08F2btEzbE6gEm1Q4GK8tf+UkS2ZZA163vXR9Fd05N5SSkPrrDQUPF
ViNO/Ucq/IHelLi8XHpe0tz1uhGgdZTsGyB3Vj0D82P+jwUaY7Yw57VDop97b0nXiNf+dFeSobkd
0f0QDuC3NE3x+mkQMomi93AkAW8wmS3H2uC286vP4H9oKb/MDetUn22oQwN05G/jv1ymxirizHY6
WOqaZIpEVqSf0zNc4BB2CnoFiYoaEe4Am9IhwpBs+UnCzbJ4KH3DA2z66Z7TtLuPJL+397UHceW/
igFwD9KlbXityHaZvzNru5VhLj+dxPosIZ/HpLs5DX8nDfO4A5V1ocfKjk3sRtLwggljfwWGPBQw
uTIv9NWQ2vdmIXiLeZnRUZazA/+TBdPkFa5PkkGO3PX7eJ7MBz3/F9vggi3ZMBlOgDDPEV+G4n1v
xQiHxbZ80wMwLmZ7vqW0KLuMpiqo+WiP18eAya/jgI4uTlCv16dSncmqlkx+ms2PlcPzEUTfzpTP
4r+HhM/gUtLzum12fSYrQaULg+z+M4jCXxtdk4iUGp5rVYyhXWcLQA2i475ZC2C6mc8YGp1JLNX+
RLLKBcxNppLkr7kM9tZd02aPTQH7CxgxWDFIwuAMR2ENapp3DpGxiXV94yoCEemehRWHSuSG1ad6
H3muz0ko9DFaAFAmGhz8TqipgP/CtrbnoziROmtttaMn/+F+BlAIO2eceUxqSpgkr+A3Jb+7DM3Z
pxvxx2Ha47xY5r6Du7ZABIcjFrPYVdaaeXxoICpZaObN9V9W9lfRjk1XWyV8Hum+2KQXddUa9TDX
36F99VRsD7tKwWYrgQR2k90AWWBQDOAYlnPoO1tb7tGRKtMWhzHEbgmETgLizqBILze1AnwPEpeV
c+xwvnFbVOba4LFE/BrISwimray0swyb0L7qc/Tn/Zij79JOSdhO7Azo0hXdesaACF9t8f0o0YJl
TPS5HZiK+8PU4PEoDQ9ojCoJxHolc8+JW27PS9BedceJEAvIaefeOQVIzAvzS4riGIGhn+l5VzPM
YunT6p0ZIxIoZEerNT3YHjdx3c24iR/U+4WcPOI/Fmt/Ydc80rHb8BfA2VoA0CAnilRM14cTr2hG
cAuBWwpXVz3gpjILErGB9nKb+RkeNRZsraihmQh1RDr5ieGR57or/8WKXbTypJU5UfW1dA+436Vk
fo8S0iNDdsbkr4k67FheXcGrT7pO5B5xIwtVag1NVA78UGqFG+bMcb7+V1Pkj+HYfV0+I0Hsd0vj
+H30Ib9kaSj+4VaxKj9G/fNggQyQ1YemCd1IkIqPklRdQXVh/Ac6G41C8AVgkGQnEUVzuFPsOKXX
+OpzrXMMG2I9mZnsP29dQyglHr64vv64KPgyWwql3gYApMFW0XOqPhRzwSfMNbLgHQK7teVxfd76
ZnQ3X+/RcnrXoOuaw6yBRis+7pv2lTtUZ2OqqWr6oznd0dwvZqfBD4oH17HDhuv/Otn27MHoJf53
Q78TucFsxs2l9aXSN0BnWIn0a7FbkewrbEKv03xLQiuuleob8ZfGiyBRqaDlvltfdDPFOiMPM+H+
l2z2/3Oqczg5LMVDSQTm/Eq350jBMdb9ct3rbZYDffvWFvImdkwrI6wESAjCGJrCZ5darfR5h7eS
n0TrWVhbh8RDId6/q4ZnNxy2Ov5+ryvVKXr/B6sRq+cnKGlum/tZdpDBvQsAmwBqBTsHROJzqS0t
nPiBmG4Ug6JkhiEX54tVMtb+y+jnBXg+kSHR/HRJxBievfWXZXmio2W6UmgUgewUz/wHNxTrJskp
N91tLqYBI+Pzb+s8TjlDRpiu/vAzRk5J/y0Iz8WUL3bnYC3OOwEUv1kly5UOT0YGet/Tc5m/koFj
YgeWB53x5O2FhmT94yWebezf0utBXriA1vnc9AJJ/mMniGX1LQSBN9g5ugkkVL/m+koAMY+R9m8A
/ke2DJLJMPRTVunqBoCL6+nchwWZb5Xwb4rBpZfZ/GXrsKiY/sm7TBHyctCqITkC8Xz44NOiD0bI
gwCY1fD1z/tBy8ly2LRde99fa0eF+yt9lA8itNkiSViSlQ68dT2ek3rs7oe/6LMpgkA50fS/rRPy
4/rZ/OItTryrGhWGmN4r5b7XvyrdQ9MLvYjYeg9HYk4XnP88F/rOrOe0MUZz7reM87F7cBuHuXLs
xSovWfVuaIUbVvfbnbTTCqemBk8lu65N2r0H6/GSFixANBLabGDVOkEQK/1gZNduJyVs7ETc5fd+
3FidvyEmOVr0QpdpuEEhahXV14a5bJLRvmMJSww0Mvlq/m53j/o4tUGqU6rSAiB8xPR5h7YTprxg
vW+QIq9465ZSTYyAtZl8iH+196FL8VKD+qGpTrkCUmpkfzIbCXFYhF2QgsT6fxeEN86BWdZ4u45u
4yJdSadYOjDxkoSInxWOc6GKxUAiguoTysqHe5WHyW5DizHl4A9m6ypUdiFrm0ElR3/13DReHs3c
FkWAv5RRTgOs+VA5h3mFjvd5clvj0/QDrdRcXjWNe7BkYK8fnWbwNt/tpSvYXpf1AVL4jFjGFJCP
3pi6zmFxasGp+YQvLC35ZZy1dru1QagkJWWmo4VE2yL8OuwBmjEXf+ylL0U+Z8xqbF7nJyOWJ6MJ
HNeXCZP436+n3sYTJC3sNoci6qFkIOujqPeXp4T4DgjWHt4ykq6F9mrgBT2kEvfQGYB1OWoMqyLG
ggrR7Vb/brD1Xr1eIOu+2sMWSeWW7yB58QxnesDekiQi540B5EOBeMEILlSwBiJwfGnNC2RswpGH
VcTodb5ksG7hEO8NzioGW6Chdu87IzzC6G6PA7Qv6QByDtDcOfwRxF9/nJTDCwMT4xCwFLVAjOex
QjtifYusSKMFpr4JqhF9JWn1buOtCfC3JUoonZHzH0CTSh1OiXd18/tEM56+Y3zYS7SJC3knUfZK
gWQQyDvOdmEHGmS/I+I4p+pyX776EZ5MNmV6XLJ5xel5xiBCL1rYAApE9tec/agY46z/uCDnLQnV
PITxYAmG1oVvoXDdJ1dLedfklxbS7rwlFOTNdl/MvcN58bi1GiRoCXhf5C3Y3CiywXgdGe0xwlyH
zSwK0iClMThXedT+ldiJ9aTztVCA0MQ5JCdRIjFOzrewTc8F/S5PFUERmHlZXVKvJ/VnZptNov46
DqNnze/sHnSljdtGCpicpHZInmUlnSJs72YjPEX9jemk2ZeHik+WZkR1ld3u5qzehvGPyHCDYShX
Y8PephHbaRo6onTxOELRRcPdE70TWcX3b4D3Qhvj0GZxlYfYadXyWdYyckmpxAwAAIuU0v0tonfs
iUINKUCW9qTIeM1CPt4QFG0bDL7u+QHMCxfy2Ii5Z7HNy8xUxZZOsTRotWjZng+JnwlKEXatTH1s
tBepFYqPaiRi8UAqEcY4Fq/rCC0yiWfcxaCKpWF+Mb/kwPvQt8DAN73Qwj+1GBNr9vNvMAJX6vJm
+vbUb5uzg7ui8vdSYRpaoocfsRzAT3j9bkNYXQpl1LeZW7NRBg5Zlh/3X8DOEr/a0UD6bicHiuPF
NNMV97EVALBsObr3vUL2mc8Xyy+kVhJZDut2y3bTEzLaIGJ2IldKGrYRa7Cwl5g7oQO/U+21G6qA
QXSe7kt9/19n8b0+5qqzc4uK3sNTHzD9+8MRy0NGCbGtjhWQVqp2oqle78rRNKvBIbJ7ghiePBBD
Pkn+IdVRbl7HpUXzX3WdDI30brcdvZLcd7E4SCoC4hPIqizVfinnf2PCZFnajASczbsB5VlV7u7j
hu8olMIxgYhy77XAe18UAuzBrvWCpTviBI0KgHwTwd/MZ3q67MkmCesYMKv3l80JEl1m98Oz2YcE
VzeIwPktzLqROf1UN0kPHblTQC8NOwnzda9FcXn7swo8AXKy2RzSp2sTX6kKIlSIUbqmMHVBktWW
OML1T2g+17RCklUun7f0eGwTkV2ZkBEr1YfyVmkdXnubdGjK14etbZVq+Fr+32tKjqCRSLrOKh0y
ww/HoBGAxRDfui0z3e9xNlIs4LbMPfeDPDrnnGSN5Th8EQdYAkdId7ynIpuOybPAPupGhc1bUTFy
rE6ta72oMzpU+q8Gfz8Ki4w4MkTkBfez8adPKp37c5G5kOGcxojQ3ePAS3BXN0u7zIsLLWPrZPoN
Ciqs2xjzxKfZAAKl9ftWX+yrLv5bEN5v7TkeXYqRfpsp4+IilUBDRtmkwcmRJ3HjN0oOTUnT/PLE
eHU0rL5Mn6pDqCAuL0Vszwg4rhMG0V+DSDGb3kFp7ztDj8tcTjrGjyCTEujiorjtS3OP7U7fng8J
VypIs72VAlGHtNK3KD/9aTEKci4c2Eao/VRqf2n6BdhSSoGuZnlgR3fmNY7w+Od2nJh8v+CELYt9
jTbUzphs1d/nTP0/Onj4O6Ihl3FXT+FhU2Ufk7UX3x6cQDLcnOxIo4WkKaif4i7I11tJp3xaPWqY
Oe3JQmkq1sLXi+4TRgsRafnWODNx06FTRbxM901iEqUPca1AA01v936SAnyRUz93dcCm9qc37VtQ
7Bc0jP4VWHmRTmOVZtRTVESgZANSqTWlk5MEcuZD2TA0KJ4Pp6XnZsUfjuKyGtQBPQ8ZQAYEL02K
e4RzTI5XRvcD6vQSjNi9eHE3Axphc4Db6IJyTeTji/bf4896R8sMTBsECsVl1zEnsnSgabUxluTO
OzUFIugGYIdsCl3DGQVxyZ1XFso9MydcF98hMGJpceV6wk6OoWR/nb/2IggN0wD1Y68VKSzQouJj
U8ZynvMtvg3sVPPfSmau8jXnXPFjHXqYZMyX2HMOvl0NLNobWxfIn+QaO5DFChNaJ2qiw2AyBxWR
7jqMb9ivLGjgYYTJn/NZXsIQLaGXqtSbod7Ii7QTvO403wwQLFD3Usf7jzoKc99U7nBTZTyzRS2i
GsxLMFlLyMzR6WSJbWXD1B93p2MxvBmvZv61WkhdduGlFiNk4XeGdY8SYyEdl57Ntn7lHWrkXmme
1YjoPHztjseNjEc0lA5VIAMHMz1YTyxYprgZp5ahFk1358ll6Ga4jbO3Pu8OQ610FldnejAb76iY
KMlcAz9djMMXq1Tjift6OkDmVmughRZbbCG0lRZU+TpO7RQfolh8t9JWlH6iaZNUguudAMvz70P+
3fH9e/59PXNwYtmSs2g4KmpH8V1EjRqb8m5YfKQBxjPv9sCbsZr8MnLHHdz65jsRUodDHq50Is0p
s1zK80CUIaixNW4OaEH0/C7wpWtLGFEUpdJ3RzgJSgzgH6pZhxgZC7tTCv/6hYL8E6+if96BeeHr
rQoEPZJ1xykyi1ZmdN3oQZw+Jo8exTUxGuHbqUBeIXJ0W+mvnrYmSyJbk/3cNVTtS3f5uXXdszb2
3NRWZORyYDRhdgN2+MsLM2dptXbkBQNOV/6tgNoPOkpXkyvLE9Ln5CDHJckn+/67XEO+WsZ/fF6w
pe8VeTDv0ge3VkjefNMOAqj4QdueqUyM82lokkzbl8cSOgC3Gvq6I0yApzGeDPeLWWQs3KjU10+a
427onm9lSgG6KAxbrbW8b4nByQg584miy2foawPEKHrAEYbCfydL5AXjLt6GuCKff+MGkqSSWwlW
oIna+KPKgLOtZFdipVyDrdKqLmlQlkGSWQSYVFyjyg3bKVW5ILnVE/rywvJHFCxK9iOHBGzrv+AL
tRkuauChEu0/xx6V4+j8r1CzyHKMUOq8qVWdqUhpBPiRx+xp5wLKUq7hyfzCgtho6z+jj3HIEZc3
YgwZryi+QEX3yOJ0GGtQU70YMxRFUe4+wNyXvf/CnbDTpW0rMQxJnmAYh6AfdXxkLZdKVXTujiSJ
HsnbWsnxgQHpl8jlTDcOXnkjkOWrzdeeawMsXLt18Mk2KydQTvMZ+VGQnud9ltylaJ9uTL0nv3Qn
jZRUxgaupx/QH5yMhe4rCoxpsFQvsiNDx4p3UPIxKRKwj85qSaWPT1obcizgtxoQHBXuakCGaV2b
NNqFgJShIGbljPufmAQyQ/IimNUlYLOB/Kf3aymLJjOD5QbBdQEyyhYj2IRdziejMB2qVkQ4ecOJ
c5ffLeDvKylhulHpxqx0WN/lMgRra6rhUh3wYrg8lF4jj39gxf3b1dOV8kfbENdBhVkbI/HGxLF7
SAHN9GJiXVa3ZAvjTJvHpOMnFZjbcx6ApW3U7kp0dAuRkyCyNFwWOq+8reLRJyJjG802JKnHadAr
Mm0otxPkPK75uqyYRQNGvV5gYa+JYM6XnONZfd4qG2CmVRtuj7QeO/1RodigOQMVbB4/sxd/sRHi
pLhclos9BJkgQ/cVJzo2iVt78zbyT2BgLwbwRbfv44XRKaW5KOPI0caRAeoAsYw6oW1nnCTIeytA
ZaG2tcNd78xMh/IAks14dtj5PdUeP5FX+d1gVuBhDqOZiXJFidjr6OWfRDTmzwJbSSnS3RqTbW8C
ROP5ReQ4mMaCsgrvAmFWQ2aJAMT2f1mDbGjT38FqEm54JGLjkAVxUobSwx2L1W+13BxQp9588TT2
oJ+MWymP91Iwm3Zz4lo/3x6gh/HMxOTwsHw0Duw4tDzlS23o2p2Be5U0qQCzq/AtDyXEFWXqfZ3o
P/q2kEFEm2iqNsrrwwbu3QZdNN0GlXZYur/QoGn+Robl86SFpyYdfAjzrnPCBYOrhOnGziZnPzt8
uLN/fVa8MacohCi4kCxpWN52266ZvOq6f28X+T5Ya1lwvv8EG1Osdyml/w81az1Vgqimbp82yFWH
m/rFBbjB6tswaY0hHBnh8pNiFkGe3Aj2rBoOMSRLaCAjl857zxJiuhnR5yJyzA7m6y5g2SEb7m8z
qGvE/YfhO1d/I7TMa4VuE3oOkTIjGXNcC6p0lo90P8LEoeCIbOE2ME4XdI3Y7+iENHdaioiHy9FV
CqYRatFnyE0a1Y93wzZl8PclHzvGWhzQgrC7DVYj41GbUyhHMi3QLwGE/msfaZTTtDJOICuX8XwQ
NUcVuRz0rl6EMkfbbvPelnJenr7IobzPdacgLt3yf6NhJcLR6zzpj7XDU7DQqZ0Lo/xbxQwUeMRW
Jckb7KOWa9QvDap9ahdP518Aq+hE0JPXpsNZEK6ybyF3TTG28+3EH1wIp8vb2ZPNMNC4osvKErpO
kOqIizAwft68DV0HNwOocSa8saxX1eG+bBkXTjgWWwmpjF0Rj7hUrJXgDs/5l9rmeTu1YN8V+e/O
UzzQmNllmcoJX2rN3l6jsatM3j5jyNzDiCo8Xk1En8rjGLVxQsxGWptoMaMLh7jPkrBaUl7RA+AU
CepV1rGR909nYbCB2sShKWaGGe78bHlk8CI5dndqaku6za/FnlDYOv6zn9jsjHWAtsihH9jl5pK6
5U7qSjKkMHFbMjjMCVr6fUbgT0Z5rD6YlwEFKYabBNhdw4BCvlTutBRue0WdKFFtNqSBsfa8/svT
t7fKH697fRCv3yM8rp9BJ1WxWgZC0/OR13MOC8/vUR37/j/LBZiMe6FmFQLJFQQdCCIg105TIeBv
dWZjkhDs+lzdLXx8W4hUHh0esZge/OpVAy7oUMU12KuiySUxfslofZHT/RgY9+XQzr2MAhSf16Gr
J4hp/ef59vNX6E0SWe9NuCZqOOn8MfdffJ6BWkA4FJWB7VWO6spE1l+efLfaWHNjDDdQiS0X6XGe
kUV9phsNqTD1ekceRLuKIJx4Qa5nSuQURh9f53mPTU4mFfNW1SEQxIz98/pOygCX44J3mpXrgJdC
WHAVPYXoRARI24NdrIQBBXBphuQ6lh97BATdk7oZtXi1vWAFlLnN1T4MTRKCirBmCOJ1tJYAVI3w
D5pE1Hn5RvIGVJ76uay8aEY8WNiH7vuGwKYoraAbMfBALQKo+nMah3fz/McuAYdebwSd/l8aNHhb
klv91vPVb2dop05znu1iBr4ooeyMYU/q+V+1WxPn/pxu1Bb4adwTiUKSDdgLjEYnHpOrY96+Xg5D
PXpgeOH6uot6VxyJTi2/YVjuF5UbigfRJ5ENnq363Qky9SQ9Q2FeVIx4vN3gMEFIV5uFYSL/PAkY
YCklBMZjyiV7RFI9cDsMeuaXyo9MIJrAahOK/wmJLGnLi6rPT3avBojQRcXABHK1m0j1tva4LHnZ
el/qUU/+RkhmbNVnggGKIAWVdj1Y6/oXyxDB9v6/TQFtCpdinPd7l841TRhYGvrTgbCENRADOOJs
TzbtcS3ZVlGw/LmTj2zCxaQXXItpnIX8u+ZcuWG3bIYnZC/IWwX8748cm8mb6IwMuAXhvECE3dFw
blucwYR8qfQT8+OG87PPXs+H2XHhiFVeE6EWXmNHZKhWCtz5OTWjXj1O/7s3i20/G8z7sHrR9riz
mdlw2CiV4wxyh/+XD7sxEy9kssLADOVvP8cCDrMEZtdRFjG1c11BJgOfhzua7z+4y5LaRw3Licd2
pjJBWHjFubsg7kohHtaBB5S+XZHXEgU/J9we0IjL5APwZ2BeOlqvAXm4FNFfqpE+D1YmUvNQsr3m
PvYXvJb8yuCrhGsShsUEwTezgyn6WqhnIg/PawFrzVjx14ugQTjHg55MeHYVg8Fa68xv5T91sVg/
TKb0RdgguHGlMk678lwoKRA15HKnkhpPQAqhhFQhZtYRtLsOJoTwFIiN04lEEb3cTmImtpL7x5K6
i3w1X8EmkNWU/JG3NWhAmhRS2MbY7LkH4DLFGNKIFHAmPQqXk1Gr9JrUfRp2u57a7VvjD+RzV56k
QvngG4OtY4PkMowSu85xRlNXppBBC4ONyVSLUGQn65Y4TDiSKEvEzFnVJCqvcRL7RNXkvOExuc7i
XZqNqOWQ5js7vYZJniSQx9hYQu8RaSDnGovlzV/l2nCqMzPro7REjrMI0KmzCmUhpiFR7B5A/27W
dOj65kZ0VC9mOd3TWmwhwUv2J/d7ibK/ysAn10Pgu513oMi/lQQhJFOQ7K1zLpDYnpsfz2I1fEp1
ZuSD/xK4DnhZ7AFCozXmrcdSn36uya0MiwhKPuUkM8vFtfFFUFQBgVYjQu3SWNr/jyjp97LB30p+
1sLXFMKsWp7uprh9YbdpytGfKHgweInzJss/n33ocEZHDAxTVb4n533PRXyMUyTCyGaBeUffYJRT
DyEuJpOeAOVUpDLKgYeCO6/PWnYp8PDXDgcFK0IYI5OEhdeYQkH05tJadznaY1tGzvUtH3wMP44u
np2PBOcW9SAB5zz/WfVGdjOxs1FUhthdJyM56UwOAbb7Zk+g+xJoVNfM1pd0cZUmRqM4zs+9F0B4
Oil0Mh44um15Y3YpNY+cmBC9wP+wrHvFiEGh80ys5reAeWMShRYpjz5b8ggQVbMJ6SRBh7DqFMja
UQmVSJZOmgAgcPdfei0n6p6CvP9TZMOm7TAziZDciWNSMd/F3uKkZFgtp6vqpsT2eBpmES1u9UDq
byoumXV+84na5D8vtM02yjbOwjcm0J69Cd4pQkqxd2RERfTNTI4xrCnCOON4lSAqPjNnKrpgtpy2
oBY96p9BMwzISQAA0eJh0eezvdKG6ooSUEzdyV5GHH7W6ZqOg1D9QsIWll0TFYslUQjVomR7n1CC
qAr60xFT3voa5DwHK1o2ARu5NQLgn2p/BVfeekCxLNQMMF9vj4/mBU+SiFvI/KyoEWFHCvS68bWk
0jfPtoLOr/GpwaR1FUxONMhyMpiDqALzvbjzvKNIwHqpgg7qR4Q8YBONHSTmzHPJbe0UpPJHKxEn
gPEc+QxtN8tk1XYiKvvYp1Eo4AMpcuVsXkApeoVyyl3+YSZAJfwGQh9ecsXLF6sLI7dAWMSFYyeh
08BAvJCFaIqtG1B7LKO1WdjZOCN88BWILV6qokMZMOso9HELvOAJ0acebSOLG1k+ZK7Uz/M/Domc
RQpv0WetK5ynsF12+uzmVTW1I9VYZd/jlfVXM9Iex0EtlkHkyaNbE7UObp5A3OSFaOtJf3bVMpYt
7+egU2PINjEF/4igvovKOULUZkVwOzIVmr0zAGl2Z5D861gybE/egPtfOBZuLy7BVe/3PxvTxAgT
jw+zUPlQoAP5bxzlnKUyXUrezh1K3IHDHz8Osl0tV2E32Qe238XTbK/7PJTh+7ZCQePCI70vAXMm
RcQdziGofuWmBwjB9KadEfrAREe2jMnwLq9nXavMaGhlG24Q50k1EPw7l3hontU6Iiaz5u0scfwa
6KOcnKXFoA8pnr0K+qbSdFo5Q8/J+pvhhgcso3q5xWWiuqPP1C0eVGX8Dzd9y2OHY5JGv+NbLX6B
mzxuw9L18XbrjXHP5NoBaQMom0EfxYSXBnD/voi/PB1M1guRjA8Kqw01ZDtSesaOeMruFV7k2wGv
CJ1IH96TGAqLKLyY2jwJYh6YJxRgt4FAegaorEHasJXLXYwS8+Ps6SYVgQEsdE0MmNpag2T0F4OF
nuQYlbiptgl502Zg6YC+bnEf5+UjmYGTW9BEuZA8P9R4y1K4N7qRiein7p87OO88Qydoc3piVDJ6
iPK+uy4/+KCl6pZRIOkfIriQ0sxIy1oL8s+hETAatmLMhQlis0gEPQQWWdbYA+qzE2hG6cRXEF7t
lA08AOVRiBQFcLQUVrEMT6Rax8SfZwc6Gd+D+no6G0YSg9+XlJZs9WMxjsqI67Z1aJFjaEtQFDnz
99Lw61q/qCPt+KmDwZxj8QDO9LbKBMaLcTZk+CYRo9xo+t1b9YXDGvrZ8tAExN8vf/nxZt4vwQfg
+A80LKuTUCkpWKjcC8VhWHc7XLbsTw7OG9t1qnZZAKQv7IrtvQI0FPhYWzPveISmbOVltDhZuAqV
5PezcCCn2PTGrCFR0UsMeSIpoJjopjaUER7hmtyF6CcmkmOMh4xmuLn9Sht3lsvOh7nDn+uXb8C5
XB1/1WHmbf6wIW/JBvg4FuyV/4DwqErAZMufHVJLjnJZi1XEvjUka6aLZsgog4vmhAq8vj6wH4Ad
cbOUkxDote6JLodzLq6wFpJmFMK1uriiVZRVT6UmI87pm9Qh1wtIUI3LzevlZAbw4Gfz8Jzj0Nn1
7nvtcSBKNY0feKDadSCgmxFoG3BtJIg4At9ekIDHOTh7cBU4l2uPVoUd5BJq9w1K3DfD3vPamZPI
+zLUzY8qnFDECLVCj1ZYqxYoRDrCCddH3yNmmtONIPdLEJFkRlP9ttM9D1xov5BiyvngoYfMb/3s
HosS5Zq0qy8g3fk5pKIxMqqs7WRV7OAuruBTPjraG2i8rBf/vPvsjlDK8foNehST+gsH/d1+JPtL
U05KldO+4bI4OQFjnByziZaiJPbAqflxX1kyomlLrI3DfotaciSbooummAko4v8vXeN0NpPc3H6/
Czk1PNBjz6DHtkJlHSnlYXWbaamhOdOsm0W44NKu9vu/vc4Rbt8L7elpXUFV/CiJWIpAozsrKk02
WPMq7wDOuj5U4glFI/1+pWrIinSefgeXI9CNv86HkYxgLPzA9jZMIF0hmgys9bYdPNFEdXqsTnj2
CN5WyUdctt4fqZEOqeWTi3iNzP2qjWRS9TTa2v5Ave8nqs9ZMdiyz8VnL0ZOT5z6e8K06lH6wEbu
QF8+BPt2II5HX9SswtRqI2VBFeR6jSHYcIVsUIVSZyaL0fS2mhCNU4BeDWE/NTrf815xBYBjim+M
MCj3YMl7jfmoRtcKezZ6H1gvm/5uK6O22TMUExXa5d1QWB/KyvZTzTU+Wq2kVF3HVYwSE9lxHuAv
sM38N392Z25vcUcLZIijPXPMHXLdjiHungUTGjeP0tOwiCXXMZvqh9p62FAbg4kx3vZDRzvTawQ6
Yvt/K7xk4meHIPcP0Sj+niSNstT0Rc7EUJ3vJRD6yJIDZJmuomrNVMrZkOl8HH8YVNA5hxLI8E7i
thFjm50tQR8Egzq2g0JUTk5GVtX5JJkwQPgCxMRSsNM01iqhRxaz2xG82493RqbaZHx12KTwA1DU
DJztRkH73TS8mtDkcrAl3C3gnf2kSz57D/DkU3oMMVI/xLnslxqurd/7C8t1s9JvuVZgIV0/m6oZ
FEOxfqeD6UXDLq1lH1+EonAaXS6QASubEx87ANaxy9J3Kmuu5uzMsEq7R4hry5jleWjVcMm6UBsY
5rYyUk7IKQdbCrCuzMYapZUY+3YuE3k2VddcnKziHnQCykjRXqAX0O4F3f1zimMSIhq4wrSiYIeh
D0bgAse+ixMNn7rW5hTdd3GOjKCDZ1X50TuPYSRKaRs2wNUCUay6XpFgXBMAnk/wlrY+FlJfe5el
JKH3xcbk6j+z1MbLyOvN8iqaU+qJ80LCNm9lsJQx2yKiOZPTb4Hz1HZlpBelFjqCKuqCuIsXzuXu
GEYIZXox0GFXbeya4o4lIEj1Kk7SPMnJaBdAbvwCs1CHmn3k7QpsCUfau32+tC1M+MfTtSek7jxM
0Qz8CHLv1+9GfG3YY/NFUyCB/N0SHxHVM2lY0rqKnRd+DyfuGmk0qvRPdYpIQ8LhCjr3fSsewzTc
tWDJsG32IvPVjycw6h35/rivxfXK5oejboZKK4WqmQqmJ6PLK+IV/Fn6396BWD0j32J4kWakxPjJ
3UgtK3h5lfFqVWJGDIJHJa7TLwol8zkupipRUvNLAkFuSejO3hjD3MD3yYWP6brEvvgpxlY98zlg
g1rWhaKC4BcOpbXpldWaIs0brX9UzuqzIUI042gTBbv0h9YFg7Vli8whPsDslyXFxNiHa8CtEo/m
/h8I0u8SMNT7OQJ1sqhqUQQy/AIVzdi6WqDwbkIKqkavGTlsrRcjEnh5nRU6C3PVkdrGntTnGgBk
wPguBlQOqC2CIbNF8bkNrgJrjO+sufHyGXxz37A5AnTPuMk/mrHfvOtQt5zuwvPVwvoR+pm9ja1Q
+df7Z+IGrf6mTpeao0DVSF6EaTLJiURibhgq+ar6PPEoYxd1F25qNJgKIDeVwaVdaOoxm5vJlC71
ToBUbscnqAim7lxiuQtxWk7Vmb9D3UcZqJ/FoFEIXPFsdD1FUp634SmBC5HDBWD/YZ5o8RAChGQw
xj/Y2tmw4ZsBMBtQcatPC8KQRanPkTyELWto++hT3OFjckh5zxBRexgxX6ARWrrt/PzP+lxhFDZ6
Ezec9VWgOFB4Wybx3zgeZvyHdTBR0z1jy5QVro5Vi/6tnq9LKPDxCkJJDyIWjUbHo7NSVffk3uPm
4BNZgyv/QlEXS6P3sTrN9i1m3GgCQWAmlxg0/cWVEf2njYTy57uHARGUYaXFr2IgPv1/v/NsBV56
5troPLU6XDp1wYEVqazNgPl9u2LiqFk5fW0HvpYyzuitCnLBjBqUdYf3hYkAXB9oCzF6rJueLQzL
dnvWE3/LUhtYylCsbpyf47i5l0rDhuYNFZ2G+nxd31PT4EbCGMP1ZbJqeciGnzGrsAMp9qv/Prbj
9DZX9VF5NiA/8F8tAfxPwsR6XpBbuijIlXUGpKAlsbINxUNWE5kOnuyCIgbqxdObZ910+8knH/VL
QbZGPCMpQc6GlKJC3GKTa3khHecWD4GGQxBKjA0jeifQOVbG3by2jYjyT8rd5mrnd/PHRejx0irs
TJ60aR+gC50vyOz999qh1vfV5R5FMR9SJTA99EepbpxxAZcuTSA/w/951J9TGd3AFS7OQwvIE3vK
f6Xb2xI5A738pmbBBoGZUBbNJLf7c2dasVTIztvufYv4cbwjfzerotbA4lyjRk/Q4UXzvfxrbcA2
9ZRRpTupOkfRFRaqPgWZYgExik2LXQHR/QU2QBSwTO+DTciZTkkabhGqJyMVunQdwIJE6n2DD9uj
VqMy+WvbumYikNDWE+wCAgBfU4Rn+fZ3a1p3w8jbb1TkH/IvVqBqbGdUY4CnPm1nyz9DBxoWOE9/
fWp/mn50MoKf/ahn6Z56JAU5PHVg+TYeZ9OnOubLlo0izvZgMPTA8kaMN81usKO2kDJVRAMjRPKZ
tu58RiQ6dDvtACPeaNk8yJshh7HP9TBB+MMyQIJ2OwSCdC1Yuo9UIs8mFcvb0s22aqI5CHwljfOB
QaRoEH5a9i8t+njHJvLLLpljhPxxxQjXDTf1h2QBw+3AKoz96PAlYaC1kMyXnXD+bBmCFS7aqq6W
w2NoW30h4Gh8x1Ek0OPtrNRleLj/LYYT924LQbgqeLqIhMAoPSXw5KCOX2CzSrGIKB6Z682KiBqC
ar+NGY3BA19h+DudYuC0OKJ/0dij/y3vey9t7etFvQY8EB7y1/42neXB690nv0xxtahcTVT3AaMn
EMkU5H4D3+JI7MFmDOT3AxqE7sYi0sVY0a5nm8tP0JKu0Ma/wXMUGiyxmTexlKfTrrFIivI+q97h
2F9HvIB8HTShtKVL4P661TKK3+Js1j6obwfG0U0dINhrg1cLb5X8oCrp2jciEOnbl6aBI7L59iMw
p1aj/hPFqc5XBI5lVpqCdl3INyK/lgm5Gqlo9H6FeEN/eMR62NAmaLc+fJZ0yJr4o7BLnhQdkSJB
1bRankg8vGSHykgOYAFleFGlgDyuoDl5UsVRSx9MIYK45PBV4RB0nKaEm4ieX7XiPIEUrHPijFFr
E7kcH6OBB1O1La2yA4OM/1PMR8ACjNRPvKDVPx6I1EQjg1O/es0kEcvO6Bc5RBVqo4ACZZ4uKeEA
0Guheyw30mNsEbuZWmahAYdBLcg2IyKGgV2WwAJlwzTWz1sseoD69goCm39m3NK3JsSzqJOAFsRD
9CVkXenWVt86ySkpP4DYk1MICULciuXnhwDcTuGIFxjvyQ4+lqNxCiHbTL/CpoqaYtE2b1XVSJry
M85bLHx7vt64dKVBMxD6ujhhvKXFD4Vu/xCANiYiXe/jAo576r29Oqz7JKKdDotmf+8j+hoUmPto
eJDoqi215Rq3U1Do3zyQ+1pxKHMboloNrL/zCV6XQWGiPWcHvbeLaQe+xjcgiagzeV4hpheSUnf8
8J5HUzEtED262mo5TPVY53G3CYgDVNS67lbG1M7byQkNN6Picw3aUILUgdzg0RKr7xS/QXkqHZnK
Utp8mBh3+rY7LFpPaM9q/vafhTf7nObawf1oFyp0XrnSsFKcdQD+NfhijG/aQb9cJSJoUQfDWoKb
SyFqpYe2G+MgjE2Mi/sJPLLubXfPu3S/jiKP/IeOUPVlRHZs6gCQD8S2BJTrpBkBwr1ZiVQtVAg2
tu3mDFSVRCB93NqAQ+rH+vdnsw339BoxGj6cpkTXeGDgyzwta2KEZ9ZVEBBDHn9Bffynu5HdoJbg
enuloDPPZQHZiOyWsmStP8yV03YtreqIA8sbueQFmvMOApJXBNV3x+I95a+zkXhlRgd/xu0EXLCS
5OHtELaZ/Uwi7HPvO8DEJP4Mo0JSjqJIT9vMUeB3mFpz5pRaw9yArRSX+DzoiKDVCYAflApRaKrY
rCqZSBxzmq/1PStYW1c5rAV+URf5DZGiL76vyGPC2oUUBblhLuIpo9nWmaySsk1rMpE0DBRbasPg
AL5J13hgYy+g3fYyGVYNcShBixFBD4UQjVdbi0rZp2xX4ifxgf1xcUfa5aG9H0p51LgGu9hwpe9t
pqKR/Q+R6YDfgcO5BrdkoiDVVtW0TFzZIS94IAnJst2MqFPVEDdJd7BAfVuzWM+xTKJSw5Sj+tRv
Na76B0bve0enCGZN03TdxGXmV3ZbD73pxzibEgquzfP8t2vRpfjahOHY+1FMFFS31f/TnF6aJ5QW
9RrUC8NmLeRJvBURBJOKNtcTJB2CJr5rwL1xkLw/NbyerGIkBFVLuTOuo4hbipKRt6JK1xNNCT2n
NZlLJWt21OT8ACH0BCJL284nRcviVotTDYIO4uiRR6tpUiq0ZaERIZkNsXC/rG5EcYCf4RT7xCAN
iX87FJrWZu9NHMZAxkwXcr91qTF2nz3KpiaKEsWbHrjQEsYmRKWdPwiInC6Ni6lk+A/nBX07zBUn
//dGmnmUGlf90ymALpRxo/kfejsT/3esp+Q6iZau32gYop5D/Ftf7bkOa+Gnz3GkWKvfrVCK9XAC
9bS4o8d9cheSgNRNZzeZOndw2UgM8c22226Ft7vVzQOJmBP2vm2TBidzXHzsbpKy5VVn3CM3jYX3
fxI/mtrg9VAQYz9GwRo8+s7a8FByRmFKE/B7rJfZsAbaPJgrkyoPSzJv8n0BQx2MS63QMcfJbJLl
YZ4GMCgZEwl0X6/PWloWe9SzMT7gR61c4QP633SdUABtZ7x+71vLmmc5e+2d9u/Bo4D3li0g7hbA
qzh/fHtdEk/QUaSIuF/6bMs26fRsRim4dE5RJaQZ0hSjEIL6r+6ZSgJjI8C33CEwkbSzmfaClb2A
GRETgyE0Sl1CEOvw5+jtU68mJQ4EtnVjTrm/v65CbA3Ak4lJdTeZyNgJ9bGl/2+tDIB/DFHLC/cT
gD/8Hei2yJMvvPZ3GYFqFysTt/T2583egq7Gvk8uPMxDxB14H6MBu1etGNHEs4dbiMKVyGZff2R+
AD9JhPkKUytC0Pp7L7hrL+X7Qim5XbgUKiRjfUbVVX47pMkhdWI3TzVIitcnGkMa/1Q8aJQJspdA
lA/XGvJUHLMHJKF2GdwPmUAlezF4hT8I/hvgXbpAniYEvJCuAN1Wn6QsFPOY2hG4UPgSRmdegU44
HdkU1WzHXYaiPkePGvrvui+g5ByPoHDmMOyPibQQPzxQcnyXp0xjjUYlbtKNX03/sfnt+/eC0kzy
CIKc4YRCxkurQq4Z7dG8PhTA2YpNBy7rwvbS7BqNoLPeyk1M/nezw5RgWLqfVdRAN/AVx33idT+t
Z6LggKrDHfnqsOASD8nBT23q1jbqsbCrTF9Jub2I+qwK2UO+t3z//7ST3BTWRtcifk9mthwL/ziC
8QjyUWlvFDZBJ4jyW5MiXp19nH+wwrrDAJpUtKpMbwqYgDmKT5T7kdq0ifvGx7FwowME7hhPLabb
30eAWp9h5LO0DZOobbdj4dmBHCd+B6I8XO3smtPaGJQ3iTWCJCxy539O1O6t/SGB/5BC8xyymRiI
HFy/soM3u2YBDarCbT5TZ+1sPShiER3F2WTYcULSZEzLrItI9pAy4TCSAND3YAa9XjLd0ajyoK61
neM7n7nT9fb2qiMf1RSkHBoPQJsmdRjIjWW0XTj6AwxHgnVeJssXqKH4ACbM/OcTkJPezZK/71cT
bMrGbfNY9/7jltIqbhz+dqHH0fzRwIIQgsJ+NRgH5RaQVuq7TPU2dh6QqxCdqBSVeVLSZlKp7IvR
9H8HD6pye1DHKs95S+DkEXXMqZK8Z6MhtgdWV7EmgB3rJvcJP3HXgftwTsBv0LQTS5JqSfGHgqjb
i3aWXH0mpWNv4goGtc/VPV26tOSQZeqQRgtL5frqAi/miq5dgOky3hht5EPT6HznrQcqNxE3Eai1
7ikLP6UEURodSkLf7bh4kboODt6N/IGzdNy19i2D8mSH2tgO13u9jqEuo/KCHIFxMyWztdy48wNk
ODtXMjJoWWmIZ/crjqhWf7QagOYttfXnRGBUh1UY36OHIWs6OA0ZaS3ujUXyBeEZ11XAbgcQ5Sn8
nQvDzLLeybV1sPvZqAbkxJ+I3ytG045DiE6h9TPKfL5WdocxiK6LszGYvcf4jI7C7YM129gHaUS8
+DvkRWRYkZYPvOIKQf9acSXU5+9j7rDuKwaC6FL+w1zCGlLrplC1Y7YeItePPyqQCG/pfCaKimy4
U2GNdZynqwj2+5fzyVH1R6TEQTiWvobYBt96NWOkroe0cwGLfSCJVtjDzrbDKF7+K49UH37d1pYR
faWUFy0JwQVLaoPA/tmbhgkdprxiiKeRJatfc5UtNriG/WCf0kvjoIQFP//VUumv2PjATYprE0i7
Nm9YDaXvY1hifywuS1N5i1zjW/Ej8psZcQVeDNyOnDrfHsmgkTy5su4dY+0gvQTuFo286+S3PR40
l9ztlINn5NUH56Qhi6grpDfPD0zJK+Z+xxiX0OdAyl1uhq3wMSs0YZ/3x66a8SZABtEaEVSGIMOY
bsheBclryEgejSV+SnIhBGqUkchdNOFnY3kf61Dep64ZYsXnC6e+iHM1ZBV/FaCnpzaJg7Ef44Gl
EcGQgQr9CeCkNwyvk/SACx/LvcNnyYAPnexRBV2vdUTKmC2yhAQMxXYcujRjlRAezhP3IQiOZJQC
IW7laqt7/SM0qNdLpAjVUOLiq2y1t6MLEwhOJ2cqkyVazLrQ36KNmQue9oDpkSD5jTzlxf8jLoLX
yDYO/2zsjzVtnFIC7+E5/z/OoxP23YygQth4FvRQgi331SeEl2WuCIFFEWgZNLaXPph9VMYqR6kP
3wEXzR3sGaqgHANRv854QcTV5sXAfpM9EMGma+L2xWVxQjYHyGyHjX93OBp/tvkSDIwTQcl2gK03
f2IxswPPB63IfsFyDr+Qn0ukgkiJu7xqZVMwtzQz9WyY4EMUZ7Dsc470J3T/cJxYejr9BPH2Xujh
+RsK/+/AembPIMvpGbC/1Ldh9eeqgu0SZb8TaOiwlksV3e2HcK2GaaTH3Qj11AHZXBKtNS5ajuuW
B89W/V2XeBt4MY+7IaMJ+lcIdGBWvLGId4jZ3yFvkFvIJVYWy6zje2VaFgEoBIgDXWdcArnp7uD3
F4kKUs1FqkephZobWggr4bbU0ldhZEE9JFv1p4lw86VFrd6g632G3lUMGB0fKVx9BM4afzJzG/NO
a++IoKq5CDEr8IEul66+0iLQm52kWNQ/5fKdaHe0OwiC2ALzJytG28QbG1cwf5pZifwiYCU8SqaD
21bA2MyWioErtrStw3a5r3hZUj42OFIlCRA2jAZBiBr6bIIEUiWD+nF7rUslgmiweZBXhcKG1n72
uxQt/bJDIhNiYsW3zLSZ4SVG1fR/xf5TFydgifp9ntHZi+Ph/hIw4xYyw1mlbLxpJPOZdo3q1CZQ
oNqVcMOv8PMAM5a8SNPrOsmucnk0xjFPHfnu01fr4clzZH6urNIDCov4QGVUD2Dq/EMnE73kDsfr
/dWBbr32Sr5HFHvAQZYzF/4uSgMwlYq/dnSiUG7+4HpYpi3F+Zjvb3j+Ii46KGOen9n0Qa39qcQl
a1Qn+t0z5dGSBcRCBm8YGiK1qJr439G8vmLtv5tGlBG3XN/ivkocVWdB0eJ6ZCnEsUCTF7DmTkJo
XHvmbSEGnyp5VLynMjJGK9VeUThKrO6IekjMiKUyhZm7YeuvGtTdfyeTEyK9J01bVdYFBlbOOzYD
9Gw85sn3WrSNcvwySTPZSaI+tvRRC1tnnzhFUZVLqLpVA9Vb5EnN1v2K/pqn9K8+ulM8Dt5TWis4
f039IjPBFb514l893TBFOx7S+jkSDU1TWi3IPwgQlY6iOBCnBmTpVXIB4JsoSrJm7nOnIRJSru27
bo1Ky4dx2fuHiTmJQ11WnGk66JXOZiSfFJNSSE+CxiktLeKaa6jWOG2XBsS/TGtWjNQCEcQbGK0X
KrTwlGcV11kJA0C405NSRfBibsBYfi6sDCrxqJO+0FOH7lZLUQBAvuUJauEmbMoKioxhP8X1MEe1
ypeVHG1J8W+MmgeM5oyBMKF++E+G4DBxWFN+5F4vLFIkYtfr5XTaiVmH/8x6R++niNi5M8V2WPMR
zsIQFiufNxUsS3wzN8zv8/gS1Q5kAObHqzfayCmhEWKXu6RcedWodR7UIZVT63LyWkiB/rVsI1zT
DwFUjnGYIcYmWIadbqJmu+OhhHnROi9Fhk+t94Aymbp1Z79+76hny0g1HVwC/RyReYFd+TZcLiaS
1RD3BQtyKelW2d+PsjhiuOmrEoKaM4VwCfgV39QmMBKN9XLnrffcAxk73p4ZgqZ8p7jeIHBFaYdD
yXTGG7bxwiSi9tO09LkONkSkADK69CNb0TM4XOgQSWHbez6jXEjhntv5vrRllJKVy+JTtDcjty48
wJbmpKWiUF1oQYfnu4Pja6/W1l7Aq0vLivwqLMtqYiRu7vOHrZjykbDA4GzPfG3e5RDdpWprRhkm
IXdIX47treUfJfyWDzIe7gqPtbhwWeDkBdRbyWEYwvWYNWs0M5GyFCHQYvi7NnnqEEMrv0DoHMFw
dgHePzQedjh26ethx2Kqo91ZzcBftqC3UpHktpfvGwWPT+es4D01U4QT7yDgJ0CU4u+FwfsuKJZi
ePSx2dVHsBP4HqHgns39DF9fbvn49LfSE7+HiW/fEwCbncnFt7jzOCEAj4mhirofKo3iptZC96ge
zyq2YpWe57iSFzEq166zprsLKwjUiIAFc+yP56wYvimOcWdzqLVeaCA08vdtS3d11g4l8OwZ3BRp
TfWNeifBa6T4ziLKCD07+dZr3SKFSUwhBbGk8CHxBui8gkKk2uJI78NDpi4rvEWzqjF7CnLIJJNH
gTOrlhdAB8DNPxyMjPfexgaGp1DgpP+DgPh/TjBEc9ydxOzIy31UaNSaP1dQ0fCyEhtXOpMtOcaK
I0KE1d3RRFNXcH7Ct50+sjI8uKvBuruvAVr2fDL4M4/iRB1m+Aozcup5eOiyU4QrhnzXdLOuP7HM
n5iGioydzkBydHWFDAokLbgePtKgQtFIcbRXIMUTkWBfEVNJHf4ztUyHzcDcS5BEQYBmkx37JA4l
W3DzB+/5TJo0GuT1tY4N73GZ0gvAS5ZPf+tWzU+yHnBezGQ9xULft26PVDqfqT4dVTR4YeHIj9pa
ELXfYgPS7CNWkeBdn2LLRhN+ZnPaHkf7h4+2TrKlsR8ExIJGDqnw7IZvlGQtIEDHwEMdr7j5ics2
0OSnnS186qKW7o2I/fLNgutAKw4Yo/bhk5u079c1cvwYFp4xc9BtxSVF44AT2JP6M+1TjfaJnk+X
yg5njtjbLksomPcl9/LHor2txALOWv2eisc84dkuwZzdiSjFTVxKFd/D5qFS8bUym7kt4Pz9bWUK
YHLXHgNKc5JrpiXl5UOzZ/z/uMAmTqvqvXuCJVWLiZwiwP/YBxxlxpJvGOj0+u1bXUxJzpawZ4Dd
n1gZbzGP1B8AXo+0Trxq6E46LY9t2lcFF2zSq0dqwMYGNyaKNqMTC2lHMfwt1PQBhvXBzZHYbaSc
XijzN2MAZ8ZO3K89MO4ZqngVoDMKXHdwtOLeNyAkKHJo6RL5NinUS8kRFcdprI0PXQfNVruR1a1m
/96F7CKYUn0Dvjv2e+y+mp7ykz4BBOJH9oLqKwHAEHxb98vq/+Q0NPKL+HNcpjK3sDCAAmn6FXp8
LKlGIjvN8NhXGfNRQcObs+j1NVlgaI5Bu4hlQ4ptlT97PmLxw5eIBqQxAQUGPfLw1hFnOo4LD9/Y
ijYRHLTZcuY2DHLpu1qHWpZrmFke8A9YwUvqNvBFaz1WKOZEOzrREKCtnYmPtUjF0b69LkZB9Rj5
MOb/sXuxFYQwW1EI7Wzt2tMMyIUDKYfXYSt/53CAeFL3a632J+Rt/r4HQjKep58EtybEo9uGrK2K
RrkwYMuYiBrPVB1B7VMDPYeYLvyildeF4moI2srE3XTMJoQPiJ08+9/P1dghTHcHWS9Rc0TgdTcI
uyF1u80xgXggqig74H3urVbuzd3wcbDwmdj6GjDCimvc3Dgh4KZEEk6ZWAJobnlSsW28yIaRjV1Y
AnC2ceRAYCJeo6obZj2uyuBkfiQmcASVsnwdnn5mKGvt4hCJfaC5io875b8oTq9sB8Ewbo1piKMM
WCtm5VPprGU2vj10so0lzpSfXgfUqXMeQPEAZ5dWfihIm04bltp4YiAXDflzdTfdSsPQD5PRieKs
q7Q0oPHKw8FfaTTKostJ8fikXJAfGFajX3g9vIFNUymatyDzYxvEgyYgjUTHM4FNikxDjHgCB7ho
mVfeToVLF06mGKU5xP2tpYAodZRaGAIiD3RlhTiUOZ5fsNSu5YTI8wwL+MunhAJLE2X33UiTbFmc
/5vr7xo06cp94nKhm+ymESxbsgsHK7oV552qpYGxYzs6aP3kJ7laMlviqK1szR+m2Nfp80Oc/TO2
6JJT/dRJPVjih6bt+9npoDvyxaOcm9osJddAQkn9VVv9hGUQpJ4n5vM4j5sYPsyDcKG8A9vlrImD
7/GiNclSSqCx2JMwxOuk0PXm7Qyc3zuqATnLLOgWxQJ5VgI+B5xo8RJOA3TOV8AauVMaRrhh+EDo
+2F7ZNPiZA1xO9I6QTZZoqLyq0H3Khi5Iq4BhcnJpY76fFqy1ln+DD2kjLkgglOo9Tpp75GPmigq
9NtQSvbY+7Si5phRTvUGo8TB3071PQmbOQJB2Lco5LHPMjCRds0Lp8ynK3roV4QG8gnD4qFPJeUG
p7hM7TcOojMVXJlb97CmAx9swHLwNR3rycu414sR7UIvXXil1gEUUCMkSxe6XQzTZ2g4mw2Nb0K8
O5h0cLKa5YRjtLCmiBxuEWDblN01vRlh3shSLJzJXZy13R2rXmabbynIbslnCwogFdeVugQmtSq4
gQuzZm4U9UhuW6DFky/nwf9UD6HhHCKDVCiYOVi3VrX7IXxl396jQDBa/I265c2aJle+a9rmvB6/
FwrvzW3WSF7qFmdeJ9+ZhzaJQc8lXJkiiceSmWi9Q1bYolOmBFoWGQVu72HY8VcoJNlaXLmg041Y
E+OIBtrnnJnnD2gVlJg6l+kA5zGK9XLsAJLlwnYTs694dKn5fuyQuQNJngXCTY0qOqUrKjNTi7JW
T6jVbXu5xpuOgob047IAX/M0Gvfq7lUMDAmsuEKOkU+j73PHttA6P25Rrk/BZ36HITF551zx2PDU
drYHHlzzIKC/fkWzOEq3/h/CN+O3dX6hosfnNFyXtXZTlN9h+ZkX8oU9KXVy8VhNmvSuCtQhoK/7
yMZ08/rKrjHtqB/PjbzDNspz01zNYf9v/pqjMCOAmW65Kk0kdgtX3pNNhGtOwDcqPPr3V0cGz/GF
1CgzgQlxrXgWUrUPXOqNVW1oBreC5xsmxckzUaDpXw5RFXZFk/J4HNC2LfGj+zLs9eF5jQo9fiEJ
IZ9hBKx5wVhXI0xMz921xiG9FwITe2Nq9glOH+GATiUWsjjlwWPHFKk14L1xZOB7lK0hGZS8Z1tZ
ITpIsgy1CDjFhUYNXJvw76ty06W4EbSDpj+FGMgXaaQoFtafUx7KmZJ9rxEdTtK/UgQAPDXXAyIn
14bIxPrLM7/Tp/ko1x5Mqi9MWfQgsYW0BBoWuVlQO87d6hK9QFx9wpxuyJNKlGZR6jMu/Vh58Qm6
nAUVVeLiXQ8ptrwuxSyP+J4SsP+0VCcFPgWB5LsdLi0LxZvgiQKQ1CVZsWrBxjlOu6wkINr4jDLq
IzEHDR8lMNpr+/SWygy1YiRpXAKZPN+sksfVpnM+DnKSMSZJhJ8j9FU81bCmoN+VmLsGg8atpLZx
T+0vG4DFFBc3pfYsG8a8n1xCEnlykAa591qw5YrUlXsnCbJL1CI6ytygbiI+mZf+rOCpH6Fgo3Tq
Jg2yZfdOUdUHlWGJV0icmDWsmmvyg3MceqqYUJ48KoUCx6EbUFZQwgcR5Essuar6KsM5MLqgujJP
zbI5kZGrSbG4xyCoFiCELMkjXAuNJ0/GFDYGedaVv+EuxgeYyLPMk36Tc6Je13p8AwtQD3UTgJKp
Zk5dahOLr6ypk5atC7SvOpk8DYvTrWJ58iXdIUl9ypDVDdJaOGHSm1Xm+kL8hRhyMmKoAstg1+BP
cBXolJolgUhkIx53aDybzFfTafW5JMH2gluzWd+n7yV6x7XOnTDBLlaFeMd2OcmWzvQwVMQ6yWgJ
9hnl0o/HJeFvR/vbCf9sg9ZndWBY0bYWZ+MEYOPFo6ZC49bboGTiHnBwp5sFO7PIz7aOBnrWWMMh
RPDI3YHCaRimRnyKtJ9ZY14EXPOM5dJ9Qe9Q9c3lDN+p1I4W8xiFIrlMK/MO57YGsT9w1F5wcMrC
Pc47gsuD9fXWrxogprG4z6nLh6/CG67wkZ/ffJLmbZpH5FdKn6Im+6ck4GLlfFO4CL0xoBT8k/JO
xB405IZ5P2UL3u/7q+si6KWIqGC/yfPREvAv3REWZB7+P0jx9bekqo91Tg12t68lU5G1UqdQOzcZ
W5hd9n8bsgoepRDMgkC4vE5+GewmUEHT/ARMl7nJKLjaSvjAt8LtWLqPxLbDLqpSzfoxH374Lc5S
IC1oI8kqCEZhavhS5I81gES9iC/tnVfEY63FCpXuKR3QpP11PdQmKA8OdAMWqkTc3OSeSt+1JkUv
Vtv3P1Y58ScCLLiINKeztEHEbNMYRPG6BopLa+/aYgCjxYs9YFZg2XXmqNoGsG16qDFj+1pWrWO5
+Qp5BxjSlWTlyeW4GTnmW01Mwj7nI63uq7Dv2g1hTYrAFHgwjpj0MKvs57gbpF8gfoYO5/d05QVN
1hQqyZLQv5kO3N+1mDMRd1BmD7J7FYpu93rkC6toHVpYiY65xcthNbI4hsTJgwiFvN4glk5nqg5J
xGg35ERmx0CTVjeCewys9umlxDo305whtft1x+hSMEvgULTFJjMIFt3jiU0SjNQ1JMjaSmviWSUm
Dbb9TXgxDqqAihmr1EF1er3Him1UCVonCKUlAzpcrUZGf3WqpiFFHeeYX438ooTL8nyZD4a7AVj+
/iJhaAati71WGus070VBEwUobpg6PBEbeKP1yOy+qMHc1qvwhHGPoEpW9iT/Dt3GSRwAJRFavfBR
3Du9O0ox5peTNWHIekHLGEm0uApg0SE/GiCh8FLl8wRjhCCA3/ZMIgLTJ3h6v/6jpWIklYMtgih8
yi0VAiWhcELZw7MG3Gc34k2DyZyUFkZUajvBwQTrRpxGDre6PB8rb4KnV5NmGQ75EVlg3E7eeNEa
t28EEJXKhueE/Qob+qo/SJDGAzT8Bb5EdPgABgL+nDngYpB6uUyCNX+/yQk5wCEWOuXcEtfn19iY
jsT1zFJXfXKUWF7p2TN1NZVkv6tj9zJQGWMF5PF+0jKT1l8jSZ5NJujlZSF9RlJJO/JnOLEzD8W8
8CWxAQuMsidTitXTdlqMHx975U+i7Bn3GrzjoaaxT9H/yRJdDA2lXUWnzHotrUyU995UEDk94uBY
kcZa8Tvzfn08Fk+SjKDNGuIGYUs2oTVlapjJobfwEI8K8WNd4F412PDgbk4czUbCKKIbZkoD52Eq
e140HedsBzVoX+lKdRTkZN+JgvGdlnpQxqV+OdHxAl9XYMq7ml0I2zc9h3hjhYkJd+XFkDQXoo48
vf+a2W6eGrVpMOJAkCe6nbxrSS4dYls055Rv/zDYrdVz1FUgm/+yvLALwj2FNc6HpBjg0I/hgdFS
rsevuScNYO7ar0OT+sE7Sip3T5xQOWSesFMt5Ss3s4126wF4wxTOLNFRH4169U00aiaWvz2zzVKb
j32IM1RXCIszNIPHvaDg1hCuCfesEaIk99xk7A7j0BxqDTJhypc+zUJcCGpytFbDXzBkP4jgNDOJ
yQNLI4JY+LfJsvSUjhpLOdogbxcJrW6kW+KQC8DiMhOBn2yvJehY4cwdXEwkiyiNMAMxL8zLL/5E
IHuGvqrF6pnTXK8g32qbR7QHO5t798Ka1jbYJ1gzPw86DdSS00/Tv+XsTO3dkSqG4IfqRwIFV2Ut
qjGxAYmoCh3y/8vkJLooMqL6e5xQZexuFdFlmT+Rf4bdofPvKUy7gx6uw+zx6JRpgvM1i6GM3Q/o
1iAhWe1gnCZLg8i8ALdOTCl42dfyStBlpqoYyPMa1/hrc9f4PgnT+eK86VaeWCB0W1ZVL7U+5UgV
hKwp83usKrwyt7Edn34x+qNCUb0OsNf7IlT2vZwdC0bONHGWPH5h5ZuzRK5NPh33Q9KY3znqSMtw
RY50OAgted3FKvBGHjVx+hikFF4pnevq08S9BeJLfHfSCj9H5k95nc9FNox7LBPQgDMpT8DsMCd9
i9ETZuqbDeuNuztBSG6zFsm0espMyirslnEZwXnYqYqRg9Nflli4OgR7oRvxvmApwqnnc03tenov
bQ+qeZ8aZXiVtykrRmuMi6Ie5xukDSTnxrYVwGJO8mJxl+OnbgE36rPFxU7p7jOZGi0cEZC1dIFk
T1W532n1qJVsci48akVKNCl2v+Un75dB2ELtCArjDl3Sjd7rg1rZ6GjAa1hyqsGbHl68iVkbGJSY
pVoJKDAX8N4m2HYGppc6g145szAa3OmJ8Qum13IMrX982dfUzQKIymBC2TIhXnNDA5LWzHfEqjmN
U0EARi51lFHxiiORi3SFTKtqfDaxRxaZQgPNi9xqVoDN6VwvZcPOaWepEpaS+TOv30PxpZUja2AZ
KWvYMjebTjNjr1ECnpg3EAAkxB/BhSXd6Kqt2XvDTnEite6CURs25LkB2NK7gNNbnpD10ecb2FwW
Xfi68ad1B4S/AvW+yGnwsGW/FOA7cjJ6CR7NWAq566SPSef7xM/j+OEm6obzULKuLgxls07MPT96
PRAy8NOphsba+oXV9DRIbU+Hz+n33KvdPDIoz5z0Cy8CbW/Q4tIUq73xYtE2kjTTnE75drIBPTn4
UYcBOaX3wnFrIsf5JhLfxGTufW2cp55NevJDrzM9WozDRszcsnxpgiOJHarkM/zPTfDpsmd4FS7V
wO+wfavBfqoaj3U39wTLZWgsPyrUOgn/f08v/X2rIj4dr3UC90hPJzSEz89dFQIV7eLjBQZ+GRtn
5YOBykjM1ZklXDITv33ofzKXrImwnWqEI7b2q+g5Bmea3GxOuF9Vx3V3sJDzwzyD4iIjIEhd8kR0
wAC1jc+Lk5SgIDRLSMYZdFR1eLccsZk0wjKMI/AJh0JmC0cPSnKc9DmJ7rWCjm21SK8FC/HsJLYe
/DuGD1SiY0LXs8In9CANBDHZ4dE1HV6R4kOwHgTN3Nyb+n5r+f+QS4/sJKBBRaRH9LQTnXdfQs2s
+qzrDjIiHljNkb/jnOBqGDwbaqUABwYg77bqpfSRws6XKjVmY9Ty2SjI8XyyedLzSxMy0uWTP0VP
vnpNmrmHqj4zOAsVZqvW28O3jN2YQIRLS5WvA6H7HRzVKEuicCGRBmvsOX7zxZX3HSAXy5kYFzTJ
ZH6lv0mnKQsI8ws/spTN1wLYZe+wOYTiYbsExUsdeHcS9JJ68E4AMVAZ1RFB3Qzkb8yskpNQHHml
89H5EBjc6WShaoGzNiZIZRexEU67ag5+ix1o0fCBogQOYCq/EjICWDEzlrDT98l5Eew0PWsRbPRP
zCNE47QKIOtRhlo4/qjORCr6TA2zCddFcIbqn2CHAbkoDFeNH1BlUGyJ8c7J6lJIld/rd2FIcUEE
IsnnAK9Poc1QfHeCp/AF4v/QZwJbTyVzCLPLzDZ0NdrwC0bpUDaV3xjvPjOhdlZzZfSL1AP7+ZSl
AvHM7ib34+6svX9ok0ke2IDgo5ING70etBLcJE0wyVZUmXfRemT1spHvxoJ2V8zR15cwn3IrJNqD
yJyPOXXwV4cMmbnbdOBTF1hgpLYnF3PcTT30n0SZbChlfxF0TLJJm05DvtGbZHTCKC889Nswu6bH
jWxahd8sRuKNT/I/AOfYQw0p2MbP0WpSFOl46s8s7UJJenwh9hpbmIMFM87ZT3uoPh67R0K3atiN
u6Wl8LgjqOQcuVUypiTdyNGtg7OtoajUyaZtoOa+3C7z83uYdxuiLLWo9QQJx3CCmkdlc5eYPNQv
rjPbJw62rvUYK1K4/8Adw7EHRxhE0b93F+zGSb8xYTbMFNMbP+uQ5ZwzRukD9MWw4VByqN6xEJ/6
yEkuHbnTjBEg12CFMpVydm8Q2AkyhG/iPam9n7HpnwTcMebwxF3F7ji6/su7Qy2FQPq0klba0e7o
bG4pw1GRCdsg3sxbVsuzotIYUSTenilJjZzeGqFqySzBzQBzE2QvseB9SnXMqHCJGh2j1bgzgHfj
r6zd4WfrrQXHBFrmlmdfFTwMkEU2CDt1vt7p43Dyzn/DnoKCU+ZEhCrnURbuHZ8WIEElljV/FvfD
1tp9EUmhUQeEu2g52o6Yo7+r9WMpFHclaDrqTcbcxeBgfNiBdl9ereWyK6tL5V5bBmngcNomxjve
4jHctdn6J1otNlDWTZSxyIpOtF7DHS3hlkdRQBAGQ+TC1BOp2ki4slBMfAGMspn2Plc55Bf2qrIO
3WDunXkfaX9pN44CbsQ2/jdzLHWgIi353IH704iU7YzFZRE8JahVpUBDcV62OATKDlepts2tjKsL
2XJVLp5a1exuXIDs8u9qi3i8txgG4VDrbcSaxD55gldsq4BdxFIGlCjG2sKuHrMV9fgWzPbj4RoL
Tp3ugqdvfbCSxLJuQ/QSfyKEINcG9pAEzbp4MQRgYl+r5mPuAZcs4hxfVJ0M8e6ii4TVquaJAYsj
JlC8prxcsClLOJZqGQYh3Wl+XOOOYmbiY4lsBgSJKefKFRZDuWDVsttaDSPZIuk3N5DaGxZumfUq
BFjzgWRFBWxHcqJFqP8en4h/j7c4E3WD9PK08GTDXlwJop+qSD4gsckGDbZBS14irnySe6T+zD83
ifptrBYN+0SVjskZ4XQidIhWWocssu7YlxLzPpJ1h7MFWOd8z3f98/aUNUHP/ltPRdcaO6GpO6yf
SxlQnh/F5168aTaPAMu4ciWkJumKg8g5doxXpTQKbl/vJ2WB5DTG5IHOf/32aN22RcEmzokZm9Lb
JrKw2Z+MQIWq/vKHmqBx697mdugzeOdrM/XhftYO3BcZ+WV32scKtR4IM9aQmVrcr5DRL60guVUI
APO2QhjGTgSfVuDXIsjj27KUP99eOU3oScGp7Kn+m25X+RcJBLTQgZp66m5kkP1biv7rLVYAZuny
vRvaLdZaa4cd27kma+GEIz41fr/hyAlJMrDlk24wwhiFx089GzGk38U0fqDSOwTR4Dzbr+p+dwGq
AfUBgZhWW4WjQgHSqmDNf9pBpd1/elSu5kv0i4KSslKM3LNv5xhsg+/RkCB72nkMWP9A9NuGTl7a
VegIwlSZA55Br4DLcQ5R50Xis3Rwfu7xmH9MnHn+UMYtUOtWXFFNqXuFKEc6vA3hpoBLS+Ecv8t8
x89jK2ZOnbjehzKdhpnmgZZyoMCU1A/VQkTbVkENs+6fuNI/3+4ydyShjTWUdtgNIAPnE07oO3c7
+3ovaE/+4qmqqfe2wP5H4e0MWpFQA3lC/0WplKlWdKPd/aAT60UuwGO/Ehs93wgFcf0QmyVLUJ6d
aNTZXJwOS601o1JLSnO4POGlUZdVzUuVd12cI29l7wb9nM+se84ZJjcwj1eM5ZSZKf3nF9OXocQF
jIo98m331DczLOuaD1oeAOIZhLIrMndigf4mj3hlCp34LQsyPkaZAnqzyWqsxKsehM+JjdLQ+4Va
mSFBivsFdP4zU/Bwx2Dxqt9b4eTRGS1/rnqI3HsAor6/vHrJkjM/3HCveh9QkpxjlM8VznZloefx
QnBQ73UuqIZDUUOATkPbo+C/h57izUK0F4TvLAv517/93tZbM6IPgOqndIcoNpKet/k62Akgyi8U
eLiB6VYAefA/Q/QvOWsx1ldizsVbGdE+iHjKh61xEUXZNhJGIrAk6OIcEnDzXK7Ly6yaRa8KVU1C
LKUoEggShrWibj9sYgV6sukBGAf/OwuDiBD7bstbHIffMSDi0mm1/lb+12xlEDjuDVOvFDBXb6LG
xTBToXe0Qo1WgySm3xrzvZNyJtZhyXoxAmqQU74kGwLmIaOfMwW3mvuMCqpubQgwUnrJajh1Q909
9DoWwMHpvkVqkSZgy7n1dzZQCX5aXrQDfQdguGlNcC3voDjgFcl1uY+lwreG15s0u+JfwMMqvEfS
H4F1otARXTJxkW81yF/deR2fmgKxv7VvxtyGmddj7vBLOYU/FqktZ+c2oXgMc+9ryy+3F0voBgwf
Yb/OjUGJsGTxwZvFRPFWTtH/Ahf3a7lrC+rba48/M0tSzkSry4cmKVnVgK8mOc3XVYRsZ2D2NIcV
NL7cPJbeYpNNic4/11mK2SGYgcDCbRp5IfCy3cgPPtuUYgs/k+vezFVw4zzD6Evvv6SgzTg0Cu4d
5edP1x2pdwh7Y2rgoXklkIyDhPYBUJt1SdO/AAJzhUj3JmhsODmk8B8G5ghh2WhPBESmulxFC+UY
fAP8+qfwNl4B4SqqHc3CfINX+z2hi4b8POQvugRDoSJrp2ay+dDwFPuSsai7BD04XV4uGhz4DysO
DjvfMZUDqBNTk8mKt4ozSkcfiqyvzvjU3cpCCedhTMd9ESE0lJYJ3wqxSpb7Mq74TrnepXKemb+N
QmceYm7ZupdxgkgkrINKNiHPt1CU7rhR0aysxp6QyaZE9Fqt+7zVBMCVZgWb5T4+2ApYt2qC6F+P
SVI2lClDQ8zlaLEXEuKmCq6yM3aM8CeeWNqOBbNPQ/UNH0DC/aDfMGF5+JDR7yvdpnZCYqf/U7EC
0dDaHX/fLeLEPT50Dfu2N8e3c3SFdAvJgIhg9hsqq1Lkn5+p/JT6GcQw+Rf6PgrXns+RAzD2WpgO
i5oYuPMqG/DuYPUBMH8VMh/lsUSO84PGSNXhKxWtYQ7g3q79AFF4HTijmjCkNRgsnVUkq8bhfzXx
Z08tslNh2c4zIx5+dP/CWddiqUaJ8/NGHkVElrneF1knC2b1h2uAMyzpedp7MYtXdXVCPZ81tFFp
1QPWiT4R9pxMT/CrTQSD+ihMxwqG8+tSmsGWoJMf1SMVTr8jCGXSTG1hcdeZ5TWdyH4OtK0YU6IX
VYHL/5r8SR+0GPkmIDle4NDSYdcmxM0e+cO2ebBoyO1z8+0li9aut4U2jmOS+EWxWvHR1umIg5w0
u5O1jQbH2n4G1cRaNIskVuwfplQW4SNQkFkj0rGT/l76h3pQRtaBXfKhdgfvQK/1K6EZRHSBjiwe
rxbPrURd2dCOSstNGCPz55hGw6xrG9MELc6g6wdLLRP0IxkjrSJOVyBjdZ1pyVr5UkcURCUKeohA
4mD1+qeKibX9TU+6/P6YOD9zCc0MwXjJlrpGY618u2KFeFTTP2KM/1Efh6mC52x5TTC917c4LEEB
ojVPVRWemKuGK9sTeltO++jZDgnk5d+H90BFYm3BPtmyFTrB2i39Rq38FVH7YH2THVozC4ucAUKU
Wj0FNkXz54DSnadeRLLyNmP13h8OPEP/InDGwdge3zPVNf6UsZzFuth3NDLJgd36qExES+XQ2Bkr
Cfys/qTDMV3kRcsGtuC1klyOCPxuF0/YZZXF70Pq7GL0R1O7L3rxMy0/Av2FPqZ9D4BtsZ+rL7AI
Sho3Ox8eTDWulpIGhsA0L8OwYhzyVRpynvweg0rx6Qg18spj8OrwdnawzUOOm33ANnqKoIy86bDL
6IAPI96xeFn9ugAOtQbpuqTJSznfg8yV2jqAo0OHKgae8XUhG8f9DRvurZc1PwZ2y4Ae6G2y7C8X
hCMBDjyWy7L1aAGIc4dlRs1M1OIvIzhD8ZrXZp4UYLuHURHMtHp6OYLGg92nTLYEavmQUdSQpP4V
KwCEBwdWa+kATbCGf6Xo9a19fPk/iogBJC4lJajXmYwOUjM6LqvkYFWwhQ6MZF6AwUKiCW8vEqlQ
XN5viDzAwkHWku+XuXuxCfZRr4WMzJx9ch3D23M8ZgHDbEYl6hBmA5ZVIgKc3EXON8x0vuOLyjRX
1Xm9Hu3ooECrihd+HL7W3VWhVe+kS0GpNWrKZUsz81HXZHB8GM3TEp6rKO+AMm6F4OqBC+HfhbQb
pSlQhqlwKzATn9RYn96kZQHbIk+aSmaAInPhAScl8FiBQaxyEGATsbY7StgPUbbtqH/htl2nuk0W
V25Ty/THZBerWMXF3U8Iee6l9JaXQAFlW3sSVOdCN0eJ3m4k9jM/dkMP+npm5RbA6F6LAbbCo18J
SFX0zOLr/PRiwn7cHV2cY9HJFE0Sbsk1dRlXgPGnpF66NG34H6yNFBMmlfm+fDx2Fc/ifFct1cZC
7qF5dSo9HOaYk6XwtwJvv1SBinflc0w35WQq6rceLZtcRe1eWrT7he7X+a+yJqMOEgigNGa8jdDt
xKg1+z3LwTGiJ1Ve34F3HjEYMIz5ZINDAnbNV+7PhNO2looIR+ea59h2DUaRqw4CtbgstnAHZoRw
fXhmz2vpSSDLo8/HdOmX55Xm1GEC8G4THNjFTFPJPTrvXD87jxWaG2xdHhIeCV++n81V7YF2BXYu
oT+25HVRg03JO1cxscORjz5fifftVcVf4CFkauxIXLm+pH9Wxl3ZYFmI/6F4B1m/lg4AFNe7sMGE
sliL1pjYiOWFZNnHV4C2AJmsXNPSoMxgzokHJFXkaIuwNIHGv0YacK5tLcqYOy6C0VlrKvi4Tv9S
R/Z5S+l67GTM27mCsuMDoPlEV2boa6mx51zZLXsh9wnXZPok1kw5Dx/gSOqpgDUyTr58J6MF7HWS
oRo2K5vutl4oRJ7HQ5JL9KPFSwhrwQUgrifzo55dFpFodwoP5I00xfp7UO8Dmvz7073I6r7IO8CQ
7RICq2VB/qbZylwt20rEenEML81wnjYOrsjTt0/gM88EuDVjDE8hCVjqUeKXLAhdgxvrQbPb0G7k
Of2jV+bOHY4W8e7xmP+HjiPBkMQP8pZD/0GBJFnZvKeOYfQpea246OFh4V85po5EnYKLETuiQJEl
LDIJ6K84MwqOMhPCs8lLaWbXEQ6Gn3s7eZBORThqaJ4yEWnL4IvSwjp45f9NxoDLK8pz+u9Nd0yU
ZGcWG95cpRsZ+sPIuIqAp+6247XX08K9Gd1lclQIRN79RoeULSLQpLecUh4hIyUojcJG7uI5v72h
r+igdU90OI/k0N47y0rKzhG6ueGmtHZV+7kZy9KQMEija8viK17HG5uMT3kDPGUv+iYosfXL0JLr
uCdjgZVt2fPnKlb6XmcDYX7rYACjhuTdkeSo7my7TxsjNC9pSBr2CoR65JzW+N3FsZIzxwuvoe40
bsPJMvsDAKL956ZMRnSQUx/QQRRehhz05cmx8wyxN8bOTP81eHhrWjyQuIflFmAbL8o8iik52vfL
OMHzJyNo/NFT4yRe8LcydzxvfVdICTu1cdRc9FOMV8bblX8OxFTdazTJanAAk9hZyBLSbdQCq4+N
Z1dpskin9VNsIi1sb//5zEDYzezkWbmcMTOsQQb4MDFzbInFrSRn1r0uYI96hJvJiM77HNB+V6nb
M6EwRAO9TpDmsnFzenTTDFMGWcGHekLzkqO5iIsrcFIJNZbNw5txVlnI9vIIDx2mF8To+0lFVIek
c9E9YfNlsl0BSy3ShBwt1WkTRZLvugFwogBUMUVsdV75wlxgClUFGJgneeiEtkI7P7H9fa4vtOtS
mAEZ9RVFYmkTkzmPIwBGWA80aFlWsVI3IQCfPcOUAug9xGbW1mliQCdoaFG4NOkGU5TADT9ANPqf
p1rdvAU0LIRC0EMK17FGQN+35/gjFdvShKEc8vmfvHRkSV+Yz809r9o+oDnFpptKYbtWlTZAk4Nf
V+oSJKOtOA6f9SITG62e8bGWE2dtVGanB0gdXoXhtYcKfHCyxaf/MaC6cDCsZXyTWoYvYWUNkpNS
sdNEtiCRAH1bmfhSVL/tqMRqCG/1zbqrDAnwqiqYwelRIdMiCnr+avMHd6EAyYSPiiAczaV9VRhu
ZdQgOB9JVPvPGUpLyDTk+JuHK385S9GN/9mdVyQiyve0AwPwevNHUQPcYhzaG5ysJ1pf+uo84VAz
2FEJwgUMpyn0pwb60y13NlqiCA+2ZObjgCzjSx9H0CQP4x1MsuRjocCRvuxxd/tQVRQezsMcsDJd
zsTx/2tDOqIQMJczMGISvhQb841LHmNLT5uw/pfLKNiMOMvqv64uRwIWTtwqZlLOaeEa7lQe/MSz
7F1z1h/WeaP6KgwUBgXd7mZC51CFqWE0t3G7m3ySY6rHW9mW0hmAPslWUkTDO+jd53tQBaNzNfKW
UfAFdArXq192LjGerM0cud+2wRJOvrVeQpXA4G8GeF8PhZvTPzxLIVECLOChdQKYL18E3SkJhXAl
8L2tCMdSdq1tsAbRb21hQdUahb/wijCCntHs1EYzCg7mVqvN5O0/iIus+HS+sQjh6y9wVqpB7GFu
E0S2y+kVII97381LK9I5SLFtiXwyNcw8ggvJaHjMV+ke16JVu0WKjOEajtiwPL6WMj0HMr5BWEVY
eRM6hSWc1NENnrgWBNw91MGOrh8fDq5aDDy7VQQAlI2Zp6tn2Q4XE726T/ZXww6hYcePMWgfcoVd
RPQFG1YRJAC39T2pMy9GcUFo0pmcPXLAIB7WFN6fr6QWnzPn1su0NjPD9qK4UVu1C46K9QqFFASG
lPLp1DDQ664BF4gQ+Ba7JMxSQ7P30zo2ojCeuqW1gInNt53vebvZSmjT57HuqB+pZ9MdjGus6+qW
wpcTAsWuCC34Efbgji+o0KxGtfmKisZyhjQ+465ArUqEHNblChAzP8LbNWww9Zeu6Uwlft4SbBl+
/h5u16cLVD17kz7QL31EIo4pvA3WKL6xSlcGFs6ZHucFUuqKYPoGj8amOAFc/W1b0h+2mEIyhzuW
jkwKFxCaYuH94ai2/zUZKIJffYYbXVAjDPT9qYRdu5f53Izj+0FOuLuuAv473p0O7rzlzgaJCJdg
/Lj+R9/0a1BkjdJTfi6oLcYzL11KuyMUgGrq91BSehEaWDNp6YqIeO/Z4gT7PZvZxuyElcaPRd4h
HJRIhigsVN43NIel+oRRuCZea+bCPKEiZpQYzjEafqHvuu3A/luKGPz3Whs8999ALcSujqIactyq
u1Xo+l9CR7OvBJG34yqm/4Ihmthe+nMQ1gX7ysWtYTIp0+Fw8FfFY1lnI2lGooeJpgihB5LPef55
U78iWFu67nuHAnO7BVVraXF5xeA1hn0KyoR+ij2Z/P2X1czeBJt1M894rz06nDwwUIP+bROjCafC
Q53nVJ+IIniOAIqWnbBBHPCKUNX48hz1+pt+1C8x2jxIVI1QEJWG+6Jbp9JtJ/fSEk6Xhjj5t6BT
isrw41CXAMckviBsGs0OUuHyk/FFsiifomrLQva0nxtaU1rRojWIQBjwHnB1h/m1tkn+p5rIo4Z9
Ani4c1U+Gato6r29J/F9VZeGmHwQRGeTrG1uHZYP4U9TsaKMntOF63kjo4oDtFqYvkb37gJT5kBm
TJzHWOh55jtkPxX23Ht8/4VQlfPY1uxhczYvNvRq7CWvNyHO6gqzwOi5HuRQ5Tafm5rfm1HOC4GQ
q+d7M8dgGCMAc3vzPd2Jblia6yR/IdIENp6bsuN/tuT8dbI2bHIJ1gYgirSdeRSl5NNlvYM+N5jJ
dc/IAjYpK1ar1squUYDqTbuCBOC4Y6mZFyz/vP/rDNJRpy81yTSd7RtHZjJDVE9LsAPTtJ1684TT
8SG5VjUo2eNONogdS9lRfrkMC9Hm0d9bpUiYJS+/YHkQXfHDVqt/HsUz4xxJlc57yObITKfyKoCd
zSFfPcYJkqty2OYPRxzRWkNkkfD38nvHm8HhoJ8f7Daxb3owhY27Ky16504EvmBEB3GaZ+537el8
BZDLZGaH4RzeXqyAI3WSdUKrBEMRVKbe9DJe+/TycPqaMM2XUiO6iPjUxsEj/f48b29CdUf06Bcz
a5vjyfJcyWmBF7peIrtnKbLsTkUEAI+lKwd0d9XRsG4AO8d8QMxNIBkjPHjQsBCayFW1D6Q/i0kf
VRQ8nKLqzsNA1KT9kp+TxmXpyeZ8S6JmEDWMOnA52cFTdP1q8Jju8jIDVb3fkIqgV0YrAK6dCIBe
+4VG4mi9CiO8DuzPkFLPN2GtfZaJ3KeJ4QXV2PS/8sG+jWMWOS5qtmGLgcJtBunlC6Mo8diOso84
98Cc0stakXmBrN9eg8FSMZqYqbKBK8XiY/fdchrJw/huKvol1uUk/0pynYq3bt6h/l8S0A1XN6Rs
hb+woVomNYw08zJCXXGHL1zmF82qB8Ils8Y2ZmzroB5Z/fU2QIoOfUBoJed0eA2V2OwIXVDEyvQQ
Y/kEuV78RnXNltig/wnojAkG2r+0VrLhe/R6rhEsDw+WCnD+K5BqwaXJQcmmQInlU5rj3XuR55qJ
E/9+lp3gkNHwY17NeyqID0TQ3tAQEEbLSAi/OqeX99qzp+RjFGtt95M7lWMvla84tGvUYv8KKGv/
P+4SeM+Blp+O9rj0lQfu9Qtzj+NfV06uVZR5pTpuhKY7wilcQsr5M8qmRbYCr8DztfvoEuvMOuqW
2/MChxYdBM4Nze+lSevNJ7Gh/ioOm/iejbnTKeYGTI8IsS/e+U1MLnNbZzF72UHdIexvDNvxFQfx
cOw+jA7Mt55kyWkwGNxGJYcPk4gxX9CBomxs5cFPXpZa2ZVG9XjyK+bZnk6rViGVSuw3lsDruQ8m
vSXzp+X8muA4ScOYUlFoaaxk1ja7V7zqmeG6K0pJNlto7wxJ8yiyXMYDJXVm4WxSI8AN2VbYGItJ
2ZRhsPrqu+0XsfSkfc+TVDe/nSmOIYb5eMkvLIafePPg3qAmQuJ+5icM9y8oP5d8E7aSlF9UcwNr
d/DgPqyEGUsQHD896v7bbBB1E2jtLf5ytU40vm1kcT8eR/zZl8jJf7f6Rov1QQA5sRBQdTuiIKMK
1Z1QK3cMQ4W72RV6TrbM9tl4rP3lR/vW9sxXfpvtX/Vkibvs1aeV+R8xplARJTTVfVy7dTKAHr7F
MBgakOlVR8yJzunXVypCj7QBYbGe0q8GAfjesF1Ij8xnPxIEnc4X1xMIMsbskUlffzQp8QvmGkVz
uJYglIugQX9aDwCLGPI+JLWelKkNHZKvfFKtIQyCJndTVOPjKcuNH9U+TyMOeQkObgMMrJvsB6rN
qh4dbjusnTZCRmv/YV4dbqwto+o5ZBu1LTxKvoMHBjxTPcDRnsGL0MiPQRfFyLv14HhKL8VpsaGW
V9m6dBEC4rsiyvyHwK46I4M7E4nbfpc/vYJpEkecHxXYoZWz/il1DMxQfv+m0LSGkvTJwn+75PnV
p2Py3I3T4kJ0hgfFupbHrmv3SqMcwdeWJckTcMqQqiqNU3GE7H1bi86aaIzpb472gVjrEcwJbVzQ
bwW1HiYVDcPy6JgJzwxDS35+URIR2h4IyLgd0lVTJrqbHPLReONiZGtSS0A6BgNOwf094VfpoToG
890mhKpqhkKOo8zaU8NbaVhJd5/+lRhBZjDnq/anQ4M9iagTUds12oidOfIiZ1qEu1niMZK5bj7X
Ci7bRaLir0LI7TmJ/lXtiEkRTFkPswnhRZJMgkhnduxOYZMjGTcdtPT6TPop1nNzEK93ROS/FOkE
GDDwmNd7yiM0oO56NTHqv87z8GCewK7C+asBwxdUtJ5uiDN+jiBeWN9WrrQtRwEKMBEieMFXPoGT
WbS1cV4o3zcpnI2nbDoDN4QKefMvbkAEjtkbmXVjShp6WI1B7isalJ9XIqr8lU3NdF9jYDSP2dia
nmnZThSDwC7OLPdcz8jQVok1eZCnaq7mUAZBwQIgPyTm+gysI0d/SsxzZu0mEyFvxaBsb+UEBL4H
IiI7/BCVaEbgUaJxEPSzSsTGBVV5VScZSLfjkc0PlCVNKBEBAYoLjlF00XBa4n6YZ45MFoZxxwoA
VHnpSa96nGJYFCKcWh6qUVM6RO+KTG95sHjIqZT+gpfHfaUizBHB4xnfYUVTkMct9s27Lz5sfIWL
7x02DnuBFo1gNITAnibIicNB5kGNbT35zjWsr7A/MjOsqzOYwEQDp2S8qb+E0WhdGaKesSpIVWdH
WHLrIJAL6WZPNKb7VVeMFg6riH493MB8njtEnPNEtQFeoNOIeo1m2ItJsUcC50uyvdOv9Tx7G9Gq
k4kWdpWSy5VtFxnRZuLTAXNAVTtsly7rzpnHztz8OLrmlR9BBcSQ2YhsHMevQ9jFOrM9cMVzvgN8
je7FjOwAIX5CxPGT9hh65xsiGf5ZVTlsGx0G3LSOsBl82i4cvDR3pWSSIawNwOS42+os6JaaX0ql
afuQGlXtmeB/VAvPMOz3rSqKOg9V6vNYtDI7IVHxij5vznKCOgqbzKyvHLfdmZWi+wle3DDUzWyO
KIgoo8QurJoywpB593NPSV4NXPBYVUBg2b03wcQuVYIjN81Z22H9fCR2fHIkciFEp8tmHkfGm8rO
ewHBiq6FmLhzUf/0+kud8IfpgeetcTZTEmshJIW+gupDBB875AjcEmKoze+v/eJPf8XlqiKsVCC1
gbiO4cQB0gMcJ6Thk0EA5euY18Bf7ReFtI+APBMs3dKB89zlu56clNwN1eWDOuyldW7sSvNFGAVa
eei6WZlayDjNKO8Xgr9RjD2CE5ujx9kZ5gEzgmUaZ7Acf2rlGySohD7RTe9xJXRXw46mPHY6+T/R
8N/M3y+ny5O/JKqE9ezOKxl0eY8eeWu4uKB9pTFhCSKrNkVY97Au4C4BVPPeQ2kbC2flM57kO1UY
/szDbREDKf+9BFWJd+ylnWbe5L4el0iqhcCG8G9eii6ap07QwcD/35BWyBToOVibZt70aypGkeXk
9h59kA2+TT61ncMo94kWawWlwEEmq3bKjpgVImlHcgusuHJMpgQC/xAiCXhL/2jAGzmSIGHYAYXR
4C2IVBWa+GWBG+PRX01uh3WECOFva+UsRLckCyZwCHEUNvgV+nBjkj7RCA7bDFNALfYkVL4XyBod
1z8Ovm8QsCAqzeFrjhqqImstTGgjNpqCA9jlPd9c9cqQGrZYCrJlbPzNv+DLwyQpqQK3bGYjew+p
EAfuSZZjXwdBG2HtYsz/EEf1gOitjkJtgbQrXYQujtbRwe4yWskFTEGy7ohMmm2ATBxsxW4LWTAz
eBKMNp73gKyueMTV8l/2Go86OzdSJyJwDpjE6G3plKlLbPYmmECTsilyt3AoRf7ub6b07LI9BCla
c0cZ7lee2Gcl3KTZhFPLUC9WZSKE5l+ss/cML1pAA0E7m2xiO2p/6SAGGVQmbU9Z2oCBmj6AvTvC
IQzX+08fBFS7JeFr0az4LoVa/PA6yK2FExgGwjb7GYOm0GCPInzeukugfKbtHfKUFV+aNUdH6btI
Cnvthy7KKE6V0R+jJpYUP3FpR/3cNPKKjDc4JO/TC2oDltp9/wsxkAYNQSi98Vcc8M7U0CYUyhD1
x6JlmSxbZTZSkPlUV+g2ejvpEhoAmAEaMfJPvGKeZrl+9IRhjD9Wtr8M/pg+NrvXGBtJApeI5Lpu
5CL+c3nKDrDnPXgpf2H9TwfIcUJcc+ejy61nk5pUK7c9DyyLEcy890brxCwaiwzqSkK5RAktGwaG
aJ8X+OjkJTJ8OkpxHTSc+TdUnzxDoLcuFhTaMsTr1avjFE7jRX4G7KkJxJtfhSC/kQvMDlYdSj1F
5KYlPRVpsH1BLutW94mO+cdBfGbsTooZk3uLyF/09KMfpONiUtbzZXveqkKnQBnZuGrWBxenI/BR
UmR2sN0E1+3Oj7I5EnbDNYMDFTeymIgPh29F64W07QONpm38LfYBNrzwY9G3tj9CDQjR2NkoRkSP
QLjulUkl9iqulVfXrD3mP5bffHbCvTGw5yNV4C+/RM9UF0YSfSgvS3QyT1seG/zfBxjtB6cp4ker
QGXmELHMyZcgOYMHxhOYy5+Jo96Q7B2CqZCxRN0QZ2SVjYytZScMO4b8N5KWgiS/4XRbVfxPT5Yn
jwDvSBeNeqVB1vwj7dEyGsOfc2jfeJ42EcVfuARq0KP0LrY7PaMx07843A4Os9aQykfKnxpXYV2+
tosW29uiYTZ31Q1IU2U8QsBBSVZboTex3VLKyrZRYHCTO+7dxLF/3frRkX8kp2W+B7WMz2zJr8ig
Fr/HlzCvQjWH9hcNPgqLWBQoj1TskNxe/jbPC+qW8mjUhLEU6D8UtMGWUIrixuK2gvUWiTjl4VRD
Jd7O4/H6gFfB/6z/3fu746B2EyV5eSnQndmEU4NtQrNJ4SldWXVVAlH6MwHj6cPeO4U7Jrkdu6G3
2K0NKIb8XVxM8L+pdYWlbaWU4liKlvYvV9xFse2PSHTPCCInTJMzSfp5V5lzExPDc8miZBCIIilb
6EXGRj/eA6BkG4oZOB6M/hmTGI2N9BH5bifR3JwW7Y0eABu7BkZYDRBv60BGiyNpOVzs7DeNNd/o
NtogqLJptPaxUP12hqxMY7YuCU+wcLAXu6KcDJDE+Q+D94mVPvQTfE1XUtHT61youmtFIwoh2H8+
cYpuCwjeC66Cvi2cnZ8OL8QUrRYJTGqjVkpINBrC2h50axd7QeVv+aVM/+rhlwgEjGBdK84X9BWd
1fiUDV3xKBILeKGv1aCn/VUsWuGSwvQ9O1hjGIf4s8WemUzVvwmk8TtkDGpBOQ+H7hfdx+7bbp4J
BjY4gVCEoC1sDt9lnUTArYdB8rMMWmlr+ZvCZUtkDAU1Yaz+8wflBxdNLlkvNgcfmaatv+HQ0zwv
bLYRV6QrHubngaJvV6PPoh1MXAK3kMFiaZEs5kuUMVXyjQknbWEzqxHtiHI2Me2aeSMF4wWZGEN/
fkLJispnrSnl+ZihTt/vzqUudclMdXoxp7Lf8I2HGZb4XTV94ttX6DBIL/fKZpNUVB9kaleF7srj
tISKw4Bt2Ii/EOO7XJj0Lqj13cjlrOPeSo7d4jCbGfpBtOFH93Mv5g50lrlugE3f0u0bmMw/ilE5
MyqaK9BFl4NJYoBOMsQ18QY8n8dmWs2HyQqYYeteOVp/6n+dHBAy3wNq82i6THB9LduD668NOOv6
c1CfKpiqkZsPOQ2yBwvcYWEMce2xPXQRsgskkwWvHnUL5uUI+XLCRkf0e1Kx4aFJ8cWSpT+xkNFV
jyfiyw1Rtt9mSJVVegv6JHH58WTu/muKKu/J+xTg0n/uxAEUSvBHnxDQ4KXEpd44H1m0PygTFzHh
CfO9y0N+ZLsaSzmb73vXZMyNrxnID6m4KbkZ6Si5mHHKNVHl4dWvbNkcNSMovdczr47AQ5oo3YjD
BXLgYTH8ASGdKneCCCeMcz/0mCj9wLO+eb3G9+lBr582KTp9gNRaLoKxjCQxyp12S7i68Yuwmqyn
g9329ramIQAqE0J1wbrwXN7H8w8DK8ewU2aopUmCl6eK3StbvARXpp5y7afwqjrpweJa9IJTUvDA
nlqQYd6zrn3Q9lgmiP44o1uqy34RUXVNAnf2ppS81zZ3QHpZq23xKCy0VRLJDLxhH/PCV4GDtjTi
Wr5k93IWh4b7XtQ5JrRWGS823UJZLErlJ0Zj4GTxeGR+DZJIz4TTih4mBpipXXkuHvA+ikkljIFC
A0gqZUSYa8HpQMHsTX/i2Vg8N1YMnYqffmJMNp6qtxnOPZ23e+/T/BDkvYXD+mhsHLp+Kj2hmUGo
u+JD/S+MMkiGg5YM4ja7+CQObimyKcChOhtlahC2rHrSXHpVYJNpqvPu/+rzeU/B7bV8dR06dKNa
/AJ7GaGfaoN7xXkV4q9sJMXjRhV7vbqok4B/DKCyEKWbhWTY1Hl7B98twL+J3l4ASH1SlGsv0Z1X
QAkpd9PyZoV7z1Mpum3e/UMFdswmzHCqKQ/9Nwse1lOfdvpgYnYXw6jH0lX6Pw5UPN2k27VcttyE
IeEdEicFOwPr7Cb3F8PW/RId/rcGttaQ8em4pfFQlSvr20a8k2ZMM3cP6lh6O0fO1BhXgLb0xQ2N
odGvlOC0KTPtWwZmPvtlfpikJkufKsb0+vUaWYdBWPMlsQQF2Fda6tHS5lmPoNDXZD+mySIoY8Pf
PxdtJ80RMTEl9+xSKk3FQh8IHG3CUXDryuZxgmCZSmxv1WYkhFPZIS08lFOl3Y3iJ4KJ51sLjRWM
wZIxcQ+UPGYL2OPOzlrmC+sTs96pvfBMUMhhRGRl5fI1AZarhjBlWdHIAAbnkrtymKVg2ZRBgSpZ
DrpLmBbEKdkZZeki/X+TmoPCMpL6j8B21o/5TXzY7UV1COOzMNXcy+oVLtH1FXznU2Ve5EtgC1r+
QdVIN44omIeeA+EmZeuYTm59omhWYMMWrn4ARhT7F+D9zgEDm1gCRRizR49XuZWnWpCVeKKH6DVu
y5VZ3REetuZ6UzJVDeonhORK7woo+uJoUuNWChZqtdp8V8h+OwynV3L4GujbL9W562EJFIQodbH1
CtonrcWgVxa+2cPLj9/RLv+n6B1onERdcU/ssSnxqt6OSmW/Fmx20Jm42zzuh2mIa5H2DFFcbQii
te6jCXcYv3QfW7Ry2yEODytG/ebIlqqvj6PlQ37kxzMnlq7zvz+6veKH1J3Z20xdCPpsg7qU0RHJ
w69NZ0aeJweYM6fFLsu+9GQG7ffNVHNsFsWlDIDU1/up45azB8mTpZbizNPgIcZ0uJWM6OKTkkKj
cukj46awkcetM6suHLWFKWbsu8/wL4EwD+YIVWiAv4oK//O2GcIYglQT9m2bjq0M89uHg+WZqmAP
NaAobDbRVdSdJU/pWXArxMFUHuaYgpBBUnZTi62RQog4UPd46dbus+d3LGoyqhN1wnHRkmTvDWTu
SUSYYQxXeSutiUfwQzSwwqPt2MZvOyw6radJo7CCP3035nWTNjcKsVkxLn0CY9ujOI3BKnWvYgsZ
kLs2JaDbAJtBLlOv9UNEzef9cy5GB4g5XM6T4J/mk6yQFcM+G9mwC1jz+MhbQsEVtbpa5VpB+pWF
mon/2bgdD1XkeT0pBwv9x3VUH/oUta/y/Hl7ywKioZpBqW7HKTyRXLU1I02D5UhTx6myXHONbp6C
IZ+fhostaqo7PnD9Zjeen64lGylNkLYvCPCPix/cjuAqF8VQ0jUbmKGcs9FAwVEUultqUoMhmxcB
8Yr1f+kpxIZ9Voilp3ArjmZebMHCsjJ5s5coHiGcCxE5DshXake9fBoFHWFAs/hskZAsR9fRku5l
QWbHrgZ26JfRmqr18bZzLuC5CzzQ0Mteud+3R5Qv85kc8Tf1kt0BoxWyverOC9mK2JnS4TOY6dAe
/DUnV+/+zyMswu8bPKTKR/1xSVKwzoGvOa6D6tBInD1KrYfcj68o6Jav4of2dalE03rODn0l8Mdl
vHVmHJCjIjqtyqzhQnQIDHS9gK45moWeEd6rvxgqL46AYCphmeilQ8AimwgHUjnjTS6zYrWOIVBN
GPYRm80KQ0BhVvBz87kiFu8YmRn5FqGDk6JeCrZ3jF69bq7uNRQW3NgoGKzfrCZfs9TP/DFz2d7u
eqBhNfIxgHCFP/EBu9SVxwiFkrnZQI21c1hZAdaGTQ3OxJAeeshVnMs/b7JRrP8x0kvauMgc7w92
4aprLh/FW3rW+Tu1HkkYy2C6UG+gdKym7uZfYRbbygDFODtrpmFTV1oCo3+LAY1Ld0wX0+bGP/FU
BuAubelCWqFhVMM/BXovodDCiPi9AXiz7rKUUXF3yPVEGtC/Fu8f9cYQsSobcfwPl+Z3j7OHjFbA
MYfrOE11XQ3iEBOWi58Iop02bLwHYomlua+j+FNb0Cdfs0a3bih6xOXdU2RP0cFeLKZCtupdRISU
riVBDLlzpVAlKMP6DBs1LttNnZWF9gnRCzk+YQeFVdlzQPW+ZLC5MLep8D8RVwD88wlHCLL7cFEo
hI9w8bKPTbBLHNNaD+kMiXnL8cofDJZXVn1J5dYNHzOKyq0aBdtymT/MOQyDfIFS+Ei95XqeJ1SQ
mA/Jmh7sfF2DgMwAva/Ix6C1RUJhCGsGtYQI+bZCGbHsKPHocshw1tomXy6knl7s3v7gTusIDRF0
ivh6eA+jrBNu52YZc2ulC7tVDhES0hN9+5cJnqQ9+pCrf37/89IGKo83bf9NTEKobuLMTcBV7Qtp
bFHeJf0naM9KSWR6peifTJkKuwrSTGYKstvg2OjC25N+/+GtpvRnxLP1N6tnHoqV8GXPLqH4GNTM
/AVWwBFXbtpdGYIr8BjmUTMg4hgvKP9cYIqsSuPjqyGCZvbtwQJnF6hXJ4uCGq54C9Fwpkkb8kM+
1X6f/OFpXZbaHd9+Hk2GVbKLYRFFJ7/ePk4buOsI5nvkWdEomn7n7k3gCmnHIqSu+hly+H1MG11s
c/fZYZc3KLq2FQ2psmqP5BGmj+e72g6eH04LBH4VrT4riQilVWbJy0WWBFM0Kfs3LD12ncGxHk4i
/F1ZkHryhUXD28leaYke1wxlDNGuQD/AWNaOjWcYBD2fWf2/cG8HFqS/tKZJcE+Kw95F4vV8j1SO
tx94BWE4oR6bX1a2scsBcXU+RGTWXEsqxOMhvudADxzQEhv5djFVZonIR9cBnwCdxJ9Z++zOPj48
F/8U9WwfMV9cEqSjeIn8suzIR351lhX3/97JG1Siq39Cl7wazV2qgxk9MI2d6n0FyVLq5N4AQUR1
T/2liivx2cOfWoriOKICBYJbU+gZAEEdvdpUHyw8/datv1tZvQKDfxa7m6Jjain/kiVu2fsPNMGw
fudKM9ZLJw56c2vrZ8WRoGuu+xNnbcdLU4pCSRzh4gUYL3qxN1XdHsRZRHe0o9fKEyQjz+wRzkAm
ZzZPfHWvTPwLTJzDkdgwzDVNg2DNjFUeGl9vJ/Mw18ZuAZCWmF36I7HehV8OFjzMKJ/XJzdH3X5k
TiOJJUX/bbZWWqlrcthbhtS9+hxf6TjGYQEXyfQ0V8lm8YoSYsaimkIi7Rj4WivO2sL1p9TfpOgN
tvLmf/uPWIdGaWZ1Jk/43n3o7WxGAglTgOLnsFj0jizTFEXNDrraQ1w62UGobY9ZCl2Sxr0uj+qq
0qZIClJJP0bAOVwSlpZl+6+XKOsFut4wtw5/xczYZeyOIIRwNMztLWn3W2HcbTh4XJCiP8RePGpO
QJ6dAxafE6XnZHcJ111inkRzvtHMkEWP3t9RhLqq+oBgbZAXLq9XEPxFCs+v8rVvTmGcrldpsF1J
ctp54saaF5Ot4nSdUl0uEkilEGMwdyAv8PV1r45XGU/2ZAvFma+DtMPXhsZP7kLVH0z+7TXxOgpK
C6YVyTVSDg97DN7DehphWH7+ivaS9QYjtYy6F/wTtkyy3g2rZSnL6rs1htTiH9oIqwg9W34xauaJ
qhKhcM9hitOoemYm5C39qyrQ2ia/Z0Pf3G+Z3wxOQ2/1u3GSYnckCNhTA6bc58BToTg1MSrlYxvF
zqbf9jiYSLOkgELrkAgV5WbdbijtcljrkFVxxHRlP7VlQdW9A4DIO5hAwtZm9/aoyBokvfYYreFJ
WplaiFr4RIPm5GXxKgECXWyGPgxz/M6ooatV+/aaE73Xud4IIZgECdGVfRi6/GHUFSaPBHaeKXZL
0jwaPPvpj8I95DDXRFoF5yAToqQYmfUAA+JQuiTAyp9scyZMGsbT06suU5aKqwbxfybOUxUAcPtV
z74KvYeyTcYMDnfHH5cdC8hL/EnwnRQtJXGoUrRBH29VHikOOUIaGT2gFxk3o+uhUw4ciJRybpij
XIJGo6nosspdnRtgBpkEZRuVQhGqA7oOkOoRrI/TyEg1O1r7rEvO0mtBNHfwZjh4RF3Emr5Ggt8u
ePtkGzG/BuimlKYTa94EcTDXX6l+hWFRcvVwRyzSec78vFMZeAPmG2LodUiYv+T3ruhkKCKE2ki3
Tmk3h/pfaMPUF9BAazMJaDJSCMD1jWCE3V2nCL2QauiutTm/fvps+zslKT3/ZMDqFjzrP+YEsmqO
J8Ro2BdDuceJmAu+J+YjG4IMBxLWFKsLxyzKWP/9Sa28nLcq6LCzBXm6f7AyDcEm83v0xNQu8JUY
YM+cai7Zn9PO4XvMhuswKPIZp7TUfznHYECtWEGSTRsBqAhLvRDER5Th5gExplXKbAN5ik9Am/ol
XoUoh3S+6kRCy0M4gbYWgsrZmR5Gyz1A+3qRmIm7qQZKnHsUHC0Z9x+Th5h0KzcXn7I0eSO3tfEB
L47M5JUdw2HwNvjwv5TpLVBo1wEW5HZghz4DkPBYDyC63HHFJrSAgz0gC86BromT6QjSv1n7VYjD
fUjOu4RXMoeIV9qINNd/crLEBWThlkkAfu+3MP0VYBxbvC3CBki6JBEly5F303wG2zGX+hL7fEQG
+g8EG6qgS7foLSK+5S7PjbeSSQMv8kOzbdYqdT1DAV3FcHfQe3TQPRv90feAg+UOcdBZSxQN2XzS
sbnelImBsXpTI3Nb9Uxo0EtTjMw28ImzTHdKVOSlOTYlw11OYmjROUzIm3fEPXKiSNVi6zslt1Jv
e4gQYgjONSF6mfekVl3W34nJIAZiLMyjTKvDD57E+62OMvfRGGISQKLJmrW9vj2O/mx21j1TUGGv
lflax/hbQYWNx3453JoSpbOJmyD8a5MBx2ew3xxAgyZ/k7ykTKU1DQ9YdOl9x75C9IHd9NexGzYB
eCFU33MySX0l+F396i3LOTWe3Sw24Uc+1YUogbeM38TufExPIKvyLn88cZu8UwhJyN6exMc3nnUH
oDWjViV2A/bcMRj2NKGQv9oH7bJS4meqsDItM2txvOiik2FIF6zZ8dLZwnqS/Xger603oPL72ClI
uygIzjQout6ByGcBbow1zqjgwDdugh2QfzXAIxFeDOlFyH2Q102FGoyo7sJK5gyF32PAckp/elKS
NKMfVyNQizupXs7BsZG/GLvFecjLcQ/H79bL1IgMVwinT3KYtsBv8iQhLsWZUARWLIeethGkyomv
J3jmpYICfMK+o6qsC8qFzKRZpqq8Xe44+E6bf2IKaBrvvP52ACRnVOZKkH54Jxql1Bt5RPuOGgwS
A6Pt7Upps6NXoD/Kj7YtoRteWt5dHFvVW0KYgt+vIo4r7OjZjnl+XpqEPKtk/lIx9JfwCa1G/Ihd
GwmjL904XS9omCDha7zR/kZXKHOikILtVoQmWWEYa87yoTlZ+XEUFaB/nxorY4tiwrGzONRTllwN
dM9LKf1bRsU3w8daQj+yV2OPFAKpY+lO4M13QCOBOOGYGJX9OFJ6HO3ERVtTYigvvobJtvIXrYhh
JDrZXLXCIesuJtEgF63clSRMjzfjexHVmhauut1lj9w8smNcpjXWKq0rFXIfIs59XHy6+4IkiF3L
QikS+77s5pCnPCa6XgWc8rOWLoCivzjrsb4JKP0YpWl9nfVwnJ/hDb322vIPMhGeQ4NV5NnsaDov
WlqBvfAMmYAX1ScdSie4PZ1EzuS2fRlWo72+geHPFEaCIJc247XCy01/pIY/PepP2SfAAD1kdckP
41tVtd0TZLERp7aPQRPfu5V1VuQMAPKs9ZI94G+lZw6mbIw4O81lnikv0QDkb850rLIUWT91des2
WBnvuGdYem0YL1PWclj5TDs0N6A6TFdxe1xG8W4WVPVkocv+qHa5s/Dwd2G8wqOsxBKRp7CiswsD
6UymoZEkxXaXPSrAjNUmCUn5csG2+JMBkaRbaWhSHf4tJ78f/2q3+q8ku33DB6G3QmM4WHGNloVc
HxQsKQc7cR2HaJ172Z48kjC+A9Gff535gtc2qo8z+7sP1IRa4mdrG26hO8Hd0aS0PGnCtEV+GCUX
2ubdjxg8UP/dUVzknQrhSooYbp5F7DYZyew8T40Kc53ba8IMQoZnzYy2SzRICV9l/uUb6XUcpCMq
WlcjCqC0FS0yeMTjdYbGtXNUkqdk5j1NeWVj2nvJQBjyt+Kasq3Tifq9cDlvHHFOeTUVGhtNa1qZ
y6LhBM/gq0yAkh8OKHmDiqDpm/puz5HUoaXTq+EeRmerMqCJiejZrFVh+y53ibx3lUMxYczJUD5h
qAnUcEbvQiH+JtFeKBG48xyhc0Naey84aOCiB2hNvKK44xXwQksLF5S0VEcoq23XDx6yxAfyl42J
loknEKzTB3TsxiEHURPvjyCh1Yc2Bo6SwaOSLRVitJ70cOUTOi+kbGUuFjOye2ZAuB9KzaL3eElV
Ln7Lm3MJZGr6keCJK2lViM3S4zwIgp3qgUNS5IZH086mlGrOdWrzPqVckczrVCZ1yUP1OaqcOJpB
3Maz9whtQefYUyn6/SMGtQxN23EraQu3j1GdCXqUPrcT1n6Vw6DKsjOd4G46mgOEzJYP8OjDyz42
cVjixFmqzmn7NUeqqWasTBTqbfjhCsp6ycvgMT8Q6vMBDQJJzvbacXmgk5BHul/RQZmaCTXjW5hI
SsGoexLqpwRrbEkkcQNtq9OnopPHg1QOPROjm/xs9mliw35gH3GBK7giSrxzo7WgyYtJpsCmiySP
2PkYlSAU9uBz0ac07Jalf3z4+PZ7u4GHdj+dvLkRw8+lNbUDu2sk9y2nVi75fMHe4YpBd9UWVjlO
p1jxXFo68C8mVKZHy3rbqK4UrKcvEVDpaFcZGB+iaCMXBY5VRXmOPXgwZLi/7yQ577w7zjw10pqJ
NkhHsAFuigAej4jVnYeawmvI79vCBCscCQd6bSkUN3Rv9b4/y7+LF8Qf+Ivy5ADI06H+xA1WEYfd
OedixFBm52oiUeYdKivTSaYQWNXan3OMi8BnVzrkkkPUj8XBwuqTAQV7Vmg3E7E5gTs5/s+AQdBZ
v2Z1skupMS+kD0welXT5/YLjZNgGn5wQrqXA/AvHEE6+ItK8h32tMP5ZuJeBr+9huVBqvzlDXiX0
dVF2ioiUuwPerxSpr2pbpB7K0dURq6y7weAsYXEd1wzfz/29MAW7Jf/eluJpHhAL3z+hPkkprYFi
qJoLuosHIAZzOiscaEMKPN4SD/kjXoJZGPZ53bWKetzFcieKqWfpTWFAf3TufIjcP0BkAxCh55HK
umY6UEkvYXsXa+7tHz7MoZpQyNDvtT1IvsmLeRmaFU1VbasP8Xvn7aZZfOGxRuzzS62wbJi+kXo6
pCfzoauz8ZkkwuOo+CmcWE8QRMaR+VVpe8hMP5f7caefTVKIjAc30GM+ShHo2i24zt8uUEH7dMTj
Yx2BTOpHFiX1UpR975B6tg83E+hvYfoxWM1Lb9GPGDRuBx4CB9XI4a2Bxi5QZQ+OKasoTUbGZLcD
oULW52FKMrQbbHW+or96FOmVWKQS+jb4d2Oc6CQ2oGkjA0O81Kdewoqit1JvAUtDcCZqn+36L818
xei1u5TpbjiaLrVRyI3Iv8XJoFcSDkGqDVGcB+oF/iZPsgWVwdRD/HpraiLfaWxYVDxm1AsjmG3K
hKlviG6UHCjzvV2PqTpvPJDoCO+y0z3qWehTf9VFrmTNUL+oB7m9Pw8M4lEEpuhSy59X2eIlf91i
zt5yhV43pMjxdmp9IXR29ZazZGQJNehXGHVokLfIje2QaYufxk9D80ADObGbcDQ2Joq94TXTfz8c
PIu0AVdZE4OJ01RWQq+bcO+AxgFMxsqGtCz+aCnfrKZagF03YJETayAD26FcKQW7+pEg5IL5geSd
TDOkPuAp9Xo1hxy8Db0c8T79Lo1LTJ2/2GjuJS4PyEuU6mp+RbYzflk1tSgPuTPlUqDXTJT2TSAq
APkM+7Kz1xuC7+eDSRBMrJruJMfa89Ef8uDwSN9RW9A5U8MEuc33oscbOcvXiym4lNfbsYvKti5Q
yS7YKMpLHUrbJgNvvmiv9i2+0CMG+eyVD6SWo6cpRKkQsEdcAuBHvnjKZXjnxuBpz8jMZ1mytOLk
FDp5Z6N2ycrefaE3pW1I6GO/c4CUVgfa4GkIa78xAUTqmzQ+3DtpE26+GXTIffl9aT5yZRbhXzIA
dABXioaTqVXe1Zj+P1MM1h5dFAu6/wOwrBtyfBwuyNK9B02mk+rKyslLKFXOLVLdyrBYNEeSotBE
gGik04DJ2JNlWQN1xMm5D4RcxRh9hs60MRDwHNdBkXgfF7Vq6HGeSpegH65Gx+BCk81ORZHXvnun
ZPUhvQbfBP2wFmeV8SoYp95ZuW/9kLVUjXIW8q/LteLtXBHiozG/0OmnxBPEMqTXSYv6SkTxIESU
gyh10QO/Jsl/MPcQKLlpBT3tkNqMYA74fhLMnc+SBRsn9K8NBkrqfKDHxPWM+75lkC7Wf6ycyt+p
y9wInLl79R9l+P5TXIUMGvtvh0LogKOKI5qvpxbrxBWO0NoeZuackgvd67wb4+ZqliQdSOkV475Q
18/1vQz2u8SAtbtHgS/YbYiBPwP2QsuhaIUvHMZYFJfVt7ltQSJ6bpPIOKSqAivtCzRJMJu9OBOn
sZU27AlTPdpZIBhmhh1QYpQRitxEwxQj/Iej4k3uHY6dCoBtRq+ZNgiF81NyFHwD0rM1XaDa9zlG
anPhSFQ+LpifeA7s3E9c25HWcyzqECfgGRU66wn1kU4DwTX2cX9PB22c4qFD8USMouNont1obhIL
lRRrhl+jb6NU3wP4/w1thMw5AogOfECwJ3kZJq4Yc0jN8cOvz4Lqfjjvc50exkg1nJSrt/aYbzry
OOLTJElGWBe0aD/VgWV/qmlf53F4F7iLQ0hPMH8R4jDlyzAsnUh1F+0CgWCAFVjr/z4jQzcz2ZRW
2ADJgh7L4R76Ym+qim3ONIGGm6Eu+mKxFsK5R9V33Lt1l4SeGeDcbZpFt9lc+dwQeSQdVS7Bupzq
KcMI64ERmL/Z7ubWU7aNIbaozhc0MBuRrvC0Z8gh6YU5TS/69XWMNlrbyVjjmTuqZ2tqxYV5I8Dd
CbRcivIStpJQXOABIahfFA/83k7UipcQEpsfZeqz9gmRwtJG4U7jmzDp8g1TQiQzmPomdTSEaIYz
v10nVekGq6P4vmR6ymU5Fg++UMky7fEs1OldlfOhbH7DezzE5DfVmb9bYVZjvj1Ml0xxQUsEGc9S
UC2Cn85+HX2W5jeGaZpikq1hejNbDOTHH06UxC32mOarmb9o/HptBMsQVkzCJGqoEMW96Fiui8NH
FQqZll0qyuBBs0Zdl628D3DRwnAMVCa05LcZcstbOiPGF7aQBWMAYZLSDJzNDoZga6X8oD0w3gUe
h4cHUqeh0eEM+Rc5Spuoulgn4wJXUlSbYlcBPeGcaDk1Wi5+aQeFG/x2Wb7uRfFLSMPq5t7c3Ku0
ZQvrhzobvhSqerqNXlRRKaUDUKMVcCGUAF17zkS78SKU9oj++ZaRT40mrGmqpVeduVN3+dfyRVvs
v0oEiPIHHJQJrS80w+UyqMjliaky+snMl6ppxvzQjtu5fFkLGhuO+R/cwLt/H5doFPDJcHMpcL1w
CYR5iJv0+4bn5m4sTPFQRYUk1cqjRFnhPODhgkJ/AbwzoztbPRRO7iGO9oUZXm4kCb437wrxvbJq
jmBiiZSTFDPmX9T5ObrFHBsT+cB41S8oaCkH8mkgaUCtbZACRIfjATKtaqGzqQxdKWCx5z2E1O+G
luNmYIiMP/9UzDF43Ajb7TDcytwPTea01883x5PUE4Dh7V3zqcTHJY6fwTqxT5w3rYYIbeYyNVEF
uvh0gQYNpWf7KIAI+i1iMcUXvwXSqtDnxcA0O1xoe8LKTTqzcuydBar5f3Xz9/QjfMKSgvuONKDo
xj7u+zJdmA4jLTWGzirVTClRadpK+PBLvjEMaL5ijfpDLkoWHgtc05rlEJeX94kkD3S3NvsARTbB
Iq05EWtfST1BEwP3ynt4DAthh2XQ7WI/EeBKce8BY0zhtflWTenYCmT7rr3ihisdlIkTMRJVulkG
S+O6aNEyp3y0nKgDsphMn8YuoYErSd6IepryhCDi6m4hUxNvAnfso5MgePbhB7NEd6vUOIL5rLaQ
pDMECnNtL5lGtV34AO4ws5ZcHrgHYTWxWr6szHUUzpXJJUqn7c1mAYjJhK9f/zKKyDH4rSIzPrM8
2olIy86VbjUaRwXX24mznRivflu27IXNi0D7DNONi4UZNjpkHBXx5FTX9av0weqRqvA2flpWfzHT
u+4z/FkeqbY7UmKbFm2T673iGwnwG2yWMTQPuptS18UfLblOWEirpoH7pREGbyWb1Vz8skbKNeRw
y62PJ3n941WR6eUZtPahAW5OkO5dVL8ASX2xmT+tFgSy/zbdcWwPeHTQIWPa+Ph/B4tUIGSG9T6K
YtFJZ1/TrxEpEG8M5/LzeEUldaz7j8SdvIx4DcFkWDgkCrPW9ZqgLDYp2OBNVuMrJJiAd4gIYNyc
bzAOwtzU5r7legX2X7lK+DsxDXYHW/jngE5XzBCljjzYaKKjhSbmwWafp6Undsb1dlsfVUm18NlG
6cYxQ4bvo0vApQAAQN2NER5Rxm5DQlqj7TsE02KcXO7l8DZwSo1mq8cYXxn4EBLRejEULizU2oeB
FUa75AQOcc6uLtZR0wIFy18w7e7HQxNRk+/to0Dkr1ZIrf31EodIjAIgAQt1xWXaxLWp7fe+Reco
3+3R/FOx1R7TfWxhTvF8opNROz2gsJdlLp9bdfyAF9p40bxdi1iFqF7RRs0Q9XPBCKo9O39KVNRO
8O6ZT1jHtTR4Z5YyQk107hiD6BCp/Y1f1QLZ8EY7+UI3srfBiPTtaMIlGn1uet9NzJnA3RXb4kw/
nldthYMccvltSVaBFan23bm1J5ajN9w+Rir6pd1FrZi+pJUxus9LLudIZoHlv8flfZwS7o1lnv3y
UZumzdVVwDQtjt2kGUpq3bC0fB9M1g9Hscat/EoDtawdJm0sKDr9rRBSP5iids01gZm8wMWDRj5t
sydDHpy41zC9jhIh86nVON/n52sGJIvFYPOgcsrF/b8dX1OGn7Y0LmyX4iZ6b7Q7RlEDapIbwNoi
S+g8mR2C5/VWqlQhoEs2JtSw3mPR8hKo/t3WfS43A2HQwsXGP4ngyU+uOlztF0Mbt662rCG8t9Zl
27S6nqEBfjOXzNiar8XW9N9cKxhbHxwUer2kg9MkdPeLFKHA4ZMzpmxXvPe4ltzsak7xXHeMyBjQ
kDWoVUS7AWlnGp9T7LjuHAqD75ix5r/JT6DeZwHDl7tprz/DMxCQLipLeZMpOjDvd4GRuY9Nd8a8
KGi+c8DwV301dLu1PbNeXwrvrEMSgZREKzM8DrAEsp/BPDinrw/6WBOzsUcVFXOv9ZJ9UZZsMZqN
OnKuFqmv4DjS+WgVcd1jYIoc3I6Pc/j66XvBjfoj6WZpQErIsH2sGhfrKXMJdr3FzLeTO9Ygyq+z
NbAMi7prMn0yP78HFB8WYQSgFIawurVZ9SqfKu6Uh8U2XzKA4sdmo6BoanUD1UDncvIZf9JDWRsl
eKmY888QzeVjonBFMqbKRZtS//HdPVA8uVj1UsgqetpSI3d7NlaUoZSCGr58ne/9sRMbFQIJBbFX
nw9HqhBXDvk63blLYBcPJy2rrLsVijtD/Cy3jym6uCMbP5laSCzooLp42l99dpjDivlKeSoNBLKx
YBANubRMCaHIOEK1SOASFFSIETczexXSbZCQN7jF/TZvybj9JAJrlW01qdvvY6O+e7t8Un8uK3fU
rtyxZIOXOhxJZ8j9AkHDS+rue21O0uAB1tnlWskWsIwIqbw8uFFueCP3ZA9hV5lV3ZYTB7ZFxUzI
d756qHwjR6njUCzz4d2s5QwkOrSXKLnAhgR1WhfbbQ+1HI8WserlDAdGz72bTwJZG6qO2C2qk5Mz
8YnI4pFSDKwxpEc94f2A4RHnQGlHZt8GAhSO4YWRSfucaxd4Gw3JIofQj7LtM8R2HhqCzR4yQ6dW
RsLuJhKKyoc6w1hAzQej94RuOIYXirGZBJdpF4DCM2KAnfYT1JcJDezaJCiMCD92wZZoEqlrDIh/
14i2y/LMVAFPUIuM+74IS+inUtTHKW95iTNJ2drzjPt4X2RAkXF5GTRu5DfthO3CD9HPkzcqVIcK
mSYEfSYwmW7oaevUO9kgXAkZ9hyciiJqfjK3z31LIzHw3qHWPsX0mTQ1zw1YdZZsLXuMcbKa5E5j
jpMhXGQ/b9eIwzoPxjFGhbY/0GmCuUN/p0PTyeNcHjOsVhTUCivoZ9ngxMLEvgmW4HSI4taMC/1p
a3RU2oBVyjj6Nz8UMLyOVpbDCcIADIDdij8ZO98q6MO8d7XzpP91on89W/1j44r1fevmz1Wjor+Z
EFZhJ3T6UiefjueKupfsn7Gde8+UVjG5Q0K59Tn7PxKEld4X30It3hWl4ZE4cnhXVFs38xn/yGhN
t/dXDLVuXtq5zLg3lIBUJV3MupU308WK3w2e5uuNNYEk5JhiUUlmh8YljVrSOTF1A4gEJtkBZ9Tw
l8z3yk4slytbdiUNupcB1q9LzYyu+1PbRJge+zkyeS3RmkTf6RDM86lSKGUMoGMqRZ+vD87U7DH+
RktbK19fUO1/qMj86L1RVLXheW7titH4+lOV9DHBNnvjNeho9z1wSYcUB+CCQriLYbmhk6MRDdRd
mLi1EI2FBWulPszrOvWPSXVdMbE1lXVqJAl5yf8I6WqdxQBXD/MQER9bIxNIiyCWgWRe19KrFSqB
NuUwLi22Ks7td0R8SvkA0n+6pLzfr+rJt659iISx9gWQdjJR7iLkZwjrEr4iffax5yDs62GFNR12
r1znSid2KZb9yUlStuLFm6GGxAS5Nmf+3pNrJgsE3nKVqqVZvPyfyFgZA4b/EmT2HDi3SUHWIGUZ
zsJOVjgF3uf0PkWq5787wHUaV+uQXcjpMn31iuLnLukUuEL9/Akt5xLJItBV+JoYAHxQFVBXQiGc
+YV4jTLL4OzgkQmLwD0rorJxbQD5Kq4XblUTK80WY6yHTuh1t58P01YgCuBhPM9VuPgWl9mozbQ8
tNoyFIxnhqObi9WTPXdNvDAzzaZT8KbncB9/tNrPNj/1qNOlA63C9I3BKQRESKMfIZI7v/iBRWq4
1MOl1k0tgzaKNTv3lug7k9LXB5ZZFOFj14ESVhE1rtM2+pkZr+ThHJokmMuba9oWT0PRXrfr8Om1
2D6kM+P0ZwEcvfKI+zv5X7uWZriIc/+PGopKpVducS74XiLU+5P0FIlEgcWnUy0V3u6XkgXIlT96
xQov4TL+23+XyM1Q7uNBOO1DSemF0C5MfpaGhDCbryr7dnBfnvvIPN4a23GHfst6SfxQH1RnuHnO
jTbj3B4++2bYufnHOp2mhtZUSuBpQS2e2RgLUjovkjySivzjQuHMa3RKsthQTKy+MZTrzZ8MfeJ+
EUxxBdMC7c3EIlbvuDA1vEPNQwtLgbqZa8AuVUeyBnj8P04L0cth8TszE3pYzaGU4WQw89DYrp6N
/boDOkKsjm7ZRWS0FUGmseqtONaWCm35a2k6qVHoERIiwS9cd5dVS7ZlZQTx1YjvoN9BdA439CyL
JZIAwPsOJd+IQppQ6sZDc8cXJnXW0z7Lt1Wiu0QmCgZdZQLqeCCBGTjYytt2/gG+Ahmc+4qJspgj
SgB+OEjtHkJMDmi/Vmzz1Ayk7NJ57KjsO7i1r0HfTWsFs1aTdScAK5GtD3VZhJqcaGM3qFnSdXOg
bcUvusPKGRrftWjQhQT36t7U72c1A7ntpAtEXMjMpYD+BjddCJJht/LCZ9538WGkFM+UFGO4XlZJ
dSB9vRCK9UDevRsn1Wnwk04mw45IQy3fO2y6Pytg07kja7gKrrCe0QWdW+qVWGKTY34T5nwNaEiV
yWOqibzJ3axSUZAkVUfSBBh5Ia2EyFkfr6pt9g4lPDvZmHO8LSqMrXb+UoNJeDMJXwAKMVtJLP/6
LU4GVVQEFh2Sd/t+kLS3ayVWGULozN2MyQwzebD7vOWMEjZSvtVcV3w5d53aT3j9YDeoOpd/GXDm
fzk6WO8a/YeHpkTUHnonMjappYjXs4PsNchT3d1OlVmwXd3OQ4EnK2qjvKWEEK4KYMH9jmK1JfJU
EDGG4Huabp+AhuX6KZaWcTZLQzwD2+a3VBRbL/29vJrNpLo5bTymwXAL+uPGeaNvZkb6GNBUPGkV
FGsB0lMGuom/WRHGVgT5yS6CRHQS1Mejyywm2PD0cXiwWeYueJyrMScMROQFZAvpsn66LzJgwKgV
vmq5f0EfNtcJ0sz9Juf3P1u/DgdoyvPQfBNYX8tkGZNEjfEyFPTmFHFUxb9zP0APFACUzkzUGaFt
XKz3Hh8EE1BPcZPetgHkGR6N9wr1SXZ6qn+Uiqh74t18N7WTbYox/QC5+g1pzBA7QgKDUbEzrOPh
K9eXMyhiEiiA+ZlV5mgKJKCsQpLQlY0RkwevV6+D2AZPe36d1WVV0Poq0KRXLnmgQ6wkDSgv9mo/
mRAuRbKHbFPFd1TlACiv87skugrTivUJFkYVKCuD6gE9ujJpYQRPu2lO2AjwW8+3dJ6JPWwXzIWA
jrxdpfZN3Kg/zddV2/VQZBfoyuN9yj97DdZ1jQFTNpcARVyXgRauXA3igf8AMwMRPkWPq8xT7Uxk
UWr17j/TIcnRL8bXg27xU1nly7wCu/xin8d4Xmm9gVMVEUCKA3IQHyArI6GuBTxPiy4x/AsTAKIW
m90BaeydBqrpNUJ4B5pq7k2o95SAtn+vmEz4zCf0QFmTKIw7nj5MAvby9r5cI2dC+Rrc1JuKKNiX
8HUeccEt6PiDWnvSD+nkXUpDxNHOUJzeyl7vxwjdrj9q8gX1i9OJqaQYX0Ni0eTjjDdDTsSru9fR
LA1C4gw01nVkvijXX0ohoxQNk8SRvVbWM1nzkA4/Lq8J0s/qaNPgdajt3yOUMwniSl+6tWfULu+m
Fdic8wh+Jrmild/0i9N0BqttNE2UM/A18wOA2GhtkafsbpExkIQOATETnMkaG4tvw1bavGNJwpA7
IW+9b8whRV0o2rHMqT77IFRoXJBI8b2tB1KlIba5LFGO/JKgvBqOxIoGh4GKWnpSyIAPTuWJ6L0M
3+jYUwQkVdHiBHWv7Ge8c1OF51EkvM75O5O5NP6YYq4hVECjOL3EOJkd/bPIJhIn4SmyEXlmjNFa
d7lixg/Dz3QltSPiMHmILQoLO/CKHFlPDl41IwtKcMc9H/T0kkPuWrW5I+D18MLa8b1nSSiPRn2p
xn5FOhmm6AH+/UrPi8CShZXcZ9ZJ9cLElJzjzxNI2g2De9zLQ2bYDZ5xOV2/lTkZ85eal5zF5+Vf
7gRuiI5DIdEUQC6ROa0cVM/H5rlfZgMS7szYPGF6G45QbVaC5HTUnGwD5NLYN3/ARmAZzhzS4vK0
ZYjHHHjFQvNnneK9I7qvvRA8wROXTmKLWzU1b86fVDvMc89rvgZcRvWd05RhUi//DKcqNAl/Ke3N
TlIDY651pfBxzddQkcs+NEUo26MV8J9/+MURhy6B/OU2vj34BF00OfeGVGJ6AG4ijeocJc49/5qw
Si0DdG36B0/TBWbVlbLO/fkYr5YIvVBCk6xezSKlsI+yLXDxXFTPl65XHWguWb7WzQgyRpqvtGJa
Ka7P6Dlx3Eqqa11jnJ+0CZh+HRa68750rMqkT7WD4UkelMHtjDnRHDJI8pT0u9UUCiFUZR30GyaQ
mhpvNusS0RAlLn4e2Z8kfLOZby588TuoYhsi6UqecjW0xThk6wZ11NIa6QB0Qe5Ox37XhFNzegQi
q53/z/1dqSaWnFSjsVYh5RCDaeFK00kgpLPdce3prJiTYG1rzCxVgkOg8nblZnEneB2F4fwGyybY
S3vGUFmHmjDONl5Qdh1I9ov9BpNSrzzpmLyZ9tIeww4ZAlwFLkWfXk2dvbDf0DFcncJ0YhZ1XRSA
k4nDfCmSvKGGP2k0Tc+lvlRHDIwFe7n0cbel+OME+cVmhkvSuZoqvmi1U4R2kBFsILwzwNjNOF+Y
r1ml+aU5Oiul0V8pd/ibggO2hTKreBz5BBxUezO0b2ITosAh6dEmVbY9vaAlma6fCvmONJdOJ20C
d7CmKC/djqRC9D5oBr2oilHdXErS1ljVv84MLsdq8zOWEdjgIAaRmW7a29PNeIBPOYADe80/7BfK
XEkalm88jNLD5DY8AJWSRBuZZFqQCf5jcuj7lcMzUq9tpGawzqSMDfxWIes/tRQOJooaSFiJviD5
eVlm6qC7aWhy7byfbeauofeLtvMVOdKjq1I64tj7cCYp0XpxlB3DKzzXnIkK794kYSR3RB0+bsiN
Q4L4TVq3WQXeEWoeZN5i+aPzifukJ2L95nEu8X25gGsqcsfstviggxDioNtQ8grCjE3cP7DEq6J/
B9nLKyl1PlC4yQTAxB0n8VchBmSPJAiayQavCNNMr7WTSUUO5ftEMep8zlzoxU4edI0+T7+Jr1uJ
MmTwwxbtO/ejwbH5mc1NCRe71ellu3YhaATqqsPaXPCFEfDFtn9zpHe2acC5m0D6CQ33pSnZN1Yq
VxF3JSUmWjYVRFQgMg2rYP3/ijLmqBvjhCWccC559X23HiGsKYU+PvnNG+VJHgpF/YTAGOl3iWhW
W9MC1g7i4q7MKeeQy47XdAPzp0voh5Wx169T33etuqOCiLx/nCvsBACDN6zm2oEWbbiTDdP1Kv9G
x++KSPnxlCWGYsGzy1g4raR/AuTxqA+QDkFgL+j2KUSbbcUTcinOcQlXse59PED2jYQtX0CvRvfd
6TVu2BBXnGt/SBv1xd3ytkTTzOcBpgp7SYMh++YY1NSGJrb/AJGB8ZzEmODzveIWgcrYKdkBJXlr
ui8eQhL3I3YRgvrAvs2jgbkz4gGbc50E4bpdm+aZfxvY49a2ZZLKjho0+LnTx9cxXMSEFgnb62jM
j7vTrP8ebmW8MQZSULwV3ty7VQ3acUCSzI9YLyAGpbws0e96ydQmX7Qd9/mTxSUMFDHSTplUP7WP
o4ShE5K6SMOcCxQ1n7e6rIhiu3ttZzGyc1pdR5VYMUmBXWxNeDaHclONz2ZfRUmLSlIOC7CM32sD
Zou6s274hg+wQUZJzQeUDrYxqWsEf6r/tA3Is1Xnf25RvexS2+IA+V0jqr21uyKaByhDaoyp/HsL
WQzhpJLTpv+kIZEnQm2cNnTB6HkZzT0nJUNRWWtg3X9Pu+569Hq9hvMvf7d+JXeJtM14azdF28pM
HBksTfQKGq2Ic/oxi6/5FI+Po3kRNQ2SRHkWb9ueybaCIpBOcFovTjsvvNIiDVilBdxBzQUJVDtw
LWOEmTdVB/H6avdGYqXujl+lSH4lmjuRbvF8U26ifMhpeHncUGeNFsozOXWXBKygFJxmYUtVZSSn
N9u3UG5Lfefrv8Tmc9wa5CJhOuVhH85MpCBFuq6DwNrBhwSUJ1I5D7HvsdJycwtD+Fn8gbR6nBvM
9cwz7Msbja4J16A/807OjnwffC68p3LVHalhUpTuy6fLcq94axQSwb0oj3aeJJMOMKvtJhj/7Kr5
2fU0bZPvQNjfkUIuqot/fmYK08cMbH9AuEbj2d2rRpzArxJAPtm4ANF3jtoMIkHxg8L28wxl2OkV
tWutVdKe24OX2gnIGXkP8cwMZ5LxxQGOCI+rLhS6FQA8hdCO7BVzecg+MS8YtMfARxytkUIlyqDU
ine5r7vwSI1l1b6FfISnsZXB3Muw+DQjuQgRvUnBsA3XeLmlr7qR7DQTdJhRkilrQv76YyL8EUTu
t74hbMbdx25K1NAYmIOMRuH3UX5SQRU1iswG1z86E4Gq7telC52DagrDZfgtokKVAEJLQ8PXQ+k1
os7WNkp3jMNOcDpAL/KaLhSDqi/17VCS6YU2t7VglWuAmkIMQk1cI5PhEeTQQ/AVgn5LBlto5BHL
mOf+EB3IYRvTjSZrNo262h2bkb65jkYYe1sxYpshGRpjQqTxiyX4xwAKM/GXiLzI0GFg1uGIetO8
ki71urY0aFA2KmvbD2O0VBoOTrb/W3N5e3iTA0YS66rTKxGciTVGqC5mgY1DzTsqX4EDevlpiDt6
N8Et1ZZZVrmtELoofTZ3EIL+/foNTojBXxsCY4nRPjbpBsEe/M8HxJLz08afF8NLLWVvDm5cCFS2
QzknDpkgeG5kKHdtm/63CLEHYr2PWguI3R6btyi5PvAXHf0v40nLbD4Vr7Ukiv8MxC1Sn/GdYICs
8Xd7H7BPLec99LfQ/emYE0Y2mt14wQ5TXSDtF55CRHV0Jaf/dKT4tKDiSNDG0rI4WJuKxQgTQU/n
jVEiNntaDxUm4egpQgeHCsWSZW/47LuHkTQlnSJ/9yVT6pjIPN5v+PdvLRhKUleS8iLb2H9Arjt6
YT+vX/ysDLIUeeM0eorsXyJvpai5+K+0MKEIaQ6m2xWJynQxGUNBn5w0D+P9jqa7Zc80QEi99J5i
8C785Uh9NvRZGnLOri38uPAMPab1Pq7FDEBseaQH74KGtAP6Ksp3l+j6O9vX1sob0rIhB4pIp98D
sHEx5PBljg4K9FDOIJeTwmPXB5ur5BPMdp9Xf7tXNfXzzSUWLrpXuWNvuF4QC4r/76AlgqEspvsx
xec7FgqxujnoIJsr9m3jmX4/WwAtXpAIAsN4iCInEw0p3sm/I/xs3/+EZn/yRzRPUBnkNKj4zgxM
zp4R3GOw5ZxAJRip0wmn7A9bJKeuB/RBeaL0Mm4A0xF6d1VUHrdcNXb2ICsHZhMYG1W8x+QhcQ/V
WH1nWAXQRfh2DRg/FRrg71vbV3kXohrY3REZIoBqYRWTSx6qFaY9URAla5+A6/CIX/798fhWIgoZ
S5AcFN00ZPLQgxPAyP0hg/1vgrZrvyOgetIsQ6G61DN/23SXd/6WMMwKWwvlmAxMUbyxi//u00nZ
QPeKAcnJfVrg13pKjuaYOFO8xscqcCK1i8FzFcXx3jKFrYwZeoVqdU/uIzJGUOTnswcPsyZbkcm2
Avx9BZXlGDCcba7PoqWsNECZatflhKhBR0GnmChXt58U7aX21bk1pmUckkPVTRXmD5VD4E6596kF
+eXFUPfFbldqXNstaoe85H1smrKf89AXjG8OTL1agJx5NZLJTXgAlejjmnouR7FOnI+VhYfrriOa
I3PCxkyXbS6oTpUzk0Dw6LfPluH2LNctFbrEvX6c/GCbUM8enUUuDibbSrKrqRidD7bW7Js7cMky
fw/Lte25l8reT973uR4OZmu8E3Ww6CIpokBiDA/Rpj8gjvboKo1mzPFyj3AbJupC1Li6lIZUfMZt
Fhl6UJZiEUzy7+SCC0GpfDessTVKVTmIFTDUUDS0B3nVc6Zbcl1td6EGXzzEqVBZTtrzpW9nNmUP
BDfn9TsSz8USyk5Bq8x+XWL8NTl5zWrhgrhC9kQtaOfk98xWXYRpmx04aHNVm67aPnSeAMFJ1asL
qAYIek1bsllwwX/tNy+8dQMVif8Ic8LfC6KmkyWJvNALc/CPCKAssXTqbQ8OqbraLsvjIKLAdHw5
OItx9TqDhhzqEa3WrfnfG1isA1GDTy8DEgPyFYVSSMPVeX1CxjaNSe5GqjeKjEHu2pzrGuYlJvC8
t1JSVvdMZ3b74kFXJ1vTvQ8D9GZKA6qfVJGgXE1SBY39b27sOp3FKWSco9/qnTEsyQZeBs8wUFjj
owHV0M5OiyrcuFyTjtDrFLmhF50kGqzDFX27IQkJ70M2aARyEkVZmfCh9/GFsI3iN2+TyhX3s0py
f0TgpEdLFRRcm9M69XW9CfjNPGW1C5Aw/NcgCLFgVwT59T2G1oxntBni6aNBcS7Ik58CXxDLw5nJ
DsCEwij1hNLkk2ombi4jcEDpxjQsy0qFlMX1uGHAkRdmEbvlZ7FFZbZ/+q4GXEjh12ci2VRLCv/A
COwxO4cFUbj/+gy0ESl3Vt1rHHTlEHNi5JQI6aIjD+NLtPf/Bq1N4OCu/b0EiA8SMh8xtClv7isY
CiIvVxErFI4YYd8EXScz2b5pUrGR+BM9MOn5gxVt3aOVG65pEuP1tzNuljRnUF4yOlX5qbr7ihIi
Pwujrhcge/WgqMXJdLlFBSeC5pIK+43xNcAKXIYvkh56C1gtPHUVz157l6byWMVuzc9BsVecomVs
NosJSci0WrOTJnt27czgmKO+97E7QF0I+W0d74yORn9oHVlY9EZxRvgM6j8ao+yhVRq81lpQCgFo
6CDx5Vve/AdBgi1k60BnMJVUNfltiQzrGu7SGfBqJFgivG4pdrXSKrMbEm3OzqfysGrqy92fIDob
E6dXe2S1kF++VqZszM0CupEz0CtVy99db8EyWCg6WRqDsIec2QvGItjmfxLz6aI4AJgxIj+RlW9g
mRb2oAlXiF5U/MXDqh3CblClBQig/4+JFl4yrXLx6m/wOtRZnsAIvNnlsXxD1b+4uolp5SiAorMB
lzca1iYFck/sr2k3rrt/Vzf8waFb17b7SSt/ugeCEVT4IUIKMjHX9tuc5EYS2d9vFv/sXXZByUym
8BnINnHf4hr8gc140oLQTDvFbjCLkWoPPVp68xdBsF+3978DS/nkHzZhQxSy04V3AlLShu28wE2d
kq37Sz+NcfWo3xUN/3Wz8SZHdxQrCKLkAnSBCrKaah2BpGhlrZe/CIiH07zsYzdUA4qNyQ1V4fqD
kXXER2US5SzeECSmmTzhabGrmtM4EuQ4nxCtD6qd9EfQOhS3o6Ie9bmKdi7+HY+ryJVaRxqnaDEy
Klu1iJpOmAPS86iX6rB+m1QDmOevMuk2/n4Bh4Keyku7/isJbhq3cLVtKq268uu020fp4bZHblqT
VxEuu6D9cZWiajtZN4Ax9RkmfQ1CByMiIsLOYmQA3Cqzz9e/5p52axfUdRxXD338V6B9i5fBrByh
8iDRpI7DNyQwT0W7HXO4YpmCwjjcQj+Fjze3mYi4yr1EQGylgQ/bp1otIo6k/ay/q8Z/oR4ZHgim
4QX8CS4Mg816/hSG1NFQQPlaVoEefcASoCZrYGdEin4uA/597v7uqebPSOWWN0sOvQ+QMzLA7GJU
OGNMCc378LPADFLV+yyaTyfL2HKCGnW7Ymkk5Spn5lzxF5gvj07D4ozBiX7r2Y7fT5vPmoQO9dFL
WxIZUVK/WDGJJbQmLQoG6XPT6pV0f4TRZ/ZbjvICVi4snzurrwlBTwI2vQMfOJIHhmiDbcRJedrt
Jvz1AsHmRIEdiV/LvCz9eP1VZjG3QkRHU30OhdSZQOj8NPzMebmH9NcBThA/yy7tHdj7baQ58I3D
OKKf7ZHa1Nn1aGjBI+1e2mg2y/qXNSSQ5ZxGAMJNDrGf3ptji+IgG2oLg6O95qh4SuafFh+5rFVm
EGqEjYRIlhkUbjXPlQMDd1Wa38dMT8M8vWnoIEyGf/Z8Az4daVkLZTthA1+FQp7sMF+2efSmGRrk
KjZUCjWj6O5thLq9W6ENcQHzGkYwRwqMUeEaWcowwywjUPMR2unAevEqaz/H34gLEyx9oxncXmne
yjgS5V1JE048/ztnSbPeg3eEpcWFTlkELIV4uXme5Fxs23lKANSpo+Z7E3YjY9hqfLp3kE2ci4um
3ALide+Lq9yy95HWuVw0bkj785h4G+1PMMT7JowXzgx3lccymLMzNvojULaB/Z7nR2EbPONPau+v
gHq/oqftvXjL0WyA5ueeZs8aIxFJB8CZc/JhTqdLZO7MjkBt76l6qBLcCBT7t8FyZWC4vT0YUXKA
uXsJH1I3RdUsSiIGpRWUiyCbr/6IAkhqMD5UXEOXIau4qdffurVin6oBeNnK8ZmU+7uuXcnLkwIs
OljBPrep4Jb1lKhYp6ekB9o0BTwsFVIFkoemfMqTQ6RqAcRvwtX6RHrjqMfSMUqPP7WfQp8xTK2/
UGnDS7yNvMc0DpGA5BR+kvnPU9fq0Mfu7H2EvkJ7nNK9uHgacTI2tmyT5Rj0PNuMoz8uB5XmBBcm
8Hj5f4nX1SmYvszkuEgc1VBu0l3wYVD8udP+njQaBpBPwIMf+IXH/GqaBXZUrdXrH7GaNvxndd/8
XCvU/0ZuPSma2KyPRdz7WbWNLn7V1iPeBqXMUJ9vzNe5TltzkDrl8oYdFl5n/R6HNuhCXhynONj/
5S4PNfCPrmT79rZvSlrN+HZHAE9vLeiLuNErQ2eERdaiRaVgnRUiMVCUnZ/p/+efTnpQslvI2Ouc
t+iZXPfeQ7D1v1YPwM/er2uDSnGLYImLzL38OYrODcVVAWnJMGPk0hEPSdHiDAjfAgH5cgPosW40
O+OIZxm/l4joKPiuwiNmB7uy1FX1au15Qe5PQhZxCQ+XfaAF8fzVbBC/gj4a/hhVMV6xAr1A9OuR
UEnp3OtnVBDRFR2EXfbMFSbN1w3tVKNdyLPXay/IL0uh+BO+//2n7G7wM+XSIR7Fs8R6cm06aAGE
o4YG0K0W0sXlu1kzKWtIpkRtU8sJxzBeLq76ZEhrg6kv+1gFxUZWEBzBJ+pWD5IUqfX14CkBeKkk
vFXX6RJbo00k9YQCi7ZzTw1Y7snus7y5c+8oWyt9KROety/LsOG2CVHaa5fmXNA4+TD+5qbKexD9
ILEHP4CV6WfU9i3mEHHBUZv/rM0n680xLspkMgCZOSbCa9swnArhHZWccc1/QnP/gK9lq2K+0n1F
xWK8yafu82e5PGEoMmVPO/tjVflUOkORFCQQ0/vytdSOQEJzqdz8qelplSq3H13YwfONz7J3fXQ+
gIXYAVf7diAz+FJQYfv0/KG83cXBp22lwiFXcZnZlJb0enEdztRAIikXa3fRFqqgCp07AxTuCNIv
s96fnI37LdA/WY5yLvjyWrIX3+G60mlV9zPlg1sKHJ2kRImsaaWxuXpJs2TWhXf262YXY4Ir/d4c
nO9m73q3M1NQ7+CQGqLg85KOBNzazIVCyQEcUcKc3B54LEnGV+b94gQwSo574QfkjitndQB/Ix00
f9vx8zYf66q9CCuRQZ1oj8Ia6hS0LvPkicy5ztoUb4kYOtsrG5OVXHArLFYXCJswSVFfU4wojwuT
MgiXugraQsa4DM2Y/utsgRHJGZgViPOpaLClFoAJMFJGhZsBKVlZr5LUDZuwFyA+fANqMRMFDDwG
106xEZ28aGnOriXnTqym/NndaMvBmn7j61JNXHfFENqDNLBs+9lGa13zJ4HLLZ5HB594I6ad2rER
cPr100n3gPVwxgYYFBcqpKwh8EHeZfkJmoo00ekGydSmF1vBDUDll7G+lE/6KmerCw6XDNuxMykq
sU8CG6qTHTyEDBlyoVvfGyG+1l4AN1fBOBtpdo8ZJrdhj1AdpCKCBRyHztdXhlNocQgbgvBfl/wG
SUGvPEhQK/9BjCQTUfNBkoLZL/5WDzdCKthuT1mCOC939r0jAHirr1IDX7MWrf2EcoAVRlsxmA64
/4mKSGfaYjn5fwwyXIx+QmOf/F4hsLCG65Zg8cnYPby3OaC4/I4Sb/6mt2BOzVsyGFHdyErtXKRG
Un3gdpDGJfSYtJEljDg5ldkKfLtmd6l+LatAnn1KdyuFYkpPD6SVni1oa/EV6DCLY4mZdxClZlYx
1ImWYdHNLA3xiK9rq36szGD9R8815SWcmeKvS1Wj2CKHQLfXiqZHs/KQh0x88gs3U5CmrxRCQ5gl
T1Et2/XpPDFfGJQvxej+vtDPuylRyJ3FgYgu80hd3nZ0DumBQIwH9eXxMwgzBNXwc/3wHHLdLgOE
lc0JtsKHhQA4ig9JrWMVYhb4itO0E3z2oXolfBOOoa5FGK88ogzVBpP4TogIKhiwSF1VNfeWFZmV
bOCYLLHzL+Ty+EwXm8hoNVPXDZLBoo3iqdLNL1AHFCu1U3KW82fO3pkBvJcHdA/Rbigx1QXbzcF/
W+ZTxVoh6uRvXBpsmvAbhmEgUsrDoxstK/9HsvfrpNzgFA2UKRo0BgDl1632g4vYTgPufQB3kuom
aPW96t3GuqSxPMc3oxgf6xUJn6wkIEIjOxkxkH+wqAUaFPO2fjq342AzRPHUyUp6CIxO8T+UpWWu
k+hKaCnoM/qhsYk/l84JP3AJUxPUhhC5RnN1F7v7PMR1il5VigU/rVU7Ux5M4kdGQzLcE9UY/dtH
M0+AsGSvwxmijR0RKrPq+kpfT5sCHRQWd+ntQD3D6HbYzXKmVaKnBC/qEPhNKiqqbPw0a9/suIg8
Is0HISQs8naMDESYEZ7D4hcZ+eIlRtN3Iy+GE6Crbu5hz8lhmoU45sZIsPi5TybK33J7Cjtprc2F
2rA/FwTNRHp900kOQ0U4Jv5qFh8Rs1WLAAL1EfDulIfl3QXATePJ95v2fIUNlKxeDTQwwYpn7l0D
oPb5auZlX2Z9Z07a3KbSjDsoUq0oCCtmZkHB+3b3qtKz5YNpmHpfe0jUOgEKmux6uDlErc+yTYnm
QVwc1ijB6ZozOsg/OUlEIfTahczt1zxyBAmfTKzwZo3IjBKe79S6aF7yPqaYSQuORpKp58XCFOlZ
CbTSTcqY3M2JLSm2JV+qGCuPvZj2ZOxy8I4xzpYI4l3JEv1oThXY/zW9Yn3OaK5HAoT90FZXkK9V
Q5NIYEtI7li/F/k93P6n+IclIGGXEM8yTv3hhpwagEoCkRJ/ysRnbAFlXTisCpwtwYs43/50CFNr
qW59DX5cwugFVAorRuEOjmmZ3O9OnJnM7ExEsC+1hR8BBZfXVKmriBwflR0/6t+pjV4LGTKzyksP
73yGx5CP/fKISO70Ev7mqf2mFmU6ngX8REKGWfClEFJ8AqSe7J8ZBJ5o1z7qXsFD3d4W8fIPsskq
GWjEbr3Ms53/s2tKA1T5QU8l0Qo8O3+vFDQkezIzMsOLyY3trobHFSxGeL7UszdtuPdeqKhmqBMw
aHB2o4fqEReJx4xEk/7acrliOQsJ4sIxy2qWObH5v+n9yr8SnZbH4zzcfH+7ToCr3mNke0pjQL5z
88nnZ/K3mkW8f/HPs4fTozMUBxXUT72rW2vLZIAUOLA1w5ehAwdqHtHnHDgJEXSteXwIrxo/rAqC
Knt9Q366yY9SEJ0LNuK7/+DcusailLtXtxPtdDxeiUEy4QCiCeSt7WgGIX2HBJSCjFALHDHcTMei
GyRysI9Zti3CTD7Mg5PTRH9cpSwyrJMSH+TukBuPzv28efwHfc/mar5YelMLihD9SN3wVHJaU/n1
2Jj9epx1kC42ZxwZgkk2Wp7gdY0/Qo3TEmeGSuwTuuLV3JvtxdZhX4dicfK4dBn6te5mH3trxzdD
xWI255QRQa1guS7Nt0ppowvENUzUMXFDRNnlWGnq3xa8JAR1hoLUGrNo8sad5kTYnrQyIRoD/NAr
fmsWQzQbetOiQ+Vyiaqa5eSRHDrOXTdFtT0XD9KKl4vLPYqkN40PQoyGVlN6l8yM3d3RayHe5ycI
R3ftSlDhStP8f8Z7y1WqYlj9pNeThRHuzTfUrjZnZGTSt3MG0VVR/s8d2PxXQbjoEDAM/ZeitqW8
qrKNqm2P/rlWgAKZqx9rwY8gcq7w8XknPnkq96mOh4YI9CFR8vhDzArRUSal7RtQy+mHmXskF2w6
82r1RvY82CS9JgwjqqkduWD8aiaYmaWcWjh0geQVnw51IKXqMnklYI9oHRkVDEVYGKDi3ZCt/oKJ
/qOhon6c0K9VFztq5mesGuzU4lcHzy0rcdE2BA8kktYxhCf2TfY3xEnXFbVkNqPK7E71/To1UVQ4
8NPKAprKaqOhenzjeYuhx1omELpdh2cnYIzt1RN23wjcJ3qCbsfdaePkPK+Ewvo7Z7WtHt6Kr2GO
pKUbtnyrb2i2zh1dlWOg/y+Rs3gmNLyidWndYuRvyPkXllGSbHGZGTT+nOw7zPy4Vw7G4b6Im0+A
3oP1bWBqmkxlosQ/ZSupzObq0ltU++P9+dN+HwwGW5y6q1oB5u9bwl4Ug5fLWQEpzKd07PO6msuE
UTOFbrzRIQxB2sY1x1lbRz2cNZcYigQC+3NYn3gxbcUaJ1bGRXj10jvQi9mFTt0EW25KEj82qfcJ
nkn16mMk0/u9jIGdQf/ZdO24HUNtFRRDGrH7bFaWPKk6GjhIuNOcWZvvuJ8Ivle1RQj5UPl3L9Tj
NNqmcikFeEoSTV1FGphBKUAj0m+Qr7ag/SBoWpBuvMPPNmM3mQXb84wz/RLruhkdqk01IOkfR0wh
7Je8KsdLZjePd+yjQ4nm2TCfX7JpP6M7ByiIFOQSWSEbQ86W0KF22imwI7t1ti6wSqBNy9Le1v1Y
wQ/S5lxD50IB7n104upglCK+8OyLY7ry1wUCGukVKaeizuZW3Xf7MzhC2Na26L2IUFbqNjX3H/Db
yjDU6o6hzqykZx0EzfldHJHSBp+BBOXH+1O7Yj9XzkxUH0YsumUdwPd34mI8+Uy+h0D1Db6KysD3
Ky5ewjyIj2kukIVo8BuZGUEC5eOPWGZ69zyTuAjwDRHDAs6cfIv7d8Lsr5Uw5AdfTSHea37Kx3wD
7ogBp0p4DfChDh1mHfKvkdMTFc0FrPWJBkU/QzY5HSvh7M0tp76CczA+hsFm95CQpaMRMEOSdn2E
F9tO0ThR3sN7DDuceZqEJYrQ9Y25qJ9VxS1dv5dzs0rvMGagcJ0oSG1cNBdWneDkk9p0eQroqXm2
iFR7XFLu956zlsM7XX7N8MY1DNb+TGMEgMfCIy4CtG+69W8vhJbfi4m5fxQiofvpzPahFpXRkO8+
C0cS4h+o02ImnfGL6+VqlQX+JhOQLNikIbmYqvUwKT2+3ZOqQGNwVbpTxsW+KB0tEIHhRWFsVLqI
cXdVobcGuZ4JP5sxJ74A/+CEo8heEvrtf69IE/oJCvnKQMOslK0+km8X8i+E3HcjBb3WspE9Ur8x
ZfErd3/0ZG8SRbKpOLLcsEfmzJFZJ6PAHY1jtxv4DnQLjKQ7F8hFrvMTbIq9Y2nCiv+IwdqqOL/p
6sPVRbkG169Ex15ibB20kFHbI7f5FGEB0BKTtTNeyz26Wgp2wYiIiL/+3bnLKei7zpnyKVeFiI17
XS3JCw9QCFuMWuJWhWLREqLmNlQtWW3wvOWHcHxbeOixIXTdY9xMD41/kUTG1YitRIZ7UBpNLjYc
et+zplG0Xbs849zih+ntrLiLvVlsSNRNtSEIe4pfcBkwyg2RTGmuOfET6k6UbMhKQM7mlW7b4MzL
enfwH3354OrWs/4ZUZisf0vCgE4xUwGeWukmm3rEWmdp+VcXQElQ17BCdbwUmrBU8YMekRvMOC3/
pjSpa/9jd3JabLM020FqyL6ID8YnTmmh4tJxx7Vn1v4J/rNoHCO0KAZUfSAH7o+McNT/DX26tw3c
I+9nSZi9CMAJsDo0EwCB51YmdoddIB5AZ7WlImrf5k6XYvU0BNK6W2PGVTNj8nipAsOnN7jIixJM
lGgXvPvWMjrA+P8GkJo5YVu8mmaks1N2+hxtEdpNjOn9cV3YHd19+z8B2CUYuJNIrbbvRUZEeC2E
rxLHfCI3unq/MTe1zZfRPOEJ3S6ibYhXnWhDpeB4UD8BaYg9NSIV8GLnIDdv5CRLm5wKUj23BZqi
RfbyG3050wZZ5qpRVWuPNAmCvWP6+FP8o8HRlY7S4aQ/1UvBqbNcs84WaJzFMMiNBvEaPdznUtDK
GITgTNqxawXCAeFDSZqLPIcQsFhpefbkwSTkb4NuwQBGbFcIv4AShXtF+uqyEH7RbFjpk30yNoL3
BCJtcubRiq0osHgbSViqUp/kZPW/TPSUv3bODyEmx61ClgwRczGSR8FyWQqvPX7Su4vxqwaZDnF8
eKk35iz1+W7PI7e761ZcxSyGf0WmFNcAJx959ejXYS1VNyVvy+AeefBbrgAJiiM4g11DOrmfzslp
t7ex8s2Sz7xdeut+GRpxGzf4odxDlernZi7rcvWDp8VQnWrAogt+HOeY1FXygE/yV5c2Zm1JmrwD
0PFZRKJ6vXWldhWanBzb3yrs5mez8I2V2KQOnM+MRGGz4RyBhHfkoKCxbz9OyxQ+5CsTULYu2aij
uZ8vvfeoydp8wGFj9u189Yj/k3iH3woD47zY+n2YuAeB0vtHxgNz3fFm9gKpHogr7PrdDJp2RIFc
2iRsWlmkZu9b2L6cMC1YdB3CVsCSoUON5XUqrYXkLiqpHCHz2C3zvzKvH+ZzU02IYq/nQbe1dZ5S
a7tfVucn5x2ZGqt+vTld/zCi5AFmnpejPav+r8TGfxr0u9tCd0JsEfQZpre1z5OVWm5hmpQN8eO5
vsR+uEw7Ndz5XBedyrZjOYBJZv4czbPy6a5sKE7b4hysZ7cQa2pLipol+coO75t76uQLrgR19gkF
btIMAi0+VeSn8baGOjf8Rr7mHfYAumM9jVHaIXQNo7ktb2/2X+qFblXe14/c0Gmm81H5/QUiH0/K
9WQbG5jsv/pTfFfFdj1bXOgIk8nUVUwHA+UaSxWn5zxpTtWAKziLt8gDAFzIIAuPbYksCPVjvu61
fooD8hPDRQMfrMX2VT83S/oGAqMuiXq9pF6mZWJCWi7KGxEAACbO1MZvKGgzVkOhxSYRpJtPFYDl
vM8rw4+MSPprfoDKDzjflmUQhpvzoUQnSsWzaQZlAOaulcNbruKzVHhhtDMqY5O1gzJ/MfWwHX2v
2ymA3vFrnMjcerTxUWq0VDUI9KeYoz40xRLfz+9uEIa17XKpJwBMqZn6nmAWkafL81mU6O+HLld3
gRp4Ieb5ttVf1/kAAHwRd2AMizXFqHi2pip+sR/6vfOcpoOWrYUzCuPTG3kvDK3u648pBoQJ66Qt
H7clXfejzKtPEzo56qmdCLgghZcM8pSnzV81LtA+9HUHRD34iTt8gp2YVYHZa9XQG3MWtbq8sins
jxo1zKhlTgUmKIQvSArc+sJEgftYNnOkex17WM2crOKjSUqlsv0txi4G/1xWBMM6MWfmj6zy+P5G
NZnNcF/2Qj93wfqiUNOW8yoTAS/tQ7RCx2rdriRTEL3qiM3yWSh8c43Ukg5zHkrCutzmFk+AMuN/
HtjPJ51DthD8QQWE3Ekzcihtdo/s17SXH2D9/zuLXELo08TfaxHJpBz776KwD0G1oJV2fAtz7GEC
sVdnGQ6gzujlrQoxPd+QbCpcGBCUBztcfKkdYTB3Y8wH3NFYjUEyc1sUjZjuxIUPJJyFpdWJMcCy
qTPxbzVEaA08Qeqh/V8+jkgFqfizit0Ld6sobq9zTFVTRBJqMYIk6V316CTgpei9bE5BSATU+5Ww
U41oJ10dDUQvCgypi5UO804vDL7dnGUoeRPA907MSmyCR1dmr5VVQuioGBUqMZcr3I3CBAonXDEk
C/sJAY5vWUKb0Q0vYPuFjAWft5dOaQpOIxYaDEBS/czo1xQ0myGnrKsBuhVX/hncg+qxxWmT6zd3
xIl3vg5OzNBh/djl9hBcfj/jGnujJoI5amQ+iBTiMa/PPuvpZDYYY6DI5hMFa/N6rOBC0uVSBylW
H+9rzbjIIjOs8snUTCAiXhy85e6iuUMjOQVS8rD3omRMgRKo62BgVgxX0jZAphUPeGoUgZkCchIx
feUmDikBgadWyySgtrBaxHsJ9HAeeh6rJCaWs0VdOWOAPh7VVYo7rb6inpbX9DXzDabxS1/CnNDS
t126WP7dRqfXzI3ACQOA97JUnWfTV7AxtaP7iaoVKZRpg8CU8yTe2QKtV9KYW2EpSaEppjOGbZdP
qPEU7Z3TzDyElC8IaXiE0SomiknCetHafdvHtvo2OLO/h7E8RSxGlkkwx3TkrVsLQ9eQVmcjbHFc
0eIuk1eNcE6HNdLVjwf0twMYXWH8Nii9N4OFpO6IhNwYx8ptq1hI34AO0aPUqtE8FZE9953bZwWY
nsEaqTcZuHq8nJs4uJJnsoggxrLE2bU5b9oJPQaLqKfM6VJAt1t9eMLEQmDhp9DV2KhcVHHHCHlS
pgc05qozJGrG0vCEMU3qFslxOA05gk5qwwfRviZf5f5tsJdCmqa7anytRCBqg9W/7NdiRD6DPifo
sEOv0BsEFlT47u75mRdfGSvOMZTH1HHmWGTbuStPJp0aiGdDT4P9SDRPajskF31M/zTTDoowdrIj
UGi5sO3ZitOw5rV7VGa91JUTyezoaV9sU2mcJDrDtwlTontcFYqO6t5fz46DMI/5yOzW7gD+je9r
IPs1H0W00xLmLnb0dmO3bil6LQGLHNraQ0uMw+WOvGUmJglMT9btZ3mFy2PaM0atvr0xYr8nOB8J
aMC2TKVM/+QsYDOGAQ6WHSw2Somvdh15UwLrjoIONSnisVqAR6jQa7NMJYODWnACzqQg4BOqXJjp
N+ObncUBYxrKt5hRJg7VImjAQFpdvqn42zk+rADX20zVdWmM9Sz3qdak1g3PCpK6TdrQhA5FC0hz
+FqEGwmNPIjokboN/0vU5vGB7I9R7tznBuc/3Kv/ZarQPa2dwnVnNoToFMufBiDtzrfAFixqglXY
O4lxTG4ZrUDY92u46DjRHW6lho1uMgJp0qjvIzqVdTpSYWX4TdsnxmYy1Y8FPkiHS19rtoDHq+4z
7dMsFHVUIk02ax3JJgay46AChFRIP0NNNfbNPI1WcdIoIy0T/P2O/qHc8Zz4nG/r/VMxhf6EGP8Q
y4P0o2lN2mIezEif7k5ApA1CbeErSfUGnhjkfJ5QNwy2QjRuzZihUOonreC0a9gCM4ehxD5UJSbO
BGIBuhMGVpywrWw34yMYh3hZ6aiSgg1NYmtKFCYbRho4kVsSCHoALj1vVQJJuCobj032mfXQXTxf
GyR7wHzQD6ZNWa7PQg3Qvca3uF7NFjJelm0BOMuUbu8D4R8lv7juuETHoIbcXp562O+KPBPWLxE+
RA/wJLGoe4FUvGXl7NdYHXmiiJuIGpsQei9BobNkH+gMS7Md7TOPxYyjj2/Jas+x/5iF2Tvk65oV
CKlegWXsFOiWl0zA/n72qQSfCurQqIa6CRVul6tGEr/Eltwyz+Hv6TRS0u5u3h1FpwxM2qhKwwrh
523WpxS9TCynZmlsUF0krktT/ve+iAPf0SuDd77xw91cJk7IcwAeyfiNZWC7Ve4nU1U+ro0kLWKz
SAuLWh7AvT5JGhz3OA0R92C+HCPIynnPzzN+Lz0EvETEKbuMP26NzjLZhInrDEOilLeD0I0IjomD
8l/muyt1caCnj0tJ8V/T+N/MAks8z3Uu6c4WUlFV6+thZuqTIIOR9a4WxsPtpY30sTJjFKZj2qX5
oss3DC2bkMAlo/bLd76ITDQc97OmWdIOtpkvy03rIJxVSTsCxqEQtT0K9fN9KtnOn6qY9sybCNHs
4N0AehB+RKxpvSBH9EOT1Z3eGbDSRKYhGEG5hQtZlA1sWwYiyh6aCUqBMypmZfChF1xntgK0wNlq
osqbCIr+OMpMSNmkKrkDJ1CcnCDRrkG9UB4UveWflwzucNyZx73vSjolKhB1dnoxDRNxv/tL0mgf
enToNTvbjD9O0PsCNRZbim+guiZBSc7mS3Tj4H+LWeF90haSVqmXiL0r3gP8b+w8/jqQlgsGIb3P
jd9dS+NytJVIbwEASrq2LbPCJxwNJrNVm4zbX5yVeJ3GgI+qASJMeQKi6KxnBwACMI27yGiOgAk2
7eXxJ2xg5aSc4Pq2mJ5NkvX9oT9bgup7UH91tgptqiPyfh67cuuoKS0F6DJkHrGNLKxM1dJofdrv
3lNeT3SNzTeI2A7NKP5Jm1HfEQPaDldwRzMnK2Xz6a6dgxzBXWCI59moM7RiKXC99VWgi8u3P804
vWFbDl5ade2uQQfnMuA3fNMjL52glGN/xC146P/Ww3H4LI9m+v50r3UZhcvGrYRGqqVhfgL1AIyk
oTzwU8/MGoD4Y/asNZgNBGzY++v1282/3oWZRKJR26D814nZ65TtNGvWxV5YD7nDbIdxIG9nvwJD
Hu06v5zd69EZtYlsWcvI6eKHOgwdnxPOSUBbTAMV9mGMIt6JzjOmrbLR1VwbjrUyVw5ygyMZ5kJe
Hc/egbjMi8d4Eo6LPcvxpGPrpDNNnVptTuZjMnrMgYtva2PUKAtw/LWWrqGctLmxnKh7K3RTryvM
aYMEJAL4+F96dzsp0uBJS80LHt6PHomlP1qjPpV5EuNEgPx7NdMMku4inkD6+mFusS2m28m1YPsx
r6ChQvuPGTJvh9mydBK1pkORd3BcVeRkAMzy9bYrq0Cp4PmSD6ruezfM4OZDFqoMgPm5kP8drfin
swT89Y0Rai2muPJAwtxYxflZu19+2wT2vZ4/QLQEYX6L6GqfST7C0BR1+zYpPDPDl5cEOCPUCWmO
7c3/v/pwbzYyqwXyJZyedh6kixIqTbuIMmHH/kOG+VhwxsQmV3rzcKd7dXCd6dpGUd9/DkFMlNnd
SnJZ5JLqrxE0KetXBE1I2Y/jxN+/K5hR7F/OWtB/Aoea916Tmez0CXJ99y1n/pjWbDW7Zh+QQwKV
/n5ki4/pOrmV4R8iUopgizjNPuYTbDY2bKQGFbISaxGoslz+GgcAgAqRpG1/PaGak+S+EtRSatZf
eBqOBCbRNvQDjkL1aL/V9pezk/pVbbMLVWW5XB5atyf4INcUwKixKpTyfrd+G1Nj/RBTp/t05a3c
uXr6UFIPeezjIIrkhCGRRTKvVs4tONizWRjC4Jd2pzrMHjt4nElBCXarzsCs626y8BHVxll8eT+o
KscZOOS6SFZ61nbrKhti7hqVeJ646PSigHLcy8DYWaIfuwTHf/7BL+fbOiiRm0oMEEOWogb+osxX
ws2aIuksZfbk5k3e9TGDYoYxRrrOz0B4hWE6N1M81/kEO92WpYdH4KCw3IBR+T+TnHPmDcJNMIk1
UIAG5rom5RV+BWPlGehTY1RTUYeikcL5bA9ykVAmq6jRGzBJFt38aZeXB6pcOkWQO6QuAnqswcy+
vH1RBLIc5ZDF0/WP3I/tFVtyHKQwoTgfi5iFygGxuAY117vHE3/JGTQZYtSpD+buymVXGlYwtOut
ZgNn0HUvManJJA1+DQATZkzzrFG7bibkHKUudpaYrX4jvcCGr59gIkh1/U87ucPcyUf4no6++yh4
Ce2uVbNxgEsbTCQi+Y2DUj2+k9SmB9iN7muhD35VZsFh8E4BhuDIrF8BpsRZYJQ3X0VO6ZidSCyA
SSQfuCo1RYYV8OJqa2ayFcAdNDf+LC6VT4SNWivUs5AlJtj0aoBVtHWwsAFumgSqRhMfvXILxQaz
tHNDBg5jAi9ptbq8hllIpvQv5WgSQiBqIYY92J1UgjoCKyE5kppOyxNeAFSIo/ZiGcZAmUMZu+NB
JBjOgBv1mCJqjRONqdwJGjkZBzuLN4hJSCt17yoU/xMD7b9SSUWwsQIDGdgCHTblOyghPmXKEr6Y
ZDGjj6l1MsytK3HIqzUx9t2Kw8IclUIAZvjnXuGifbIGWkkzxz453wJx46M2UqkhxorRC/Wa4/tg
N4mUN0IGnPg0VG6dmT6QE+1GVRk/24k/psHQIIHZsg3Cq7JQAKABEAssDjyDvwh5RAxDL24+cH01
e5oKWT48WLZQAezONcLPlN1FaLCgz3PT5m/1auNQwu/x5MszIpAXiRw/4CrGwFQSO95peVS4KjjM
6th/QWziQgQEpoACAvC2HA2g68pJpN+Wgf7hEoI2GRv/MWPZK9xtNnBDjejJk9Ks30z6PQLlzkQr
bs4R7za/WZr3kfWfB76oPyxL+K5TTfdRBhl2taaBqutSMqGbvPplPyeJyFhqAvACIcLI19PVIzU4
L70YoMd1Iwnj+nwqShS3uu9GtTwAvbt62uSEkIU1LrqGUxkZ0+wL0pBpC2j2LGadaLntH/3Aqn/u
jJf8j9N6JMPeJpBU631FlW5ivRgOT+VSMBSU1CEDbCtkK7lxOe9C2M/4V/m/8RWlImn1J8MBERUI
29w5ehSG6TKIeJZPyMqbnm3GxhTyXnCq5Nu3mEqmoX6/ugqlg99An+5vX+IHmk0mVxZPNpskPDG3
YPvt2o+VxRqADo2+qzhLzTnPLII9+qmbvzAvtcwWdPmBjhxgo8apVNYuW3ULs4yoWAODlbA0AyF5
c5ppaOW+/eFix+ppgo73RxXLdU4EQD40WznO+3smXV0pBMWcMm+Rk8dvgOpSMboUbHWosnSWSvRR
bXoWt0LsF+HwcGgq1R4pC+aVeVUC1oCY/TBv330KZCFg2fRbNkz6FrlJ4IA/RXmlrz9/L48hkua7
/+Mdf3bBtjWKImnnakTX7CccbM76QYRL6/wKYnDFfUS5V02sF8Of7yGj/7cj6JOjuk47R0/xUK4X
dRU+nqAZ9LrRbNFM7aLjWTg1goJAE73L+o85ZFx9jFdEMkdgvrfngn7OEzhlzsDC8bPlE78bHqWW
tBZXy0+XQRe9QVoPWONK1TsKQcnCYo0dXjhSkaQ2UzSOXyvGyfacVmipOLgtxXxQvS+Z4JinGl3v
cAlAso+j4u4vm16WyAc31YfT7p1aQl4sfYWNpcNmjD7uoAe6gSszKIRfULSHfU/7H3B7cG6ej6yT
+IfwaQ/0QvOCh6q/w5ioybm0ivAgTSG0dMNEo2DR/zjPC/8EXmf62YuQ8dRztJhSTf8NDL/mkLeE
IZ2VUsY6ZkHYdLwePcQmn7Ys/XR+U/M6+eSONgRUgl45kPgFLbeQR/z6nqkYS9PO0RJeFuTW3kk5
BUY+KxSw8Xm4Dz+I5rz9cGzbzookmECYuKHCSb+cSoZiG7qdUCUDr/wkV+mU7Tf1/L79cTsqqCWL
JWrH1iidcvypsJpW/nprgfuifekDnLru7aM7u+jddnd4YdHYRRb0AetvgXFJ1ukvLPo+KmVnimDG
sxQLCuDc9TyHeghgGMrkV9TvWRB6VRAj9/H4Ih2Y/vyjQZ8r7tpUsMFO8HB2BS0HUlRoQdirbGI+
1d21UPVbUq32s1vGDyCpyasi+VGWxpZcS4qh5zr7XKxwK9iud+cR23ARh/nPpASql4KcqtpQQ1v5
JPTQ9WvQna5lntagg0+0DjEdje/ZgI/m3oOmxkfMhARggXUH/inH11vnb1nvl9ij5lO1w0ijsQtR
Zkgpi44nrQD47Jj5qm0xSg2Lj3ai0o+qPvDXhBnH4CuoascCMKMCIH+7UZxuqLbdhltpp4LeZnwd
56ZlAP7fNUuP79/bxEwz+Ex5uqwbtOlpT0SRK6HvIxmto4IhN5EdZ49tSIJqkjZVdhndOtxv+mIF
7VmlyhkTexFkYaYFFftfX0z8f2lOdCXtOkp/HT4dYimBttjeMxTB4JFJR5DWhOQFuhiuhkJfP3qX
jtRiSrZm0kDW9swoUkh68r/PAknZjpi3087viNJK/Nt8OMXfQqlpbzgjc4NDAWPrNO1fzXWdt0bq
1aLdCHu7k3wMyMjAzvoFr1cb4Sw/EGJA9pWXgEw/BQuw5kp0T4G6SBdx+Xj23RzOMtJhoSg2iGL1
+6eF3ebnDZ8bUEo0DJZBfN/wFQxpK5MqJdK7nRzzMEjp6kBa53AcAFjpu70++nq8WjpKlgwVyNBZ
ySSft0LMlOArwSc/+h/bCdaWMUE4H/GnhbzporawU3vWJ0Rt0gT996NxD5Rzs1duaAP0atvsuFZW
s5VsH1krDltH5DOD7CRX4txOcLMweai6p1LKwBc/oGZkzWJ7ORroJv6hQsbOVbBnhqcmCC/8PmOR
CaT76JqGWUxTMRySCq7C40XZXq7IXoyEIo3RVuHBdZIogx3w4CV9w3STjTUmwQOzDHq2kXTsSkLh
3zR8ReXi6kwrragZcQa753BlEiUQSxM8NwDGTNAThuZo1AfbpVN0P+e5v5kViZt9hXcTMYlyoUQe
Ac3GQVaCRrO62lKTt6t9Excv0bpx06HwMPelpMC0m7eoRkaH3UW5P+9TqqftFrg51KvriU1q9M0d
GYqMN/lGqj8xro8lThOYebQ+GxnVjjoKG6eSFAGgWD8l8z3OfZCY1mKo/O8WJG9ZtZBGW3I1qMiX
VltJWP1CP7cb/ukt9qZ2xgpjY1WUpN9o3xcpY/6SKDq1EfHxsAdostWpkMTAFJOoGYvP35HjsGzf
RJ92ZHMXlkNFyugiEES4roWJrDv1jE/Vkc1kLaTi55hcMVH4Sz0PXHU2RggeoTbzWi5yX+7yaPIt
nd0SpfHf7SfAvA/WQTHbCqYgKEnWGY7hUtckyc0RsGNVLlBiQ1Ymdmzm3X4WW1TxdomZjncEsstv
W68SEsnxTjyijHeQcSGT23hquC6N7kR906TDC9vObj0miCNsEmTwhSUbkyz6dXxxVYX+5IMz8yqs
WkunpjKxgtbwYPIwCvcdPr46bAbt5FxKKDoQw/amHMf0hFAo4pyKo3uU5waVGoeA8YYV0Eby77KN
pjTKQCkIdKai5Hcv6q4o4zApzyCnSQdQ20jmNyE9HRSu8E4geXGJh+m5nmmqXMbdHAwWvl5a31hB
OGHLos9Qseb3vNRsjogzixuF4zQPbgJzg3qkx1LRAdjkBgvij4oTqT+YOImj2XeeOJd1o+3V8lb2
g8cAX27ZR4QXBQS29Q8OjCMESyC50peY7kzdOcfV8wIQVzMiHOKMh9ZK0qQZ8gpczSdUZgY1cPWL
WXCe39KGcyoxyOYVFPAkClTUQkBqFLAb0P2AeZBnnWuIkRTmUKcjsGa0eqBjbswLdR+KwXNbZkb+
enP/ohnDUlYf7iY9qbdTVScX/bVBRr2lxsm7rVAR+kuELj3n5jxEmhR1NEsaWwDMV7dDkRR/nsT5
8LSEaAOOpJ03L2vprYc8UdxWFYZgfghRyay+eIxEuVEPTeZZfhJNw4HTJ+3Zp/jGJTjXXOqN3LN6
xTdOrtP76kRgKQLWDGHBQTcPk+aTdGmTBjNABjGE1qwNZ2s6GY3Nuu43yN+sB7Jm1aGyNa1UtL/J
AYN2Tktrq0qAX/ogKt2Fax5bKH4QzPdfMPXzQEl9X2w3EENQAmqTAB9oRg2syxQgBxpwnziZSBjD
RuDYHXX5sgX2+ctoqgLdyF/DfFG2n60lSOiqpprZI50UFaiJyAuAi/1YWDejxeqOf7/s7J009V0t
w1PT7kQbCsPKvfgEGiXr90XWEhD/8syzGFqOtbQdEMtkyo47z/suf7ZpVlIXjpTKZ+4/mEmz77sf
7hFSMNECS955lnc3T0AMskMZz8vms5gm2bZNlfadGwY5g6aHOWN2YKqpWRXgRcBgy8Jnx6QvFANL
9Rsd2PkOUbN6w9Q6YrD45w8HvZK59tqQ6oaam61cq2aYHbV+H1FnDvczyZ7KYw5pMOutNOiQdT2+
gequazFo062v60BKGLGCQDjEVg6tN7fHUO2XJenG+YnD3aRGequaEy9lkzZp17GmNWbs9daDMHWi
tUPFlK/g40qZ63+xmjLICG6yG9h1xJDqd2VwXJU7Qs+nQI81Wid3RAZxhv+Kv6KO3SkkJ0LlSCPE
lRyGfxfi5D76xoTIhLwVHbe6z+yyUSH1BSdvOs+EmBk5KFgGDPv2XIOsXAKsVc8leRhTEIhnfjAj
dLTHMeMo6tcBmHY2YtD0fiHP5xl9O7hZwZR3GEJCCoTickKHcEJkyLkT/8jYQAcLxnu3Y8w6nO/u
hPf1sNBYa2gw9qhuQSeBzUbjeczvIGK0VPQppwnLxLXHQIw7SM5dfZdaiPT6FoVNfdi7X1WxczVq
nzEz4wZanEo5VwvdfF77gLRWZw23XbBOXGiAZN4wlZqiq8R93ruEawmZCvkyVtv/87mNqg1rVmRS
sRp1+VMdl7lh1HGPcDbJ8oItXmVj51ZU8gEhlbqyKvH9CZHBN9hB66Mk2M6/1wTCF7yzJ8yIh1zX
LivQqLaWSq2VKetixel2rwLX6C9dIziUuid+3Gg9RKU/U0LysFJrZp3OGIFO7oBwKlD/V00FqrmP
CvIoBjkp5+EmzUyHESjtiq9uIRDliOUsYkCLEZWBEWg/hkUCI5Q9uiPIrLRBLVgLn3HEL6vuG7Wi
faODPv8oKWrJHhffxwzfkpPU3nENyq2NsGD+zvUnaszZWUsRQnhwKlI5dUJnsEhzhlMS6AbkuHoU
HkrBUEtuC/AyW4KU44IOv4jTbWg2bwRu8FGkUbxk5YQaN8IJ32k/rSn3O2UVNkbWUixTQv+IUbOd
h8tXYKhcJ8DHTR0DkNTDmTp/4wzvWoT8hlSPv+BixLLHzmltSvmclI4ccq/s7OxqYuYwNawZ+lr7
yfOLLNqBUDS+Q/cpWCIcB9GV0xd4kUYcd/Xjw7KStNCDABx+QqGMW54pVAv/XzigTbjbFMI7yA04
tUQO0XI2cpQBn9BZ8VpyH0W8eOFJDNTQSko5ytJ1hqYBbpqTXoMiecd6Sk66Mu7tlZopKQ+NIUPj
dYRvZpTx1/c5VQTl3RoOsb1D7rcwsFMy1saZJPsmvWXAN23SRXoND2ZY4IPZhy1z2fzPn2vIDB2W
hR6j5WnGLS/GSPDpXd8lNaX27HT1zEgGA8KDsNsoXVpcFRt3pB83iWA7ncNs6Q/o8WRc+aHmhD6h
EhwDG+1pmfIe6QhZF/YQ8WohjbJeIeAm+K2h3m+842Co4YszdN1sLotXRg31RPXVxzv/AzFOTdkL
iqsl5Xv72Bk8zMmIvYPcoYoaordQLrwmMLgniwdatdWrMZDOwZuHg2/UvKwvL8dqSfbmd2TFZ7Jc
XA6AWiZ6Wg386J0NEVWIwMmhomHZmChHZ8dvqRMa4M1bCOQ2JNoANO9ywHFBtDt4Aj3NuK5seQGu
nDYTGzaz4GAOEAsdanvwg3k0rq3YfIBCIV1VhmMJM6VuetkxOiaHdBeGjSMN8lLOJCzBgJhptRqU
nAubMmEtog5XneGVTSeQ7meJ6YMHnSPudxKJpPR+PYvqL3WabxByBJLSiA9DAiGPCUw9m9YH+Pl/
v7hAQIW4J/lnG6DEIwQbaviFvh6Aj6LGFQ95bRW+HNl84AgPkZ1V6KfC9G3SFBaNYc4HL44XpNzp
XfLG1tXg0SukXNYlNF/ebc2oCT6ibTkddJc/ZjNcxidB0XZGGOEJzN4ug+nFWv1+rnex0/VjkpPF
2d0SrB6IUFaU//McEjsHUTsmUE1eWzqCiPV930y2qAAJxg434aqwAtfQxNP/ApF6FpVdHeZZS2pN
apS8LJBTBfPOkBSSmA+ioeRINE47oAuQqsjLNGNzHmSLoYpU0SzitCObV2LaRSVDfTpvn9CcgUkx
UFCKhiYTHdQG2o3J7k7mo+HD5nLZjpthqQ49IZBaXUwa+JQJkkhOaHJdVO771kSS4uE54gxN50Eh
33ou6Osoc0Cpgzh+Aq0eURq3AGS0Zg/635hxvlCaoA0FqwLwOP9/LuQLk/dOpb0B4E4Bhs933vFY
8yCiT6BrhutVgmJ5nQLJJ+7RsE2JuzLyQuJwYMAKYrNUPUA/IOIZTR8Dz+4oQ6zZaly8oOWBi9lk
C4VyeZjAmAimalPJXhgrs1t8sKfsWKWECW2OrS0mJUsvQLKWKNgSoHsqgm9Z89/s0mcJT4tvCNP2
end7kWC+iC//tmJvRPf/ebbKQVcqlgNN0/8mbGSVvw25d+Ou0CACRpZL7HU2JlvOjLbgZYcrqy7+
qiipgetz5txHLaqTnfn8rPDWn603Q33yy4S5jMl5XEPEVCi90AAIkyn3dmDzKaapvWn1qMQk8sVr
ZrxSsRhI8171hdPCmmDRdy+AUF+MBLL6/D59hKl9Liz5bLofXTxI89UF4FlwqhboofMCabKlIAyc
V2GN13D6XT0fALEgyNMAGr4sFBbkP0MkITMGxZg7g36KAvxuAj4qb0Rkhf3ahKBPSvVNI0q4RbLt
bXICgcLc2hVNxXLfxO1nxL/R/L+II0ySBcmfg2oCmyO4PKlw/g69JMPx+f0qex/NoWbsw2iQ5ulS
jjBp/Qgz1x6wxzMSI87pwt5/h5UGSL6DD2/wvAod+h97K7GlavRZsZG4KifkNSxsS+OKe35xp9GA
+/V+eN0HpFXvZXCfmWJuIx4CdBI4/ZKHXmTOHNCkw/kSEGmR2gMrgeglrC/uSE22dHj7Y6ZeudWz
Q4P5Xbst0EcbaYYTZ7G9bvSzOdqV2iBz931LeH/zlnDfugjoFkatrLi0YVKGbhWdG/ojwR89uCqK
fVzxZwTJjg3/rLVaF3HJ1cs03v6+Ou25cjvlwROQaPzTNGHRGMn7nlHsp3jIXJEoqcHNjeRfGnwD
vl2xRxyrn/Cf+O+3YwGZXedQHdXpDrQtsVfycWmwa4IBwhj/ydf19+oNdW92HiqOg4nStc7wIAWy
eroIS2qnIZ3sUooHdpPLHaESeWycHmTlmA32bRvFKVt9ZQuUlsH9CuwEbRruCzVjfTWKC0M2CLdt
E7j0IoqnIURcgp14OUN7h7zay4ufdcrdhYnO4WFQWK6+LjhPzeIKXSVwFqQIutI4Swbhlzo3ekJ5
1miGlDzpncgTNcFS3Wzl4oUcp5dGZnG7uC7DVNZnNDaMgE00kX6TLlsotTFLbBg5mWE+SMdJ3vlF
VUWJPbtGdpTqNjBxCTY13DcD72oilTNJsMfysFRhwDZ+qqaNuxHQmY902hy+C6xGGEs+lwPd+oIy
V7ovr83ONrgej3AKnO0qurFPrJE6VUF9iTuiOZ6m0jPY7YJ3yab6tVI4EpGmmZJh3kMDvi8JuBDh
ftksfw+pK/DdlB5JSH+7vM2tx0XNdDLbUiqOa2BSZYpW1KavBpuZHZfdi6KR2J3HycGfOIbmnJT+
eNQmBH5PZDVse1FlEKNH4yOWL95QFEGh56AWLVmKjfLYNUBX2f5evPE3/Uf0RfbUyAYWS0Htaceu
rbbOBuK7m+BUFTm18SPfgsKilEEh9KAQNn42+E9QQQ62F8NKWffEmDepfuxIF14Ec0wSfxCP1Jds
ljSLrVXav8ba70qQ9VraQyS7b379Y+uuJwaD0rDaNkDeZlBvkaaxKZxTsLL3a04fG6R1ok/bBQ5T
t4QXnSP4F3Un44f9wW8oVgSPRqQMXffDU8rf0OSfDP39oN3pVAgxuWcGauzPQ5l+tWyqzWVT1bJ7
MZL8ChCxx9qRgRx2ff0wwQAcmsnA7oWlA2VEJp0qB5iaDItJsbWyyx94xYGv3K33qlpsx6DQEkmt
0zzSShVhJpXYQBKVpMJhBUrc6W/RF24/xo9OvqENyA7UONY4vGLnC4F1QhDT8/jwLk6e4ciJBiN5
VHrvJb8qwvT5PGi+eAJ0+O7xUrjx1W+8D9aQfWUOtw1dgIIo9Sa7LdjhV8VEO/j1U6kfzM+h/2YQ
Sn6VXWMaORIczUvHuBeDRHmot/GfaS/pc86PCMEr8XFw1g5ny46yX32ykcdb7tRIhb5Ndk+pvTis
zZxsSV6/1zBVVgUQiOotRtWMR0/9t64PIZyAwEsBg87oiIjlRkPacvII4hasvY8HVjByUEIryVs+
6qyUPAkYESh+E0QkK5fFUjDgshAD5gAFK5LnYK2lDGd3DgbtAPvfQjGT5aLypl0kMRjOcLdBkMUi
RoDRdadY+Z49A2oqG8freTDwuWEB3HfvclCvr6hfQ0EQwIxOZhDUC+JibjTACiFNr58Dtatovr+t
koml2Jtf3kNZbbQ9vQ7v/73xFosZEbMeuOkAarLmPNAOTeWS1Zp104YbqHxrnljJvghHnYxe9t27
QZwaTACWahu72X31OW7BqCRhmOYomHOQaD0hqKbQCCP9TVr/a2ATC2V9a4l+cO186brkA40ciXsu
ocWoudAFZjfuh0ivwzyV4gy3E/yiVaU8TpegnhjDmxhWC+z7QOgNMXCdczRxNCk8uiYyARZilkbF
Gk8jlBJkAwhQykzs5t7iTtCeRLU+wSncIFS4Vvk2LTWvzsl5b/XXFcME7kyPLzbKWJOJLNfgURxa
aKRr/G4lluU+D85FgW0+Bo/WsmxVx/BnKAcEeA6nFA/DkF5Zs0rQgOTs92EjUvEy0xT2uydvdmOP
iv2M6f3GxOnO5+wm1XYY/xwFIEcmzr1OAWZ5Z6KEvpvfB53xkmroa6uZlr10kcAT7ewi04FZTgMp
IQlcE05fwCVcu+b+CZYX8StsowX/AVw1fm/Vgb55qwIXukN452wIMmmr/8CftZ4cZWhcQXLmyz2/
28N2Uz1dx9g7x7tqx9g85q0nxTWcfUM2oBl1Envl2dF6IhdkZL9Y75D+n/MfWmopyio9VZSweoyO
9drZ5czUz7HBl7EBKb781Itwd93tVma6jUa2/HXsTd6F1CsQOfsPNxAgUEGfJgQVAMfwB7YQE8Yd
UOe+KGTYJyBwmaxGyotd27EnZPqtUhOcRPp4FkzWxRPb7E2VQBtobS0uVxZKj6KTcyvP/me5h3F6
EkHYIl5twvef42cnusGWC4SRgE6KxXNlib6pbn2iEPyxltFZlfi6u4sFuhh/mhWjZU++YUMGhuhZ
45QxMIJ+FI7m+ATvmkoWDYOGQyDDlo7fPkX8WgkCFaWLspvZ27zVHCDIt6vN1iAgBOhDLm7cAeuQ
g9EYidK/V1oS+yewdcN0fsGpC6zMOUDI9PlznHULEL7IWNlOlobGTghTWMVpKeFlak8b3xTwxvPI
HxNYjsr2Edt1G6qBXc3htmHcYtM2cSzPs1J06gJzqWA6l0z47RR8/ChWi8QeuRj/63muVY2dYs+Z
hK8n3k6r2KZsIJQJhEqQbDSmqbvgqJ32hdel4NG+yJYmZ1cBA+mvKEDl2Ck8dCknGmeT1/wwlrWw
2tgMz6A5oY4oiDRJm3VYXmTB9sY2gtqYFK9RUE7LpCEgtIryC0rHLcpbRBst2eCLVN+G1bka2f/3
VE09kmGTai1AEdcPbTC0ymgwPBWi8iaBuPjMeRRRc97v9fvvJLORFaClQpKFBr7qunzpQ+3hnMfU
XhLItyUdOz5gE9rWE3Q/d4hYYYVfaAqc7c9ALCngzW8C4Vf/YZI669GYgPegMMCmwziriad64eys
9JOkuyLa5Aqs4gFG4L4uxfMv6Bl4s57NzrBs9eryahshAbNQstv8XJjPI2+08oq3nwYLrSpoXuJd
ZBuge+r5lZ5Nz81YHigqsP6xZpfae1OTqvKMfZSCvrYh+ut29JEMrEL8HNalL6axShvIpo6oOPuX
0vv8/HvuljArE70f+3ppIn+tuOfU61IMZuYUnptuH3Q2332oJPPaKsTAOdGDmsgv36EJIZvE4+q6
zLAnqU6DTpSGtGULd9w0J68XVopnKwjBWly9TYr5FuU9gZa95Yfzud56YSMl534mvcxgN8vMbhPJ
ybuDsqOa0gxXZKcd5zY3HcTOOSey56FMPRyxdhEsejn2rllmHoGera2WAEl+RmIX3PgasPL/IW7F
7mAWn7s+FD1+i+rhDThKaOFMNzkO7tOIhKM3qK+rZUY1WRxActgiKuXI58gUE5+3J9YvzIHBdBr/
V5nhefB6Vrfv4px3uA8g0IWRpj5OdwZrK2Ex4XeQpj7mKxFGHpx0eli2aKGL1yI7XkQrpjUEK3uN
Iy1azwfnyX/5z0REgshJQljfrA2LXht5JLBq9vPgH5Jr3M37DsjgExK4Ev8fXALrjNVPMidmswps
aQKTev/r2RYyGlEXHxv1iNOidJlaSye3Tme+Bu9Q7Ir4Dh5C+t5sn/+Y7Cw/ck2IizJ5pUc2wkjQ
cZ/qPgFZAxYluZ120ZRN/FHZh/a7daL4o8fqOv5/4+nSMMbQkTOoyMfZEO3VZrTgBPQf/6ZYB85O
UqO3K4P0Uvr1VGlNmEUj6N5EosioS18R+Uq4YjTmgnbKtc5aVGFQPd0YJiX5PjUxXvJe8V6DrKYH
mIvzA08pVKdATv63/vb2C7HisT0fARfG481OFHVMyscWO/sNpz/YdnGu0SBpT++dtvid2V0Rm+ge
8CRgvx2ms9XBx663mtJiQZ1YMdIEkfQQqhyW+tIgl1Q2O26YU8FwNtKVXbivEgGKkMeLxaUzWvkd
8M04jXOPB3c51buwTuw1RqF5jV+/QDI16UYXuTpyvB9lLX+uPlGuNL3Dq6DrMD3kP/aaSRLWDsnr
7p0NrIYDkfhDSV0XUwTayEEGE61u5Kf5z1b6+bx4XNtBfCr/WAAB6iaY1BIpYJAt0hFWxRmUNiC5
T2AYiEEXhnkpzFxMsI2qXuKsalLY8UwWKOR8bVfBa/I1srjpG3Omo4D27LA49TzIpCv16+xHa/Sc
pjhGKNRffk3LU+B9mYGhTMIKKxM65phS4x9+7EtEUig7k68iyuuctf+uX7j1YLaO1wMb70//xIG9
jI6If3TWksK3FU4XoxmTZGex7ds9bcqW0hxInxFi2XpDm4BwpIsqIVDL0WZsxv6DCnxEXyoGMnvw
7d0stxR6bizfChQ0Ic6tSn4+lfD2KtWaG2yHUJfv+I+czouLVPkD+EebICPgxbIQ1gzX72BhIp4s
VgtgGrL5RGOEYL7oJfenVz9c35fGRkj17cw0UoewoHWct931mAXds5gTAqlcUE592RaBwJufapL4
tQ1+b5Q4nofRrXbaZhHjSWW5dFfe3KfxLjg2wJWOGf5D2yQTPWlW74SituGYo+yDn78vsao2MGSq
1g1g2yJhV8HSq9Vmt08s3IJkkcgEfIU+FvCixgxh90678ogfCDE2HI7HlsSZex46Q2K6kkZWQbHe
J+0+XJNsdA3ZzypLkoIT/8X8+8UEtyUhIcQ5taZIO+9QnNvZq7YuIzS2xjqrN5UoBkR0nbfF6LpU
BV2cu4vLgK58j1Sz9cT3qvyI8lZVWiQTFQYIgUwUZQ9LY9bCXVuRu6jUBGEsZbHAHvZNSkfPiFa6
ire+KTBXkfs3hEVl45IO13BzVI1mmoHAYXCHQ9w/du5F8EQruWrI86yAWfRjlPzYPMwHpFzWXZur
UfuSxDmdrar9SnjVUk2LoAJ9FkPxbcimpXiBbVY57CqcAaHW5oLpz178P87vv4WY4WJy0m7VJDsG
2fFu0kh+259uRdfUh5hN4zmSe+GJrgYMJoqywXEsHhpfJMrCaZYtmYkU44yz6l1L7wApRyEv/7aO
Fh7IkH4pcL1tClm2fj7hJf/2ZRj23bEnvjUfJ7EZrhhAVfkq/oXIojnn49ARYw0k/1qL9KkhTT0k
5xlcHFOZ/G0+mFgHvy2hZdoHebp+eXGZR2GtTKnmhbKM3GGG27hWOPYrvJdrMiq+eOcaWyxxbux2
wjY8ht0twxfokcO+WxlthFNPtJ7e5BCQRq9qfPkc7IdqWU9cEHLRaECnq2zA6tSW14tQwxXP8/6G
LJGWOW133idQVXDEDM5CARjDI7s/DjYiqgiKbtMRI/jfqAs5fIwitZJYLjO+e1iloy9Tb2IbE7qh
RWmVoZzSOYnoGaLo1JzszaAawYkKeZBw7ekKOdCDPdGL9CqUUzSMXHNNINXhRGuU4WSNckMpnF+q
6/UbnYPSLW59EMj+MCl5b7jli7KlTAbvfzCxP+XxSSwsDnFIjl7uHYqg9VH//GDlok9rzrWu2MXh
copAyCZwYH3ujUWcBTaHZtc/DDABn1bwLxw81zVtX0FWY2ZydIbP5AYe12QC2KihgRlcjXfMSlaP
eNlJpMjND2tLJQuvVT0uTDa0bRPsxZW++XcQE+2/AGZ1KlyWXq966lpJ2o7ne4yU9bUHTrJMk0Tq
vl19HqWPtZf5eO6AEVyz0MBvtWsnMWZVtUzTo0bXNB7Jpi/VHbncS4d4CGf2oSwlj2htHmc1Ne9I
YYACDrOkEFfrIfxz5OQm04GNowf6pWv6W0I8/5ntrYqgvJId5/K+gjUETO0qXNYS/EJfdVIWIHqk
IZIP0ZLtVQ7eLUgR0osgXmDdkqlp6hbOVOLLm2hCjE4zsQNRsLHunZA+oL+Uww/lFdKcBKE9a57g
vQe4Y4Qt9cifK5poS3Ylwkyr1XDd1Bo9x4zmU5/wGqgvKTUX4/rJMtkFaKfK3P3O9t0+ztsXnEat
DN5ribk0ZBGOdx1R1ZoTwvL/+dINKeH5+iNUBHgYZiBHqAlMQG03pObUUDDEBfeIZTrY8p7eWzxH
h0sCCcfUSOEBqLN/n+P5kHUw+8eg2NUk8vgej7I+ovnPTPI=
`protect end_protected
