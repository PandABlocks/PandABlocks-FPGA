--==============================================================================
-- Company        : Synchrotron SOLEIL
-- Project        : PandABox FPGA
-- Design name    : sfp_udpontrig
-- Module name    : arp_layer_component_pkg.vhd
-- Purpose        : package of components declarations for ARP layer
-- Author         : created automatically
-- Synthesizable  : YES
-- Language       : VHDL-93
--------------------------------------------------------------------------------
-- Copyright (c) 2021 Synchrotron SOLEIL - L'Orme des Merisiers Saint-Aubin
-- BP 48 91192 Gif-sur-Yvette Cedex  - https://www.synchrotron-soleil.fr
--------------------------------------------------------------------------------
-- IMPORTANT  : THIS FILE IS AUTOMATICALLY GENERATED FROM ENTITIES LIST
--              DO NOT MODIFY IT.
--==============================================================================


--==============================================================================
-- Libraries Declaration
--==============================================================================
library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

library work;
  use work.arp_types.all;


--==============================================================================
-- Package Declaration
--==============================================================================
package arp_layer_component_pkg is

  component arp_req
    generic (
      no_default_gateway : boolean := true;  -- set to false if communicating with devices accessed
                                              -- through a "default gateway or router"
      CLOCK_FREQ      : integer := 125000000;  -- freq of data_in_clk -- needed to timout cntr
      ARP_TIMEOUT     : integer := 60;    -- ARP response timeout (s)
      ARP_MAX_PKT_TMO : integer := 5      -- # wrong nwk pkts received before set error
      );
    port (
      -- lookup request signals
      arp_req_req      : in  arp_req_req_type;   -- request for a translation from IP to MAC
      arp_req_rslt     : out arp_req_rslt_type;  -- the result
      -- external arp store signals
      arp_store_req    : out arp_store_rdrequest_t;          -- requesting a lookup or store
      arp_store_result : in  arp_store_result_t;             -- the result
      -- network request signals
      arp_nwk_req      : out arp_nwk_request_t;  -- requesting resolution via the network
      arp_nwk_result   : in  arp_nwk_result_t;   -- the result
      -- system signals
      clear_cache      : in  std_logic;   -- clear the internal cache
      nwk_gateway      : in  std_logic_vector(31 downto 0);  -- IP address of default gateway
      nwk_mask         : in  std_logic_vector(31 downto 0);  -- Net mask
      clk              : in  std_logic;
      reset            : in  std_logic
      );
  end component;

  component arp_tx
    port (
      -- control signals
      send_I_have     : in  std_logic;    -- pulse will be latched
      arp_entry       : in  arp_entry_t;  -- arp target for I_have req (will be latched)
      send_who_has    : in  std_logic;    -- pulse will be latched
      ip_entry        : in  std_logic_vector (31 downto 0);  -- IP target for who_has req (will be latched)
      -- MAC layer TX signals
      mac_tx_req      : out std_logic;  -- indicates that ip wants access to channel (stays up for as long as tx)
      mac_tx_granted  : in  std_logic;  -- indicates that access to channel has been granted
      data_out_ready  : in  std_logic;    -- indicates system ready to consume data
      data_out_valid  : out std_logic;    -- indicates data out is valid
      data_out_first  : out std_logic;  -- with data out valid indicates the first byte of a frame
      data_out_last   : out std_logic;  -- with data out valid indicates the last byte of a frame
      data_out        : out std_logic_vector (7 downto 0);  -- ethernet frame (from dst mac addr through to last byte of frame)
      -- system signals
      our_mac_address : in  std_logic_vector (47 downto 0);
      our_ip_address  : in  std_logic_vector (31 downto 0);
      tx_clk          : in  std_logic;
      reset           : in  std_logic
      );
  end component;

  component arp_rx
    port (
      -- MAC layer RX signals
      data_in               : in  std_logic_vector (7 downto 0);  -- ethernet frame (from dst mac addr through to last byte of frame)
      data_in_valid         : in  std_logic;    -- indicates data_in valid on clock
      data_in_last          : in  std_logic;    -- indicates last data in frame
      -- ARP output signals
      recv_who_has          : out std_logic;    -- pulse will be latched
      arp_entry_for_who_has : out arp_entry_t;  -- target for who_has msg (Iie, who to reply to)
      recv_I_have           : out std_logic;    -- pulse will be latched
      arp_entry_for_I_have  : out arp_entry_t;  -- arp target for I_have msg
      -- control and status signals
      req_count             : out std_logic_vector(7 downto 0);   -- count of arp pkts received
      -- system signals
      our_ip_address        : in  std_logic_vector (31 downto 0);
      rx_clk                : in  std_logic;
      reset                 : in  std_logic
      );
  end component;

  component arp_STORE_br
    generic (
      MAX_ARP_ENTRIES : integer := 255          -- max entries in the store
      );
    port (
      -- read signals
      read_req    : in  arp_store_rdrequest_t;  -- requesting a lookup or store
      read_result : out arp_store_result_t;     -- the result
      -- write signals
      write_req   : in  arp_store_wrrequest_t;  -- requesting a lookup or store
      -- control and status signals
      clear_store : in  std_logic;              -- erase all entries
      entry_count : out unsigned(7 downto 0);   -- how many entries currently in store
      -- system signals
      clk         : in  std_logic;
      reset       : in  std_logic
      );
  end component;

  component arp_SYNC
    port (
      -- REQ to TX
      arp_nwk_req           : in  arp_nwk_request_t;  -- request for a translation from IP to MAC
      send_who_has          : out std_logic;
      ip_entry              : out std_logic_vector (31 downto 0);
      -- RX to TX
      recv_who_has          : in  std_logic;          -- this is for us, we will respond
      arp_entry_for_who_has : in  arp_entry_t;
      send_I_have           : out std_logic;
      arp_entry             : out arp_entry_t;
      -- RX to REQ
      I_have_received       : in  std_logic;
      nwk_result_status     : out arp_nwk_rslt_t;
      -- System Signals
      rx_clk                : in  std_logic;
      tx_clk                : in  std_logic;
      reset                 : in  std_logic
      );
  end component;

end arp_layer_component_pkg;

--==============================================================================
-- Package Body
--==============================================================================
package body arp_layer_component_pkg is

end package body arp_layer_component_pkg;
--==============================================================================
-- Package End
--==============================================================================
