../../../SlowFPGA/src/hdl/slow_defines.vhd